PK   �<�X�|=@�=  Ȍ    cirkitFile.json�}�7��_��D��;,n��닐���lKa�㻰���n��$۲ס�~@_�@1�I9�=�V�� ��D"�����"����f�Eq�K�XN糛�D�o�%��C��m<����nW�۷���������h��}e����Y1[�&<)3-��ZD�PI�d2�4ay�QD�����Oo�''��W���}���q��<*9M"θ��)�(%�0�g45Ʋ��p�3�9�
^�9�4�M�ȢLsS�<Mmýe1�����nY��X&���Zs�X~�n=���HK��H(�#n�-��:�"�3��T橝�ކE)�(��Ј�1�LLy�&&хHr�J_�MF)��
F󈧥�4�s�9WLe�>&���)
�ZN턘��R��QlbC��n�%��$fDX&��̕� n����q���/������]���)���Vĩ�[�YFJ�������H�v��(%4.U�ܶ��a�[�$(bIp�$C���LOY-�Hhf��Ԃ��I�2�y.c���!��If׼Y�UZD��"�i��$�̂�W� <sZ����YL ��瘦���[X��*�mٔE�$�ٹMEQ�`��-D�ԐIFI�i4d�2�jHu�PO�A(E:��"��Q@%9j�-���E��2XY��Y��[�3mŌV:���ր��4�q�U��8��b�6��FF�h�x��ɰM��"5���"QV'��i���4#)#��@bdӾN�W��(3��-�䑡EY)n��L�P�k����NKJ҈���6��m:+Ydˊ$%<ѥ@6�=k �!�#�)E.S�[� �uj��e
j%��F��AQ�["C��a��H�3߉�(���	̖�QM���H��̷�@'"\�ȵ�|���b�#�)'�I�(�s�SzA';����ݔ#wS.���K�\k��	��2T�P+|�4C5��M��%�l�J4�uߖ2|�z�\�·%R^�$e$il��e������*-�!,��-Q��z��Q&}��4�"}�Դ@5�)$���%J�(�kM��h_@�pʷ�@M�P��L�<`*$��
�z�D��mN ��QS�3a��F�
����?���P�\#ךF�5�\k�g��>��=�LaFD�h�D4=0��>�訂h�w���`���ڇQ���e$D6���p_�A
�� ��B�Ѳwma�4# Z�4�`��Iq���hZ��@�3���4ЛѴO�z�!Z�iY@7�3�,��F��:��V�}��o�+�S�9 ���L�wEC����@�3�8Ո�X�� �bѷc/D13�0��Z���#��\m�QRheRd���z\�aa�Z�)�>���3�p��n��!Z��3ȅ�+ ��Y6J��Z>�.���(�>��
Ӵo��'1g����̷k M��^�'�}2h�Ŝ�P�2�H�n	4�c�ڷ���U�PN`Vd�T��>˙�������{#w ۾��4G���" �y_��>�3��i�D#�!<(�,��>�3"pŷ�`3��7`>��3
a��q���� '��Хc��M��r� 0����\��2�D�h�,�`��Fa{�>��1�nj��D3�H2��	f�i�w�
��|n@�aL�^�",��0}���O��c����`F�w�&f9�0�iT�X��jڥ"��w�2��_��|���j)Kd-����U��#���j�,c�'�P��dTg�Ġ.xà�T�EZ`����8�
Sө0&�^��)�ج1L쾂���!y���jL͍�SO����-�DS�a�	$��a��T�4�i�b-ܦ@�(V��H?��tʄ�u��b�,�*ŬB�J����Eō(��TS�8M��u�B�R<�UŬBq�g�5�à�W(6Ek�v�i�	�k'j��ad1#�y���ъy�0�X�A� �59�ZW�x�OUF�0(5��%���@CW56��1;��P����0(�aE1F��
Ū�y��Fq�J���Bq*����0(�aP,�'��bF�0(��E���bU��4�欩���*�^� X�A�
�b�̶F���4�]+�93�]SU(6q���q-DS�2J�0(�aP�àX�̈́g�FF10���m=�z��P�aQ6P�aA=6FA���y��408 /��q�;|����o��(�aM;|sn����44�tج��K�#�͓/1�d��.0Fs��h��p-���хF4>���7I�=Q��
4�ihР]v�H}�l �4�ox\��y�=��9�H�0w`?���܅�ۉ��e��h����5l$�p����X�&"hX��Q!5l��;�e�qKd0i��'^��� �;�,A�B�@�n�y�F�;!@�a�Nvπƙ����8��p�#P8ư4�‾�����J�uи�a��a���ã�-�4N  /���A���@7�a;�G���Թ~��'?|uyv�:��#y���>lQ��x{>@ݵ��s�^��U�u���Er��� �� �� �� �� �� �� �� ��0��0�%a�K����0	�`�$�I�0(�aPL��0(�aPLà��A1�b�4�i�0(faP��aP� ��A1�b�,�Y�0(�aP�à�҈à��A1�b�<�y�0(aP, X�A�t��b�"�E�0(�aP,àX�A��b�2�}"�e�0(�aP� X�A�
�b�*�U�@f�0(VaP� X�A��b�:�u��(��^�k9<OP�k|-�g	�z��%�4P���Z����Z��z��� ^����Z��z=X��_����^�v���r�G`���q��^�k9<GP�k|-W#��_��q�^�k	3.���z���5���sv���rxW��^�k	��A�]�����:�^�k9������Zj�`��a�u���rXzC]�k�^�k9�#��5��ü@]����z��2G0�k|-�5U��5��0�>@]�����׃��]���#��5���sv���X�@�k|-a�� v����Z�/`���Z����Z���ql��uU缾���<&l|�a�(���wIV����|����?!2l{�݀��7�ަ��<�#�ed�$LӨ71�iLaEPMcr+�0yj�f@�b�#0-�V5�Ӵ���k%T�>���h4�.�$O����D��iTd�S��<2��Qlezi�4�XE�)T�-��~|��~k���υOB�;��S��IpJoµ~���w���%OXR8y�m�z��uv>���Q5�U���J���r0��%��9���/��G������`ZF���M4��Z��ޔ#z�ju:�Jo��^�{Z^�#:��-����e?�p��=-o�1>��qI�<-��1�{O�@��^����"Z$�;�	�����]���~���(VP��+Q1�xs�u��k��,:�/����毇 �������x�0bU`Y����X���64a�ЉJJw�#�%>+ޢ�8��A� ��P�pb��>��P�`~�>M�{�zо���J���������u�U���Q��q#ϑ�{�x���u�n��õ���^��ֽ:Г���lԯV���['Ǔ$�N෰�E�yq��Kz��k��\R#z�X��j��۠����%~�QN�<��|�{���}3���9Lu0'�s��`.�g�30��<���},���p���k�O���Y��¼^On��t�E4�՘�~��ɻ����|���oy/Z�N��H<{�l`�A��O��Ҙ@_�a�1�O����1�N�M��y�j�s  ������qX��=�?`h�i߹	�hYp>s?�d�i^E}��2�v�IyH��b��s�i��Xߑ&̵���oA��0MHd ����F���9�9����`������YO�����'�J�7���E�~�K��&��/��'���	߸�}\"�� 6��6��6��6��6�p��K8��� �9��!� ����5����NܰQ�{�@���,y�~�W���:V�|R�����ѻ|��1}�!����n�(�^w�� �|����X@P���N���NA��i�|\x,\P7~,|�LG��U�!.s�Bs�>�g}��s�=�gc;�.cs@s����9@[��^g��Y�aL�� W61�b���xA������b/�3� 6uH S,2�� �H$�g �O�l+�Vd���d	�CO� 0���� �kd��K��3��<2��%�2p�<$�s�u�9�?_$A
�����#���)7o8�_ �2k��'4y�uG���44���� �Q)�0F&�J��l�� t������f�Nws6��zs>���f��s�8�\*�� q�LH��g"@~<�����-�D��9x&���^�a�T��u�����ʼH6�a��K%
�:����b1x��@r�T����B�+�T�0\`s0����)،La��&f
�6?��M�t�;`����y �6�m����w	L�4�q�LNg���&t:�@�:_|]"��l�'<�dOx�9��`S?�9�f��.��,�?� �H5<�5��%�D�l��  SF� �9* �Rx�y�6�����SK/���f��/���@>��v]z� 0/�N��K���\�F���T�Y,5�{#���D���N5R��Z�:Ď>�V���TC�Y,���c�����.�O5V��jt ��>�� ��ég����`G}o���K����݈����;�u���Ynp��d����s�;����q����v=Ǳ��Oȇ��_�E���	�w�lW����gh�A.���rpc���t6�]��Uq�x�y^�u����4�y���mŶ�[̅�<E�g�|��A�u�è��;�e�� ɎR�L�:�`4��`&��#��O�n�9��X@�.��CT�>��g��.�9�o9�ևAE�o� �[�j�#�Q��]Pǘ�(���.���S�V4�8e=�F�0�U�uQ��tb]��2,�Y�����jN�3���Q?0��]�e��XIͱ��KlX�cQ̱�X`a+���QW�]�ƨ�V��X��ь���ԇJ����	,�EW4STn®�L1&����t�]����X�K,�%�ԁ�+�%Ų��3����區U�V�VX�*,N�
�S�#|Q��]�E	{d1f��=��.h,�5��b�=
R��J�J68@��!X:Q�Q��4hu=�x�z�T���!yKb 5^�{{���N090t�����G`�k�I
���/ ��C�`r%��0����?

`6����.(w����²����j�U7���
C��{`�b�����S.1�Ծ�<���:����б�@�v�P�S����\����? hu���� j/t@�]���r��}ȡ�I�c(�r��N�.�P;!0�
j* �IKcX��)�D*�q���g�Cx����p(w��^�[0��, �T�I ��u!�l8bf!�P�)�������z�t�*���P|�Te&x�
8��4��@�����,���+0��3���	L��/��^��@�J�i���.X�&�0������ �3z����fW�4wQ����\�<��ƭ`7ry��nR�lw�����J:W֘��PH�Cn%����_��+�^��W:u�	W�u���(չ��i+ձ:UU�ZN�DV+��o��j3���j���J��*1q���ܕ�w%�+�]	�JWB�U�]�����p%�+!]	�JHWB��'WB���n�+�\	�J(WB�ʕP����֕P��r%�+�]	�JhW��̨]4�Ĝx2߸�<l���q�,%�Ӛ-�x�ee��,�Vy�k��J,%���l��VO�
$�����U�^�E�2�FQ�u��g��<�:�L��ϥ����aW[!XlR;�k�6��`ق��m+Ѯ7f �M�����"{�$"����E,u���SZ��L�d���<n(�������&��v��$Qb����Zg���A��q��ɚ ǤF�ɥ����D� De�'Do�]�}$� [�^��>�Po��b�v��z�[j5�ߙ�����7ط�v��n�o��p�0�`ߺ��c�A�I�S�j�������j�'���≹��0�>�[l��!X ��vs��G��r��K���:s逹>��Of�1.2�q��MhO:�)yt���p��2w��)�x?q���p�ww���×xoq��a�"���HQ�����쌍�r����+�nG|�z��6����Q�Hު7>~�fn|"�"��:��D�Erv�������p���y���'�/���Í�p�ͅ��S|cs�� v���E^�ؙ)ߩf�qn�r�ۦ.�r�67̷O]�5?n|��E^���ƷO]��?n�G�K�
�Í��q��u���S�xEB�X� G�f��aޯ�z9��8���=��b/�.7���ʜ7���������hR4�n���M����f}(�H��7>_"����uU����K���ݻƭ���7����{�	Y?"�Gt��v��#�}�׏x��X?�Gz�Hw�-�]ɆE��lx$]&ɆI��l�$]6���3��Y?3�b��'�	 �b�[�n��n9�������Ͱ���Ͱ���Ͱ���Ͱ��T���g�;d�r=��)�-E7X�]���h��h��h��h��h��h��h��h��B�&ی&�&ی&�&ی
���ی�ی�ߌ�ߌ�Y|^H�����aeTrww��:+�w���INf�������4�;dZDV�,�R
�yj��e�-��~�P��m<����4ۻ}�w>,D��iTd����<2��Ql���pi!��mꊨ�uqץA9��KaK��Ɋt��]���7{���g��y��^}�r1�/�i��J��ϗ��t>�"��ʤ���cc��T
[��=��v��$�:WT��&��'Y[}L����#ir���?�Ųj��o���*�euE O���|1��$5�7�(f�EvW�{��t"�ZY.7�"$�w��&v-i�v_12Q�B�z��N&B�!����T����H�y����N�o���<]�Z=���v�nȄM��x�޼�����X��j1��W̒��{:��%�{p��UL�Ǉ�Ԣ����|7��b��Vz�L}�,��.��]��nQ���tQ�9[YPZؼOfe���b��}�O�\<LW������=�s�D3�������Uy�r�H��2ʋܮ��舱LgNX����]��- ���K������׻�Y��ުh�����!"�g�ԓ�-�)��ΫIdB�8�j���G5d"7�dTZ]�`v�$��$��՜c%EJ�ebW W ����a������
���f���Q
��a���(`}X�`�1�>�N�j��< ����LZ�:�h/]S��{���KԞ�^"�I��b�TE*�Ke(��ĠʺMJ�T���>��H�uƴ��3;}D݉H]��t=���Au/]w���u�\/�+���+�����=�>��d��DGc�#���>�O D-��ć7Ӭ�_K��FhWv��PP��Y�'�ڀ��6���j���hܔ1 2�MIXm��TQo1�7i@�I�����������]�^���������=d}��!�CoYz�d���!�CoYz{����Cև��>������K֋��>���u�[��rw8����]^,ƿ����o��Y�\��w�oƯo�y�7��B���8�L��H�J��0j���_����������uY#�=��"Jc�"^�e�r��ТL4'B]�u��+��Ќ�Qg�-��(Iuf�mF�Ҹ�Ŷ�����j�p��2,�#ͤv��(5q���q�ڶ)�;�|>��pU|c��������wӻ|�fFKEuj��b��̲ř��)��Y�tc(�&��|�⾘�Ja���Dʝj95"2��)L�e�%q�����n�,��I)U�[����f�rC���,�$iB�������,/\9w��߭߹����~��������/��IUz���L����/VO�|Q,��g�V]�D���]���-���'��2�4�#�%yd��eǆ����b$!1qQ�,�ˈ�G��""�ɵL3CH�1�S���R���ځ�sp2J�R%\d^�&m妈h�.UfuW�*cq.ˇ!��_��e:���b��^>���_�_���z����^j*�ӯ��G����j���>z���~3Z��|1����d�[���.~�O�V���/{�_�_�-��n����>��h��(��b�r:=��fE�L3K����1Y��7�,y[�/f+�mf	V��l5��~]�Rܹ�_��ğ7��w������i���������|���ӷ�V�����r��'�Y�]��̮�WE��^�� \����"���'-���.�~�oF_�>b�xĈ��������nL��}7��l���w˪�Ȗ嶌��I��j��t�g���|��z��\�%w�xr�,�7H�MM�?uj�'BZ��n�������Ȋ��Q"{7�U�Yd��bU}klL���[��]����r9�-��ׯo�������W�o_�z��}��KM}�,��n��O^����w�Ru��J8�z������b��w�ǯ�������¿����Q=�";�������]�x4z^����d��W�=��O]vQ�m��������5�ݫ�o_>�v42�ݏm���r��aQ�$��R�y��.��p7�ޗ�����.;�4�Y����U��c��������?<f1ZQ?Y,��F��h����mf�􃛯]�����v�klׄ�M�߬��k��Gs�Krgq�W�n>�k�=5,�&�{��+��j���}jgn^��\�����F�5�=}�u_��b떴t��?�����W���F���J�:���_��z�׏���>�K�__�(�Y�_��z�{�o�s�~���z�׏���Ϸ�<�`W���Z�o��Dv�ݟ���j}T�خV�l�RˤM-�O�����t��J�S��\�XOգ��υ��}r�ȍ�g���M��j���|��^�|W��蛹��z��o6���\�����m�*�7���QZ����_"�&|����"-��ܖ����M���#_6��aVmx��Vu��[��[����ţϪ����FɃ�l5��2[�g����z�߯e�x��X����n�V�=22���чwN�=�������?&S����[V�F�V�s�6-F�/���-���c�Ȩ���+K<���I����Ѵtm<[�����Z\sx���}7{�D� ��6U��ed6���U%+���ͺ#;`�����-3�ʦ[��m=�W[�ݴ�u+��f�m5���Ɗ̽��aiG�_�������~������ٮ�yq���Hl'��o��d���.��t*X�UV��)��ս�U���(�U��5T}��g���>�h�i.G��1r���]�ˊ�~:s�V7=���߯[ܐ4�~��r7�����ӦB�_C��y*h�q���4*O%E��L���R���z��	>��]�#;W?WTQ8IV�${�����&�����z��kd[��|Yum����jj9W��S/�N�������?̜�kmT��˧�nq���y���~�[�h�皛���v頻�����b�p_�z��k :��Q=#�7U=ʧo��ĵ��|�m�
�^�ͳbU�������5�[���ycǸ���ƚ�}[ӏZ1�#Z���[�8�Kyݙ���;�(~aa���|�^�;V�����Wk����o��z���g���ִ٪|{<G_|Q�5�S}S�p��ilO�-���6������v/�n����C�
�,
��.�����6��h�0s+�]���\|v�����[������p��l\�?�fⅭt�Q���j�m��RL&��#���V�� U����۵W���g�*���u[K�͒�6���F�(^���y�������w�wN�ȧ˝v��VD=������⃛��5���_�u� q8�b��l��O+X�D���=q�Q��O�J�j�t��82����'is�:}���4w�}iK��w�k7hOk 6Gg�a�zg��;wm�}�V��V�OV��|�?��p�ͪ˿U���o���QeD��d���8�xZ^�{�pu��(����a���J�+[�ў0����ת��W�j�+i�h�lnU;���wE�Vv���w��p�"�$[xT��U���ooj�v������ͱ����}��va8�n�-��l�X8�ΣEq�dE�����Z)��Qg��϶i�Zd��m�+��P�+I�dt��uk�w���|)M��PI��{��ld���[�է��r�,��Z�(�����#��[;��;��ȋ����}�Ύ���ta�>L���ޜ~�*���V�'��O���E�~��%4���NG܎�()��O�y��*�Z����ݞHɚlT?m��?;�����"�a�-����6�FS���"Z�:��wNk��[���k���x|S_�}�B�^�]6�=3�X�Ε�	��v�pJ�w�b��Mb�xH홻�V��W�F�TG��s�!�~nGêv{�m��6��ͺE��?��lh|S�M�n\S_N��{�m�*d�I���gz:���{��i��F�/e�3��]��I��y_#�m3d�z���}�t���vy���*u�쁫����m�<>X���=֞�Mfj%�U���k:3sI'L+J45:f��1!LL4��"Ti�}�f�tW�F	3&�I�#^hIR&	gJҸ��5C�L�k>e�6G�y0("�G��I�7kG���VJ��ϳ�v?-"C���(�8�Ls�zʛ��Vm�ұ���y��y���D��b®s�^Vǡ?�ܟr�r�P�'B*jT���㈘	a1R�΋G3qIJy	Ig��pJ�F0�'V�ĺ!�=w���H��rJ��I%��\���KA	��%��:;O��4�|��h��'�}v1��d�p��y5��<��O���X��X3ܮhN�����Y%F23QT�m�a1=�L�g�2Ml\�����n�2%�\�LE�yT�ª�"�#*L�|�O�C �ɦ���L:OWA�Q9��i;g�=�Ǐ�ld�h�&���+���4!�۱+##i�R��D�L�eZ�2�SА�ޥQ����rہ&��K�&�zl7ډ�J�ʟ�=�KEP�yn�M�Z��
��ԩՔ*�.�[K���I�j͙���箠��Q��!��JRr�p�q�X��cJ���()��-ͭFQyd�K@���J�"��L���ˌ�	zI ��;݄�v�AX?Rb���͡�D����<�̒���V���S��S����'$�9�*�VrS6�(�V,�B&��>�"zU�y��d�w/��1�[�-�_�'���z��=�{@5��3�n�ԉ֔n����e��O�VyĒ���&+'.���A������8�/.�z������;���%L�ⵅ��q�D��H�0�3���(��#⤈��Ms�Y��� z�$��"��c���'$'B7}�)�zm �&p꡻���uq�� ���q��b�ckBbM���l&���1�(vc	䍕����������GĆ�����	l_?�/~/��p7�,�zX((9Q�t��z�>��G�2e�Ө �Υɳ(W&/dQ�����@�$���m���f��Q���Q���Y��e5�� ��Z���!��?�uI�e��bC�%� d�V�$�Y���>�?�YR\If�ކC���,���YD�"���6�,Ea�R�y��R��D+e��XaG�7}[���q���H1�F1�\^�XGy��$˲TeE=9@ow������BwY��+̶?�'�D���:���J�A��I��O��W$�7eTM���i����U���|�
����Gf��;UKw�ܴJb*'�DiH,���e�,�EDK�~(�=/d�Eǹ&�b�9����*H�cu�z��˨�� �w��8�Tw	��"��L��/؝4�m��A"f�T%�2Rշ�j-���!޻B����i[�
+5�\�i�����yԷԶ�-&	_����z}�ݭ'̵�pfEU7�;�:Ы�CMk�VE�;�E�F�e�����d���-,bs�!o����
�\�ujG>��7���}��@�ڰO�|pIE�Z����ש#���E��02���u�V��=:��8�'�A�[G�U��8P�f���.�IfQY�쐈F�����(U�[�j��Ds/S �JSNh��=;^������fh+�\�tn�0����*�
b$v~��*1��>sn��n��g�e9�#QV��i�*.��Pj�u�	sq��=�A8)3^o���z}�{�[�d�Y+'�>,�܋0�����Ws�����d��*ׁ��\U_:��0���/?L��;�-���4DW��w���pb�19�x�N���)�[�;�Y��+�/�o�x�(V���9->�hU�{��.��|Q�Be��:�������t�N���rJ��ne�6n�V{���Z$^���������ϧ���d����w:�^��|���NCK������Kn�ڇ�#�P�QU`=�*�m��̲�����7-� *˘�<$�x8 	@<(�����&�a����< �� I��I#$�D8 �80�DP ��;@DA D �`�*%�dN�Ҧ_�T>i�x�B���f40YXiFO#�0���쥊=�� z�ʻ��D���	�v|>M*c��A[;�L�G��Ah �pw4���Ah��;���Yg������T��
 ȸ�� ��Utp����6�������P �R�V]e�9���n:�[wOӯj��gK���AɌ�I4 p[?�� ��&XŁ�!8wǪ8
r�oQ��x�<�A��H(f����8����c/ �����lS�x��˃�.�ZT�)�Q	ًٴ�����\�<��#X�*h�+��<��vgpM�[oO�ۯ�L�/;�t�a}��HvTB��\	�G�v]T��>䒻���o��x�\i�=������r�uail�m*BD�.�&ہH�G��S����X;�AL���y�N�ś�D�n�r�lQyN-����d�y�>-8B��7���xw���O
�������uV�'4@���#��ݕ��O!�d�ͳb��ua:��_ɮvkW��Z�
n�44�6�Ϝ�9^O�d���cu��vUt�D���(��@�@�*�:��#X��|�:tK�$��-�'�6H�Е�WG�ve���PۉZ�E��h�Rz��Z6fH��[@E�p{�rXE��.d��u��آ�1�&3�I�,�	{q�������W'Y�v)o�Y�]\��<W��}D%�U5ټ��Q��z\cu
إ�Ђ�����]�{��kA�Ф�����J�G��S��zD��q�bs=)J��<5�@��"��T���¨�6׫b��������H��V=�hs=N�6ZՎ���]u�3��M���0�*�] �9�<�a3��t��U�Ѷ��;vl� �? ��e���Ք�#���^�,�3���@ Y-R�eH 1N��1���mْM3���$A~�*����Z��Y�6�m8��4w�Ƌ��V���՚t�  �- Y��@S�۳GH���1���BG���ܝ�Q'T��i��&�ZT�-�r�Q�~w=�侟=�j����ؤ�b"�2�!��M������IU��u�{וֹ[Rj��ͭ{���e@��-��'P���B�*_�m"Kh�,Pl�x ��q<<�5 ��6�S����H���v��Uw��qE;>�{rJ�ͬ9, ��y�;��J����ނ)��[�M��z�|�BM*�uOӝHf��W�Zי02�^�p���1(,���s	�-�N��,nP}AjM:��'^�@E�d�yHۅw�����^�f�j�b�ON����{��S�t?�d|U$��T�5 %;��67
̧�'\
O�g�،��[��_�����|�i� U?|�H��i�`�#�cx��0~`{��'���	T����{��Z�*Oưf�$4cX�e&C^o<����a������*j�y��Ҙ¨d��>�G�����#��Kv@P�W,�.�Ad�c�����a�^�P�("'�Ɏ�zo��AN}5M�do��9)
,��.���nX�(UH�ܥH���aw)rZ<��XbkM��`M�BĚ)�X�k�w����<��`>]'�Sl_yV��i(�I��	m-2��*�ǔ��f!�V$#$�V$N�F���a���<�ҋ`T��MP�nC��y
��бց_#pZ����v�&]P�5��P���\���P����x���5��<ȡ&�w"�O5���ԧ�z�
�v�>$��6Ncg	��]<�C^�}�%���qw�G�7�g6[T�V����Ǔ�B�&˒(-q�d�6̮�4#)#i.m�W���+C�u���(��X� ��e�ס(ydhQF	�7��
��8n*C�� �pF+3�-*�4�O��%%�Kh�D��<J��Ev?IJx�KqEh���.4�>�z�5L��j�=����.��`��=9�n6i���F���������4��9Ӏ���l�Ls{ǺB" �A!�3nw
�O����<Π�~m�!�>Bn�y&7􉛊�ȍ�o�HprK�����o���&?��`�8���v�)�1��{<�h*3��qXGz�y�[(p��Q.!�hQ��]�$�<Irm�|	�9@�x��,H���#X�f��;���̓����D<�%��?J׍�����g�:��]��JU��^�)�N���1�t8z.�g��d��$����2�Rax��\���1�$�t�[��ŧݺ1ey�]>":3jOF�x(!�@�m�P��P��o��g7I	��4����Z����>M�aROTm�6�%�����h�S	� �h��D�#L1G�L����Ƅ���z&�m h��M[�u�<���L�
4�����#x�6u��q9�-1(� ��@[K�Ѧ
���f4�ǝ������'��Ⱦͧ����:ڲ�C��ʗ3�B�-���:�n}o�d�ivkF�$n�m=�����dm��%8�hF�:E�4��S���6sP}�h� ��C�^��@h�e�	�#�B��-�l;)*4�����aΤ��dmI���+d�#b���-������m	w��ZMJO:��2r
Б9�:3Aӱ�2 ��T�~/8��ث�@)�Oʡ�{7\+��'����M:��{Q~����4�[�<v�ZV��S��$�����������u�����b�_E�zV,���~5��l����PK   �<�X��(��8  �8  /   images/02932828-f6d4-4923-89fb-67d65ebd103a.png�8!ǉPNG

   IHDR   d   �   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  8kIDATx���T����������tX�,�(HS�(c��5�ؒ�1&�3��&�F�1�?1Ѩ�1��i"(�.,�l�;���o�웶�]��|ٙw�}�s���<ߘ1cZ����&�x<��z���K\\�466JKK��=!!a��f���f�w||��{���!x�#��1��|>�< �\�r���>�v�q���͛eӦM2e����dܸq2l�0ٹs�����	��}�G�ĉ���J^y�)//��=�IIIr��'˜9s$%%E;�0ٺu��q��.�E�u�(<�]p�:,��g��:9##C$999�x�m۶Iqq���Yd��=z�̜9S���Z�߿����K����g��C9������'//���'�0s:T�-[�_�y��Jee�A<�~��f��ٳG.��2Y�~�����KlϧO�>2`� IKK3g�޽��555!�A��Ғ��w�O��Ө(P�6rݺu�t�Ґ���v��an�U�J�ٳ�lٲEv��%EEEf�u���Y����3�\\��� ���s�]�}�v�����3c�p�n�4i�2��Z���^�>r���J��/6���gAX��t�0ax�R�%J9�t�$(u���Pޚ�������_���:�\��B���w������a�\���ZxFvʆ��n6���q};Vw�%��W�^�JAAAȯ���S|���c�����#	z��!cǎ���z����iJ�=�!v�#F�xAW��M�� 7ʶ}�����o�'�|R=�P����
�%tvn1+Y������� �畕+W�"L�n�,�e���V�Q�������ؕ�;,11�E�[��r��p)�*�B	��-�N�����P�W���9~�m��N�ͼ�_�כ<���
-���?�8O���h��TU�.��w�q�lۺM�9��y�	RUY%wnO�
As��>عc��=�9����o��V`��+������J�,^ I	>y��G���e��r�7N�Q#�ˋ�?+�e%���$��		�fa(^���_���%�w����7r�5ט�7��>K�K6� H�6;D���}W^ye��gϖ;���S]q��΀Ҭʐ��������<�w���eM��*�q���Q�Ƀ�Յ���&3$>c��dű�;�H�lʢ��d᧋͹��\I���y���/iƙ��v�_�w�<5w����J��������7�IrS��Iz��́����n��{ｆ((ʶv*�W�=�c��y<�ET�3�^8X�A�W�ҴZ���:�h��47���5�����|��/���S��رn�(���o-N�#�:TD{P$��߷�rK���.�j�>S[[kvKT>j�js�bn��|<����5��Zb�(��s�D��Ǽb�]�yc�ӑyU����<+,�9cΫ�dT��?Z]ǹ�����;�4�n��V��+**233�#��i���|�8��$:�#���A %H��<T� ���Ȋ��KmE������"i�x%��@��;\�S�Ϯ�x�i�\�y� q���)��=���|�^�'i=�IF�A�OT6�����2���U��%ez��U��KL���C$C?]��MQ�G�EM��Ç������޽{�sss�a���)!��Y�Ǒ����=?p��G�e���u�1%T��Q5���]��SZ�S|2�~)���J�����LK���ee]��|��t7T
 �-�d�s7If�Qr�ٿG���mPB�{�ϲo���'�Jz��뽪*��I*<$���Ȁ����؅�����d�+wI��)2�?��l�����3Y������Œ���z�U5��a^�T��e��ߓ���"m[D��[�r�jY�R�}II�T�6��a]��t���O>	�!2����������<�4��q*�.S{dȼy��;J�/QJ������L헱��K��s�qSJFZ���`�������u�����oB�C]���RQ�.�L+�Aj���ŏ^#Ǐ��+�"#�$9)^�A�U�2��5r�_~*{t�#ξI�g�aW�W�H�����#��Z��m�+����3��"��d�jƏ�"%����ܵr��W�ލɘS�	��V����by���� /��1N�����0���s�ƍ1-��7L�q�5*;??�:%�uF�c�~���F�t�l�ʽ[d�?����)�~�̙�A��_��dמ*��'��8Z�N*W^��,zl�L��{%�N7kX�]@�ؚ�BY��������՗�nvqCc�46���3H#?�l�����e��"�}kP��Ƹ�V�;NO�d�+��;gȌ�#���IWs�ޯ�k�3S���'ɱS�ɅW>*k�H�Cg^e�+7��P9�}5V�}�,|d><�-�!!  
��+d͚5F�[�X�s�GV�p�\|Z/��w�HUu��`���x|�Kj�z��F����˟�8KN��aټ�e_g-��Y�>W�x��?#U���t����X��#�u�����o�>C�\����͑�+���#�}N�+e�[䞟-'��_��o��]R]� �����>SN��)5Mr�n�� W�����Ø
(F(EVku+FQ%2�V�u�r���l�XR*��U��g���푕,�Jk�fq��J�F��x����صߛ"���w�a���(ݱN�K>Tb|��Pb����݉�e��WL��zD���}^e�;�͑��r��ce��RIJ�Ib�W���o���
��/c
�ȅ����T&_pgTcֺoX�����m�H�ٴy�"����2u\OeK�RS�h��#E�o.uv���2E\��x�����c&��?,������
"�UVP��C9�l雗��v�Ab,ئ�n0��:i�yґ����[~��RY�M���z�{?}O������ҝ�7r#A�aR������Fe��N%��H��
�%�>?�(�����!��&+9';IW\�Aۿx_���K���{fF���U[H���2�G��f)��kŋA~Y�Ab4b;i�A ��/WeZ�N�8:b��F���)���Fz�<��&��Z�+��jw��8�i^��=UR_]*��i��ϙ ����M ��� i�	RV^�ȑ}5F{q�0��y؆�����o�x���vC�r�Ttb����j�So�[O�Yţ�L"R�qd�e���wX��7G�����;�c�9
�)��l�X��I��'����d�`w�d%Ii�#GXٰ��D'�V]S/{�5J^f�!�X���Ȗ�k���#���Ęf���� nϾ��̍�@�y�{J�^�r��CU��5;ο�@�����/��+�T�iI�Ĕ���q�All!�66�	՞�gw�1I>x�ߊ�:=��	#G6nq��p��~=�)�͖��G��[�ad�{�)QJ���I ��d�V�]�!���n�2/ZV������K/�dvq��18��6�\� �3D�y��ﭒг@R�bz�;
����	a�92HTb,̶vJ��Qr󏐵��ǞY&W\|LP�쑝���k8���T�?�}�����'�EU{q`�6N>xs������q�!�8v�@e��Ab����:o�ߒ�䌨;�Y-�AGΔyy@ޝ�Q��rQ[�<Σ�q!�3���(�W-��!3���"Db�˗/7n�~���D���G��)SU��N���~�%2lH��x�H��X}i��F+���*O@�Ϳ{M���i��g�Dod�^ϼ�N�_y��K%;;U���V�-I�NB�x#7�r۽o��M�2튋̼�1��<4���W����z�����a����Ӣ��IP���R��$�3j�s�q�ع�M��(";��w�5���1��s&ʇ�+T�M�|�=�6�䆟ɏ��K.��x饚;���o�+�z|���6K&�^�lV�k�1o�ae�)�����1�R~z�q�B���ei��?�#/,�Ȥ���80ٹ� kښ�"9���W�LQ��@������a���r������t�/��q0�]��u�WO��ɓMX�
�j����c�k�-�!~��������-?��L84K�A��(��={kdgY�d�<U�~�ʪ҃H3<<�^�g��e�A�O7���]��'d☞2����k���5����5����Hbz�Qm-X~�
�_���~ ;�����O�}p�Y�#�z�� o�U�e���s��e��s���B��!����6�*�.���a y���c.�����TVmZ!�%�ū�+}�9jȑ���� ݽ��i$e����Kzn~б螷��{����-�d�ƥ�֢�FcJ�/��3ɸ��m��H� �9Vr��s6�K�C����Stޕ�p�j�_W">�aه��)�����&\p���I��w�.��]Ch���hH��5o��o��0ZZu�f��p�sN�d�%�.��1��*蝘�Gz���~BH�ə72rɽ�:QrG��6GecD<�1gވ��y�b�~��!8q���®`G����x���!?D�TĘת�!;"rq�o�і� �yc�3os(��ɶ�����,Q�z<z=o������jYhP�����/���Ӎ�E�	~~��a)R�v���E����(q���^��� �|w`�d6R'h�[�*B�6�9������!>���3���o���  y֬Y&I�"DCT_~?��3C��_~�e�k|q-��{���>������<���Ki�A�cSe���ciA�x�bg��xꩧ��N$�p�Q��裏9�q�Fy�wė é�hb��8
C��;��c���ůApjR���7K�����p��/�ɲ���D;�7E�Q����^��J|j�7�oSF��!}����/�-/�چ��d�z%��(M���)��֔G8;էc=��c�H}S�|��"b��_r��Y�I	q��Ty|~��'5(�N>"KR������A���2���*�|��s{��Kf�7��U�9���	y\����Izr�؊Z���b|��+���D<u|�Y��,,1�fGI���N��u;k�9A�"�oR|����OvD�����+.�
�A���� ���Y�Z!ߜ��hۊ��Uef�����Se���^�j`�D�')�����^6�3��=vH�D��mv��\T/[����2@L�Щ���;����ʥN�N��}�y�N��t���Qį�V#��$^��6��������17��=L���k+�̱p��),k�:�����|y��r���ʱ�3ewY�4�[��D�����d����g�HB��7.5|�-Z-�,t2�T-���|;fJ��i�qf�r:�Z�1��}�RX��K@liu���b䎹%R]��w�V P ���c!pM��KG�׉���qeO�yڮ7d��-�+�T:�_���JaSd��dx^�<��^5�[�`��v��� �����)HX��u;k���c9A��� ����<�v,�\e��x���;K䝏ˍV��/'�9�^�Wf�a[EM�k_���%�D�n�wV���"�Kuek�(c�`��݂��sXЁ���,�3�$O�VR٨�ϰ"V��χ�~����nWM�N��0&S��y�҈�rK���ݶeo��M���f�F�o�,��Ň���O4i�6ށ7��؃0�X �6,-
�@�HeQ�Zv�a"��.�!�Peez$H�Z�ŕM��R)�j�0 ;��:/,n��}q�>٧c㾌;_u��=�g0ySii2x�`ٽk�,��m�)�ѠN5��gL�8o�*�^_Q�\H��=��A��פ��}a�HGE.���ms��	b�ymy�!x[c�X춋��Dbˬ}�D�����t��ҩ ??_vn�&K� �A�u��1��'�Hz�7��dm�]'��WF�q���c᰽c�
 E�,t�
b�]�z�!�������-Y�dI����s�1��t<QE���铝 /-��� PO�'G������w�����~wbY�<�B��p��4�����	��������5t�Eň#�����)�h4��?hA��x���Z�I���Q���F�N����ފ�#GP�H��[��t��T*�\x�&�Ǉ�E���_��C�Ô��q��E���)=Ϳ�T~���)Ƶ�9 �;i��4)S�m�����~���:*C��
� ���Ͱ+`Q�k�_z�%�e!�����,N��ɥ�^z�����T?��F����k+Je�jZ�(˸ٱ�Z� ���6��țE�dD�d�^�a,��D˲�������׾&�<�1;(4� �Un �$\�_ a�wךh��w�E슺�f��o6!QU��d�aCᮓ�6W��?�Q#���F�ފƮ���$�m�ԩ&Q���g�}V^{�5C�0�C�������8bH�	}���Mmz����V�I��ũI>��iʆ>X[a��l6Ao5 14�-J/��U[��;�m��� �J�޽{��ˍ>����4�>EV{�]���o\'9i�&"�Ya����A�a��_W;y��FTq°tc��7u���� {�Du����!�	'�`�`v�]�$p�� <���{�VY�&h�oeC�BeƤ�Fi@y���ii�.��B Mz �%�<�Z�*�P_A��A�����e��bΕ�P���������p0Z/o�ʛ[��<��kd���6Y9�,�E� w��/� 6 ��&���o��8Ot�kdA�,�Tm*sd��4)��aCh^�J5�c;'�Xe�ʭ5]j��b$U�Р��H
.{�A�zx��ϝ �bx^rH�Y�\�E��l��=tGʝ�4�U6D���I_௯,�)�g��66ICWʐ@�������3�qKM��?�|���,+V�~G�xx�	D��xB��q�/�P)o�Ժ�]��į�@Ö�u2�"��+��x;�z�+wrb�a���W\a�	���'��~��"�����J ka�s�8n���W��eJ�W��H�����yb?V�w��&��������#yJ�:��r�9Bl�8�!h�C�&|�nۮ��pH��SO=%4�a�!*A@.>({�UWy\�=�9�m1(��x+�A-�uҨ���+6ε�a/GI3�E8��8ix��O6A�-E��dO�!R4�C�����VXTѵZ��#���$^d	�N�������V�ߜ�D3f�0:5�0J�8�7��_C$W>/����T�;4Sm�����Ę�qy��p�z�if�%H�� d�'7���:�Ⱦ�f��ۘ�߻:/�P]�~�_�n|Ʊ.�&x��G���r�6Y`�jS����G�L�/5����$&����� KA��1z�"-Z�
G��;��T%J/բrt�3_a�"sW����~9�2�_����u4v����+��X�:;�o߾f�����i��v�te��5��v��`V�*\�XIZ�Wv�8�`&K��Dg<�jXRhB?4U�	�l��7���j��
l/i0�t蛪��jv��Bm���׿6��/���}�٦0�̰�o��4}��H9bB]���#z��o��b�X�P� b[F���S�e��Ϫ�C)D�<�'K�&��OV{�n�z��ޙ	����bR�
.uv��nM��I�g��|C��j�W���Թج���׿�e���v�i��B���QG%O?�t�	`���`U�$�b4͇��Ak�l��3X��d��&_������l�ߐr��#6E�Ly�G6=�N���~]�]�Kl�&�Yw��	P��!�C5��&b2ā�ݸ���y.���Ξ���,Аȟ��C,��!ҕ�Z�Y��C|n�CM��RGf��6� 	v�8���Ů�,rT[3Z���O����t�R�ԅ%�ǧB�v�DC 8qb����:a��r���,-�=�fţ1���0��`m�0��cL��d��GC(�� ��"�q���թ@�8G�?���r�uי������T/êº:�C��
���O7�%���af{���`2d @T�'�1dՃ�}��mU����O�el7ۢ�g��tY��p[���SM���|`ކ�]bm�zWc��b��`:��7�鮩�
���������m>.+�,D��hP�T��)kPA�J��v���#�EL�ú�dk�ݠ���[���v�,��+�m�(+((0JS�XY��ّ������{g���a'~Za�%���U[�=���j#kI�ț��V�1��p�WWB�l�r�{�����$�6�j����Im�u�=XS��E�z�hCMK�aSM��C��@�	lu׉���k��ӛ����x=��=jQ7 ��x:�[w�6_yp(Z1��	p4v�mj6�W�.��'O7V�b�I|q_"�'�����&>`,�i�B���iӦ���~!KȘ�-f����9�,�]���h���� ���y�xĿE˒�������w<넁8��w		t��w6��-�Ƹl�m-+���&����T�v,��]��] -�^cx��e����i4�g�ظ0��}&?����,�lMp�E�����F�W>�L�vZ��΅��.M�ˌ�n�y���Hqe��+�ND��c�>����}Yx<��ᮤP�`����m�56BC�dkjM]`�4L���� ;X�''���J\�<�JEVzs��ek�]���B���D7�K!$���3�L�O"�c��H�ƽ�lm'#q��d�*��,ͱ�!�7,����	�9pRw�pX<oر�.�}�!dH@&�w���z<�|�ȅwה�5Y�!������RS��a���\��0�.�<ei����.�/9o��K�/�$�{�P���4&x�ǂV:�!G�H{Ƣq��.!��{m�_�I!� i�x{�����n��p��`�I�t������ԟ�����$�ט�	�o��¿��`ߤ�m�����E�Ŝn$�PI�h�Ð���%)�qR�
PA(\�+�և8'�H0;���$�C�~xW!���2d.B��¶b�V !|�&E��>�������� ��XI�����C�����o����>:S�\P,q.����lA�Ӄ7��X�ZSx,�R�w�{�9I��V�Ww�#�����BXԨ�,z
v�$��w�$������]l�F1l��-D��LS�X�Dd�2'V���Ǫ�k��;k����'c��I<c�;������~�9D���5�6w��Pv &y衇̿�Xz4���<�yYT6��Wl�1�8�:t�|[92� C�ߴ�0v��Ϧ�'Ȋ���M.�g���Tn:�B��?&~ī��P/��îx����N�,`[!�݀��7��w)E����1�4P�+?2E`{q��V�k:9d�U�_[Q�dǻ�b��|-�f$�� �S�F>�Ġ����f��զdAc�˟e�� mX^��d�����.&��O����|o�Q�ρƌ-S���QwESk��n�#C'���Z2≭�0B�o� �$����k�4��x��w�I�c�G��`�;���R��-m��Ml�D��_�u���pv��:+�DY��
���"���h��:��v����������� ��u[�P��@nG�u%X�XW;�ŉ��x��fnl=_[t�=�6���l�. ��8a���Z�C�䴁g<�wSM���l#zsP΋��`�0L@*�M"�z��
2
Wms�O|����A�;���
r�P� �]���%���	V;�(^V�0L[�X���ɟ��'�$G˾�
����o6�YQ���j]�:����,蟓h�������^|e�-�}g��dD_��Ѝ�������JJ�z�}YV��\d�8��sx.��7��Ұ����~����\�gN�a�uV�W�\]n¸Ѻ_��N�|����f{M���;&��,V?�E����vc!���j7Q�=�����o�&y�^(AL��D�)�yn��R�~��=eцJY��ڴw�uB�W��Ū�� �WB㯊�%`��*~9���i��<�m�s��`S�_~�! �qd,��?��pm)V8ķ�e�9O����������:"K�_W�+��$���J0)A�+�X	QB�`�B�:*9���f�,��)��b�R����#�Mׇ�n�[��|�?��O�;��E(�`q������t�����R��g���cOd�����،Z���C6�ݽ��=TV-W[�*��}��D6;��d/Z-�*?�<0<� ����;T~yzaI���_Hn�(�nvRLA6V=����-���AHV<,���u��֭w5X_�o� ��c�1,ş��e�������'�:�EJY�J:��^��Vk�(M6�G��B�2��S"���� �2L���r8lZ~�.���~� �����w�qH>/� Ų6��|��̙3M�
q���7&?�	7�tSTyb�NrA/,�ՂgFXP�s��qJ����%��#�#�ߑT�����Gf�U�+�7Jr�	(I��%��v���!;�`�P�ЮP����?���L�ܝJ�*Lw���p iu�4bqr�DZ�-`y�[�a�õO8,���+��-��>IF��;�p'Ũ;hXoji0���x��z������`Kz����TиPy	\a�>�q(�/�����ch�A	 ��Z�D;��aD.q�ʭ����h0�!ׅ��?���^{�r���{┅�G40�l#�V�uCa����E@��� ��|�»#E4����
{��z�3�zDT�L���J2(�z���`;`��4�[*r��⻂�c���M��n��CU���8�Bk$����b^��:���z�T��[a� ��L�	�/:Б�� ��K%p��!+��HU�_��2 ��!q�����u�����!��C���i)��w�)�AI��\�3I�q�v���I�&9��h2W
�;݃�CwH�dAr=2��*$X��U`;ʡY��G�>��!������ �d~����"��[Kq���x:�Vo4)�MF�#�Q�I���=g��4+�a\���z
�J��(�tw�sw����fL�PB��G�駟JqQ���^'�a�+�Z��m����~6!��+`��+���o;;�]A(�gzp)���np�Y�29܆; �0)u#���P��kdO�Y��Y��*�b��7A��7�4�����r2����<]3cL���-�����o�����M2�n(sx�����3UgD�#A��X�$~�Z��H�:ݼ�1�0�L���	�$����.uH�)vH��5F���D9�= ٰ)� ���ļ�n1l� ��d3����߲i���47��Vt��c���pD҈�ҍU!Z�7Д̨�^'N�)*k0��`��w֔��v��N���v�!m�	�����闕�0Dj[��rt���;�=���pʑٲdcU�1\ t����-��&Y�&�3_W�+ٚ�E�(ma��6iҤ��B��
� =)@ H�0����n4��`Y�nք���&;�E�����O���Nt�O�"�.�	fB��K�`��IT2���w^0Sc���t��t��-�u��K�J�k�"�	E�g�u�>$<��Nkw֚RU��!Ć@Se�T ��^�:�N���;��|�ȁ4l�R����f�qh�x�E���1/z�V����ɼ4� �V���0�9�͜��e1���6x�(c75���cu��7E��B��9�F�H�!�$<P�jGյ��!���n���������=���Bڏ�3�˻���\[~C�u�RW�}Rp�p0;{�ؘ���i�iJ��h�!��.`�3�kk	��t������ç����������?Op�G�6�ڲ�X8�E;��S�ۉy��sQB;�� ��[�����ilj}��RR�Ȥy�����벮d����Om�\[��VbFgǒ�F��X��JQ��,"�L|�qm!x5�$�KCRRR�^�DO�T����'��r0��Ma���w�3�y��k�KQѮ�;����l3v��n�3����W_-Y�Y��ܹQ�Hj=�~�"��?�P��|�56+;K.��"s?�T�_�|��m������7�a�<l��n��D���Jq�[O����9��2���*[\ �b�)E�DxVO*ՁiJ�F�y[NN�T��Ew&�JZZ�uw-�7��ǻ�yw�;��n������ӷ��y�Y&��M����7jēE2$?_�y�9���/͑x �X[�y�̙m�Yބ��hԿoU�?���[%*�&8����Y`�w�!+����(׭7K,vɐz=�Dmm�|ec�&L��OG��A$�G�p��	�| cC�h�� ����x�� I��v|B|̱�L<)QbE��=

Z����>�r�s����}uʔ)�_}�U�k���)���AN�Ȉ�
�ڮ\�T}� ���Z�J<F�]x���|9!�r@q�/E~�4ü뮻�:]W�lYү_�Dr|6�DiP�<r��1 ��C�@S��J�B�)}��:P��ލ��ڇI7��~o��������L|^c�������<�a��(Q�Z�飼����u>��]��������q���j%H���>��?m�,��񇑛d���J�A,��:.-���uXEQm�@�䣧���i~Z����t��ȓ�L��4�o���L6M4��L=�p
�yْ%R��H��k(!�B zø���j��`���^�'e��z�=d-���%�j9<i.] �c��c��l��p��ז:p�v�9�����c��Y�<(7��"[�6\z��6oR�۲cG�Z�>b����a��ٺO��k
��L"GF�3��5k�.��8����}�ň7|���6x����{�rsH �M��U��'�b �?$d��(��\��O"{���N��'�"��߼�̂bAd�� D��o�86(�����bR�k3H���hK<0	h������f{�M����L����?_����h�����s衇>AT�7I�<�0D��曏�gK�(Rv��:CU����SSS_��� ��I�2o#��DA4��JҘ��~���7�
�A@������a�}�"�.�}B���� =B�O���l�~b�7�t��7��A�%��6���x.�3�-[��3f܊������.**���c��`^;��IЭ��^��:�c�٣ǲ�s����۷oϡg ڃ�E &q1�R�~�l��ްo�D�Õ�g�,�Y�f�����E�O�0��)�'�	�#��Bj/���XA^��:���[шY�j] ��g�x�\�E�\嘚�(q�����ڍ��T�w�����>~�a�����n�՝oP��	�:0U���"���^��ICYE��lKX�;c�>����<^[ K�=���3�!|�q���ܰ.x0Z	�x�qӥo�L�x�֭�`ڥ߻\�u~��{�9�d5����e�`��W]e
1�O�S2��P&M�l�s����:|�OԶI�{O5����ȸ�ɾ��ED���1c��{�>37����S����N,Q�fԇ��6���@�=	�S��֣U,l��`_��
?묳̃�7�Y՚�.�f��#��;��ew.fơM��Z4��-��m�b�y�7�P&Ƽ mlm��a_[�w��X����^����� G��>3�S�e=��S�>m!Da�^�ν�xFp�BR�'!�8»U��X�p�Lȃ�'uoyV%+���ʰ�`�Æh�ikYm�$n��p  �@2Id��؍n���Jq$���������ޛe��ܯ
�q����]�=Hp�柬~[�a�"c1��n$�k�FN� A6���^�wV��31��@�� '�m��9��]�| ��j��f���ժ�zN���w7����hv�U�16>p�B��&��}^o`�/0v�~�u���h8툽��� �u�嚶ȳoR�����[�B�t�uy�1ʧ����Tu��3Ϥ�؏^|�ŧ��8�t�6�f���c���o��\��+���cC
�u���=��L��e:�P�|��7����M��`��f$�8�U��� ���3�x���u�H��={v��D!�x��Ǔ ���ĩ����(!c�{T=�V��y%z���_�W�}г�}W�ࢋ.�")Ĺ�+ڃ&���UbD�E0G���� �`�灻/��_A��A�|E�n_���W�f�A�|E�n_����[�V�Ax    IEND�B`�PK   �<�XWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   �<�XK���(  �(  /   images/1042b8f9-2e87-4dd7-a644-1e53cbd80f37.png�(׉PNG

   IHDR   d   R   ��q�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  (|IDATx��]xUղ��O		B!Bh����ł���P)*�x�*łPEi
�"* E� ]Z����s����t��y�����ee���^{��Zk��ʆ>|�/�|x���ʀ��>.󱛏5ο%Bi���+|�'����Z����A6��Gh0������A�V���7i4Unn�'��4�1|l�c�n��$��tvVԧ�~�@���ΟUd��)22�֭[K?��s�ڳgOz��������D�o��o���J��N�#������o��իW����n%����5��o$�R>�Acʔ)��c�Ӂh��/)=5��v3� :�5mM3f�,�^|�E:v�X���]�6���kԦM!�ƍ�ڵkG���'�VO?��m�aY��TvR�t��[�z�H۶m�U�>���~��U>�xV��+Af���h��kגV��_C�5�*<��;�`�S3Q�Ս�b���'R��.�a�74}�4��uez֬YԼysQW��z�A o��&-\�E�;H�#�i@�F���Lb5oc5�M�o��֭��&L�N=z��aÆQ~~> ��)$HOr��#11�֮^L��مj�� ��ʄ��[,�4�C�&!��,�!?Eƍ���?���lڲeK���ر#�����W��IKK���p�]w��sߠ	�GSXc#�K�8��,!f�JU�ǧ��oﶔ��C�M�a#����>�f9��^� 0઩S��d���#?���l�wو�d2[����%%�ύᇎhь��U�6�Ez�ͷ`���'�,4������#΀V�a�}K777���+��_H��	f��.\���Xp�,ԭ[��{o��{��> &���o������s��c�����;��$wwc#�v�x��8뭷โA�~|�G}���h� KĞ�y�ѠK��U�P5�/�d0h����XV��6��\;B;vlg��8 aaa,Yf�O�>}(66V�j��;���x���{��ǇN�:E���>m�49g2���W_���S�~�(==��S��s���O?Mk֬)t
Ч��B�o���Ξ=K��>�5J�)�#����˳�����6l��;w�4A0�_��<ځ�������A����_j�j1�[g���3{ǋ�A�~D��9���Z� ��<#F��� �PS,W�LC�:mn���G�^^I��=��A�����L� &��ݺ���?o�����;�̃�*��K�.I\�����p�R#*���������w�A-[��ƍ�'�|B���;͜9S�شiS�"�^��Gy��}�Y���Ç�`d�8l޼���
���<�w�3� 7P����S�Ӡ�[� �7]�U������2��w��{s��Z^��ui��Q�����?�����#?�ԟo�~�j1�V�}��Q� D�%����W�@�x�a��5�`����~�^O���y�Y�&���#�p��U��'
"�����Ӑ!CD��B�xp3���+���ôu�V����F�Qxx8}��wԭ[�BUI�.��\�B�1yxx���ۅ(�
�S rrr�p ~U c���#Ow+3�*sTZz�O#i��ƿ�aa����^�1����1J`�6�q� �޽k;*A�> H#p��G����&����]�����Bb��S?���fb���ͷ�C��󡨨H1�x �̣�>J�z���>���]�&./�P/x.��8r�xi���؁1cƈ����rr2͞=[	�P�V�Zt��!J׮]ŭQ������>0 � l �Y��u�6������c[]Ｚ�>t��׊��9w5�{u$�N�m��L���ky��S�
�v3q����f�0�l�$k��<��Ru��%���%p�?,#=��ԩ#�:t��z�)��E�	�Ce4l�P�>�]n�w�.���p��m�&�R Tu�X���p���B��n��"�W|�|�]��Ni�����+�^\.z{4�ך��k3����q܃Lw�L%/�+���LA��%dƤa4�ݵ%>���É��9V��{ԪU+AR�-DE=z�֯_/z��733S��ڵKw���i߾}b0A����"�]�dI�AG�	&�Z���9s�3��� ���d�IK�.��PY.��w(�/ #�k��Ы�.|jy�z�/p�����^� '��ŠVB��^�)�����"�3���"Y�1�1��ʥ��z����* 95�"�s���BCCE�aG��@"��U�hݺ� _H��4�;w�سO�8Q�������/����ʒ�` �k@��dʃ���{��"O�J-�ݙݽ�A/]N�LuU�k����ڦR����y�&�9p�� @J�>}��[��+WORx��Љϱl�OL�E��Ѕ�Xz�f���W���LL���j���6�K̦�a�iƾi4h� CT$a?�y�@�#@���F��>n�xZ�*�����I���0#�[s���s>���?s/��@UQ�Z����,���	Ԃq�_�Be���_ӼwޥY�~�L��=�5L��t[�ϔ���;�|}<A!�z~�-��4�K�c�a�6̭It��e����h�N@�^�Zm`` M�4�Pe(�@�� ��	U�$��I�r�����R��X'55E����8j܀}|�r����.�h��W+&A{PRJ���F�)K�=x�c�ЫoΠ�/M*�o!Av��M�I�R��J�I=���+��%���[��K����-�m��_�/�eb,ᛷ����E}F�'�$�[�l������v�o�0�@����_�>M�>]� ���ԩ��Hl�b?@(�ָ?�EP��O?���ɓ'��ŋ+L�� �ȼy���	OP`8Dm'�1�Ƶo�dW�X&����e�#��r*���L0�w��8���/�m�iS�ґc�C��H�T��̖�d�h��3�vd���o�n�7��/� ��4@����+����@��/!;q�$� �( 8�T� "zxx�<==�9 "�4~CP	�VU����ǎ�N+�ͥ����Z���<��q���0�0����eܦdyҤO�3r{�{!��رc裏>�@��~�~�ݽ��zv�Q���Q�Ё×���3%27n\�_�)=�P�sp]�UA�A�����2G&A� 
���zO ,�)�;w�iH<+�B�ѧ� ����,�`�\��1�B��V��n��1�'|��,ں�y�5���ͦѣG1�/�_1�1����h��RTd�[�9YM���ϓ�Rbփ9��a��-;��K^��D�h@~��`��r��@E�5i�D�M��p�
�|�A�xxw�O�i�z��	�@h�--�YY c"�B�`ђ�i�ʏ�͇��[G�}<�0jQ�)٤��Ґ�'���Lp��M*Pb����z��O�2�Ll#._���HN��� �t�"=��Xڻwo��\axb;v��EI� �D��)V�ZE������8�͚5� Q�@,�<D�#G��{+��� 0"�=rg`�G}�	��k���ܸ1�3}�j�ɑO�f�B� ����' 	#�t^�ϯsl�$���Õ�N@�/�g�3C��_Ib���p�xs�"�Pg�"(N </���A�3CZT� ��O��X<���dqmO�<Y.#d����H�"����?�˒ ��� ��q( �T��;�P�
@E�&�p�q���z��*A:���mى�3,�>��������Is���
 �ڀΝ����EX ��'Ӝ-��m�8-�Q$�K��[q;*:^f�Z�х�� �V�]�At�r"{/E�檛7���� P����l,7m#��O��{N����8PS�IVYGODWۀ�ס�/?O/�X �	�)3��͡Yܞ>kۆnO���,��4i�zu)�'$��h��et-6�f����Gt�j͚>��zo%�q�"σ�u�O���NƺY�ڇ�k�"�b|�a:%F=��5�L�N�!��1�`��bұ����O6����5��,�`�Z�q�#n��D�5R`���7|�\k�6P�OH�c� ����J�KA!�Ǹ��,
��/��&m��+Fn���Ƶ,�	��NF��+W`G@�B���ͽܾE�����b:��G���ׯn��u�ۗӔ�k�8�icj�6�BZFPj���L��B�l�X�>�&��qO��؅��Jۮ�q.2�٭Ζ�>α��v*)�VI0�*A��1`<Vk�فrgj��{�r�F|����~tl�~
�W�4ZGpeb]m/0R�>R��]uj'�B#�f��f�aE�ʥ���Tw*U	�o�VEER F��}"Ƞ�F�)�bbdf�Q�.aԥC(<r�Ծ��.\�8�2�,)��2w�Z�9ر��l6�ߏ�N�1q
��b�s�
d��h�6���}�p>�T�?���_�<����
�j4�龻�QRJ��߯��
��J��/��A�V&`�����#��E�d��~˖-�Z��E�.嶗W-،�!��ߛ4i*}��=(4�-_��D����C	��jIGD��*#Y	>@j��5�
�51"0��Zvz�z	r���C���d58�� �`�FJ����۵��<R�J[�m䤐�G���O?�DC�Jz�H����o��t�x
m��2��K � K[�n��N#%+����t�¾O�9G�� ъ�wM!�L�炴�rO��(�c,6C�%��4wJJ-��Ĳ�`�%tu|b:��<J�i-#Ճ̆:x�ef[Ġ�5�Kލ|i�敔�G�9Y��r]C[� ܷ&��r	r��:z�<5k&`�5��:_
m�]�, w7:~>��|���t�_ ��Ӡ�(�邖�Һ�h��=ɨM�Q�����D��e���_v��Ke��߿�v��N"؋ ���͛����W���`6�G��eɲU�0�*V߹���Nm�4�<A�����&n��{��1.i���Ȣ��"��Z������	�:��l�;�����?��p}�f���eA����E�G�#y�:�B9B��lZ��6���S�
@j�{nu��^8�J�a6�v���!����,���Z5z�xY�9��"���m@�'Ӻ�eo,� �_5j�O��#�PX����'��_~�ܗS�0[�jޖn��_���H{m��V����+q7�¼� ?��lv]1��'��V��3Kp'�\���}�� *:|2���E���rK�Z������N��+.qzZK��.]I�:���^m�\��]�f�%KD?�j{��Zu�%
o¢�˶=��y��M�BQ ���`����6��e���
�Vk(%9��әT枴nS�kJ$������n#A���Iz�Y�N���gCm+�8&`<iƌ�@��ŋ�O �y� �dk[͠�s�K>��6Pp�ze�-� ��Fz`Pw�!a�o���L�$3v�l�Q�J�ϮQ�?p���̕t5�˂�h�~X���̾%	�Դ,�!�/]��N�]:�̗
MW(�.������ykd�
V�#�R(���u���?�諯)�o�1����\6�P�i*�$)���RR��+q���E!�qw&�pd�8�� �;R`.!a)���<�@:��8�Pu}CO��F��&O�^Vԯ-��Ҳ��^G�	��(8��l�/V
�T��e9ԧ�t��B���E/O*�aÐ�ܚ]�4�=�M���,�n��<3v؏rs2�Ա��a����w:w!�0��䟀,eZ�:���F�&&�:�%+k����&%���{�x+����R��H��Y��_k��Q@@��7Q����T/o_
jB��t��4�:%=�D:��1Ee!��/Y<���~]�l5Ġ0N��pג��W�}K�CV}�C�nI����JZ��j	0�>_A���B��� G��<C�~2 ����GU3�7.��GǑ�Wm��/K�7PZ���^K.�oɑ:G�{��*rө�;w*Q̀ ��۷��\qXX�Ϊ{�` Ż��ɧw}KS�N�\VM񲰚���$����̾���ի�c������z*�����?i��C$*{ȱF������t�ԙ�+�N�(��=�N��v��O�>�nmu��Y�`�{۶m�XX�
���5qBE4B��.�	�r����ceَC����h�hQ��B�ۄPߞ�����^VAZ�&Z��}z������B.���|������iԨ�+�ǎKW�^��|z����bt4-X0�Ə� E	���a"�=s�>�`1��Ҕb;u�lŋ�	�/&��?~\�IiP!����5 �ޓ":���Gi��?R������ɦ�����
nN�}O6K��D\h6H8���b�D%+"akmi��RΫm9�l�wM�y��G8T����d�?���u����X�r��+msS����dbψ���݀}�Ӕ��Gu|��n�^�������<j�燩���9A�\��X�e�~Hy$���"�����vE�����yw>����\�aw]]�!�Z��l@��JG�y�c�t��e�����{���>�b�	2d�T�=z�\[�z�J-�@l�%��xq-������/V����tѶ��ߒ��v�����l%�=Fw�3))9���$-Y��Z���ɦ�<�tAF6���l���(�E�o,��h��1;q�z�(���}��6���j1	!���J�ö�T�+=���Ӫ���хr
�Myt����C>��Ξ���I�^ڹ���9i�6�9�*�_8���"���ɭ�N&����̢e7�￻�I��kD{������o����O�=]�����R��ftp�Wd�ϔ-��+5HEy�����:�E��Bi��)R}бS�7�mJJ8O��l����+1�U6���"�#C,�"G�U�p|��.�]�M�i��Pbr����Iܶr{*����$k;u����%\9Mi�ژ6�JI͒��鳗���"`w�v�iU|�C��P�M3SJR���k���R��ܹ��
dG ;1v-Y����u~~~r���Jm.w�biP!�@��ň��b��@����H��UŚ-�Z�,�V�]�����꜋���Ħޯ������Jn���ca�����bYڴ���ma�����{b��Ƒ�Sd0!Ω����<��!ԡmJHʠ}�)���
d�޿�ԙ���k6lC
��\�O-�nzvmAV.�5��n�my����2ғ����,Q�(OŶ�O_ھ�JJ��\V��a��q�X˖�J���bcα��ei�),t���D�.�����}m�����@z������y��k�//�Av�����rr�{�n?L5rr
�]���Y��a_$�2,6-śԴc�^����;9]-^dYI΃G"���k��昖��ʧ�m���gNҁ�D]��R���S�:wh&���_�����?�,�o1�'��MH*Y2������ϫ�J���9n�#G�3!�FT�S�r0V�d���~IjAJ+�W�R|e��@y�������`��'ٍ��6�SF|}�ng�l6�c�=/� %�rQ��P�U��0�lEq�9�V�ݻ�Th@�E�po�*S-�F��B�T1�~C�gGmL����o�7C�C�ŪZ��rT �K�.�.ٴiS��4����ϲ+R���V�\����R�܄ �w�T����!����Fӻx)U�ր��fp(�? )�$��x
U�p/T?Ey@���T��H����|����hIP.AU�����i���P2����駟RU �bw���G�Hp/vF���ʨL|!��rM���k�]�pA���yX=��Zպ'�G��ؐ��[���}\��U*dCP��-��m۷s�m�k�b(..��
  �t:�&Z,6ڹs�����-,��Խ� �����N0=�(;(�������!Ծ}��@UmJ{@J0^ԏDU�#G���=S�{U� � e�{~N��t
��b�MF]K�{�L��m��Q���Y0�u���R��P�Z%�{���m;˂�+גh���왔�����MJ���D�k�}�qYt��n7BA~�A�G�!������ҙ�U�FR/k��Bw�d�E���_~�Ev؎|�K���⳩a�]�I��@����MK5ُ��l)��ku��kD+V�Z�(���U�J�X���nڠ��u���-f��蘑wP׎aH;�rZ���ݽ-�dK�z���~��(��?6zJ	��-yulJ�~'�Whވ�}�.!"�=�C	����ۆ҇�n-�� n����шWfOV�Uu:�oF�~<@�m��H_ج��U���ff4dF�j�׻G�賟�艢E�ʂ
/2bh_l��������&�����^�[u?u��컮/�5m@��삨�R���$������������9w��@�vj��d�HH�����F��8׽C��%+�sr>���ɧ��n:����e+��^�vi?�{�9 �Ȟ�{]�^���9 �B,���ha��<F".//�I~�Z��=�%�S��<v\�@��-�<���E���b8Ƹ����q�v>:V��Z	���[����i�F���u�?;�չ�2��3�&k5��sڭ�왞n+ڵiR� �X�Ks8���j�Ie'7���߱~��#�6�_(%(Q޼!\�ϼ�t��ycD4����q���TQ��pD˸��9�/܌���ԨU)����`������0y�c�ɒ�ձT��l��c_�ws%H'�J��f.4Z�	A��V�L�6������Jߛ~#Ad����(��̙E:��.b�G��n�b��-����H]Xm���\w�&�� ��蟞�o�'#�i$)ɗF������@�Ǭ��E���� ���+`��F�����]�.��&�U�"��r���=���1(Z��`c�Z�z�ծ��������g�2��T����������!�(�'j��bQ����=pO7+$���4���{C�5�Z�s��aO�\6�޵<PDx�1.�a��q	iPA����A��0����0�0�����_�I������=--��ݷuwmOO��IxNa\�{p\0�jL҂�@�|�Fk5���x�k�c���,����B2��x������Ú�����W��o�ဆ��0��� � �qoY^O�w:��E$���v���/��fx�W8p��V�fb4`n���P���c��cQE�o�yL��1�~¢ޕ9�Jà:������y�u=�]<����k���27~����H���0� �E��>=Zu�{�䱯�[���Y�1w�g��v�vTw�ُ��[n^~77�C(e��P����KҐq���֎��8z����w�� �� A �~��L*�+ۇ���:�������w�Yy�t�9b 7�������ᚮ\�Mvi�t2R
���`�;ѱi��n�i��%=� �Ut���X%��!r�
h�փ��=�JX�wu7�B���f��o�� �m��ȭ�4��`�Z7���S{VVQ}�j�xj�k`�}��x�p$}��+�A|yr9? Y E����Xf@}_���_���%�����ԬI ���eAx��f��Mg#c(��æ`�����-~��'$��s�ЁAJ,��賭�nץ� _��[��5����-�q���D]�+�{R ��T(�ǆ'���K�
���� �N>���P���9*x�� �2��@�҈P��e��8`��
�/!p� �;�w6�^���A���8�g�bK#� d:Q�ky�)!��D*�@��oUrG�P2��/�T}����H�`j��ue���2��"�T)�����B*�HV"{�t}uavp/Qqa��g@o���H}�/��@"�	��G�ߪ|� ���1��G6����J�A0�_�8 0J���Y�2�HT�z62��L�e��=�#���������&@�W�W�Mx)�7#��tU�{"͍I  �E��$�}*�0 �w+�3G`7�__@�F��j�`��C�|��:9>Z����;@Ea U�@LaFdq�<�� �:0��)�+pP��2ҘL�کL�&\UI �`5�1���R����|A�jj��?���B����M�OV���a��&�T/ s�J}un� B]����
7Jf+� ������V�&���x�@�dR    IEND�B`�PK   �<�XR�\"# � /   images/16f29068-8fa2-43fd-94bb-aa3b1aab738c.png�|eXU���B��Hl�"���H��Ҩ("ݢ4H7X` ()ݠ�ԢA�.�\�t�4��Xx��>��o���9<g;Y�9���1Ƙ��/+AJ|����J޽� �9����m{�\�y����-Iţ��zT�5����]5���&�0VT��ԶwTm,lt��1���6�u-��-����`0�0��o*:���l��b���/������q���<?J|��yV]"l�G��ׇ��?�8\���ʹ�>��N��p�+�{�+�=�������_�~����R�sK��0hb$��������!]�\��|1�����q���q�.I?�_�~�L𿯕�pZ��E��G���;f������!
�|���X|��`y�<"����F>�������j��Tv�q���FD�=t�{�\˸U-��k�V�NF+p��G�ڗ�+]�(Ǵ�=���}%��|�tB��I
~9O��K�\Nc�u�������}�������\O�D�[��oԖ�����
����}Hs�ş��r��8�\W�4�DUTT�$�ns�nľjܑ�����{��b�i�:0g?�cձ<V?f_�fr0C�U��q�+Q\�~;
�c�#"]�%�[��6�N5�]���^֥2��e�(�%�w����{:�{0��՟b��X�Jh���v���Tj:"�pn�G�=�`�?h����M5��AÇ�a��.�ka���i�_}����4�*���硗y�%�ڹ�m�e�T���S�99<�cS�0+̼Pre�Q��r�:�:��V��R��\�~�i�`�KE��Zƙ�t�^d�n<����9�﫩�����x��Z��?u���.q�J�<��O�C��~0����1���vk���I�q(Yih)`7ߑ���S��cf���{�/�n����Ɇ;� ŋ�������M[����ϲ��r�Vʨ�4b���9`x�G�>|8bʹ/�8·Vp�����T�]���G�]��VK����rT�:,������m�i�;t�(q^k}K��DZ�os��X#|���c�fL���YF�;�,�rg�DN�d���zz�	�����_t����?6����x���kf����^�r���oTЇ~Vj[^��&2X���������I��2��!JJ~��gW�v���v�3�Jì,���y��%�K�g�&)�����X�R�o��� H���)�@��E�E�8�~��HKZ���*萞�����l49�!��yRN(F-�`�Sfjj��{��=�U��|-?��ϼ���րo�.�m�|�1^��r�4kf������t��7�\�9~��)WY�j�(�l��1�����w����;�q �`�q9�Sz̤/.>~��u�FX@�w�QJ�$>t��7��".˄�ّ:��I���1�m_��.}s�QS[ے�_����.�U%��QO��7��#��.Z�~]�͐�Z��_�^*F�g�;��O2Z����UWDE-��֎���O��|�Jj��2��}[&�ʩ1?T�?�ՠ�E�}�'�\Ŕ�m���5J���4�6�xJJy��]��z���A߾��uPq:'�(��f{�Q����n�������j���&-(���w�{��VJR�YH\��CE'��q�#�%ڲ�>t�;V���4�c<<N~)�bґ�DLJ����Vo�M�̼O�U1͜y7Z�k�f����	��}5�{���t�>Œa1X��h�VQ������h"�`m�/��ā�yb������]���Q���8���V#.�Xz�Y�i�y�~�*�`��f>���B[9�(뇰��{A�M����P���gy\N��&I1���2�~�R�?Rv��.�λ�jZ��C8u����lK�E#�!������3���D��sɁ,*̬�h7����젦u���ʥ� ��?��a�����]�g�N2ʶ�l�����6�fp:�Q�:Uc02���p���j���"��������ǔ�n�|���v����o����s���+׮u/_p�o3�#Ͱ��D{O+�������^���]?�P�Lll��K���z���Z%��3a�	��&��v<�)x�"b�԰�-��*���%Ǭ�*�y&J<�z�6�������qj��sv�B����P^� ff��tB���122�7�A�]��=���t���k�`�3MCIK뉔��]��� 6 �f���KHH�̃�����X�S!�K����]{�UHZ���c�D�b���`��<�mH�0 m�֡b:���U���3�K�$������_�8Ե_��1�@�8D�V5''�ߙ�e
m1n�}�����ҧ�����w�+���9ߙ�xո�0�����ry����l�B}0Gp�T���P�t�~7:�����S�6mfҰ� A��c��������"��&���55S���'�"G�f��M;S�mms���0����Gp' ���g8{Rղ���o5G
�t0����?*�G��_8�fa��W�ڟ���B��`8���}������k$�Q�A������ܩ�$n<|���
l���3�R�K�.�@:a���%�F����n�9��75YZZJ/u�J6�,�PTS3�ō�����L���з�ii�l_*���Ƭy&��h�d���I����<�נ�jwo�[H�D8�;�~��K&JD�Ν;R���j�F.���x��F��s�>�N3+)*�j~o��x=L�Կ$�C�\]�殜\�m�������z�I�y���!�֗�0�س��^��@��F����
����]�2���܃��r=>Rq����̡�������C�=9�g���<h0,��j6�_���ryZh�T����l��H���jzw3)m0���cR�^�
�#�x���?(��c0^(9#�V�����P�&�������9����.�^|#dvk�G;|�����?,��r��K���$�X��͸��ı�i�~I�7n�3:3�]��~��[�áQ\�u�p�}O�|�ΝW�!qk3]a~�?~�<���#q��$�.<�D0�����T�繞�FK�*� +�|�J"��o�(�H=1DLIE�~�1��:�P�l��+�[��8p��T���h����G�W�3^4�#x��YS�Ы�����[k�%t��Al��iOVbi孟>�G�;�Ȏ�z�C��2���͉�.pv�����vS��s�.���Zmsl�.�g@e~���oQ#y�B��4��C;��D*�(�E���!$d�E�?IgBogci�5�]��鵑�V#U!AS�#��J�#�����J�ZԐ$m4A-�@A�-�X�k/�ˉ��<v2�q��� y=M��c� wp������DUs�F�O���NLL�wgϣ�o`U-�/y��{s�qz�}�%.�_v
E�7h�&s�B��J~���A׸c'/Or�oދ�nmmͱ�SG��4�^4�@Q�}Q8�z.E9���ʥ�i��:u���ԵI�>ϓ^��!Q*Ϙ���{e[��$/�w@� G����F�����J�'���(/�6T�>��75� ��S���M�BР��@RY����U��{io�B�ܽ`v�'���k&
�.��q�&У�"�&'ZA���
::s)��=��/�#�(�c�C%[�kE�mW	�����˒�~�/Z�����Pq�g�u=�A�>�1ϘXr���9MD�:�(*C��`?��xQ"H��cAAAVOC6U=W
�*C==����?�ܵ�K�ҹ��М���쑯}s`�߿�r(��@AW7Fܗ�9@,�(�X��1=��0����sXSpQ��G~��zi���Ʉ]����T�E��'PY]�N��(ϵ�u��mU-�˪en���h�`N#�����������˗5S��||�7o���K�X��ӣ�$�@aqw�S7\D�f�>Jd.3/��j���2����hJr���J�N��k,�%T�)i�]��~v�-T�ɏ�'��[ ?H��g��o������:M@M�|�y=!�J��x��T��3�Q6��p�۵��&�k���&�N`!��]�b'`=��)�(+H����}�������Yp��A���|E��;'	��
߆7.�m*�X�{[��[/ʞ?ޔ�-����"Ք�y/D�<U^=�_���.2�N�5��W������EK�s&!!���ᷯ_߿{�f�hr���&%%ErmrJ���|��5�>%6����>�y�s�PO?m��P4��/h�f&�]�n�p.^!��� H綡`����ի9P8Ǒ�;���E�jv�{`�L�Z��K*��J
�����m��.�C��l���R2J��n��<<���2�zd���:�(�>��#H@�q�ę�B�EWxxV�	�-9*ji=�������fm߶�JX|�С��{��xn�.e=��.�	7�q�Մ��qbe�����䅯$�r�p���jߙ��f6���4@���}�N�,�����*�������ՓѪvЭ�� HH���L�3��\�|꧑��ngj��AK �Sm�TUNc�ɀ̭�8_i�C�$b�(9:�T��Vյ�HW���յ��9�/rX0 O�H���yii�ظ89�-���� ]*��S�
�Et��r��NNuuu�;V��Н��T��:`K�D7��'�N��_af�����������$���i`Ev��}O��J��U���M�z�8�|�R+������?�`�Tmb����y���O��y"�P@���=���q�^kW����ȭ����Z{3-�!`l�� 6��0
���ϾH���Ť%�r��EZ���L��I�SK�G�~Q��P~i+�jq��<F��m�Ӓ���.���n}�����:k�w��K��h���9A$XYYY�@�üt� �� �7u�-e�f�V�	f|uVRR:�sS��$瀼i���YT�ǎ#�s�i~�F�Wto�E8�/aw�*åKW�����s>�̱�A*��`H���M5��iE�vV�˟��U]N�x��Kn���W�ѣ�_�~9>4?7^IHL��311��Xn#���Ҋ�e�!ۑ>�ټ�|U�"zs����&G|E;�sD3F:ޚ��Z�\�㷎�N�
s[/�2��nٖ��q/	b�HLMM=�t�%N"�3�� 
��7��W'!�E4��\��:-%`�vM��ׯu55�G䍍��ы�nť�6L��W#YO�8p*!>ŵ��i)��a��J)ʐ�/}IO�_U2!"����q5+�f���n&�4�@�l�����fuBt�g�Xd*̢����W�����~x�(x'�_��)�le{#�W,a�e"��P1�>q�i�E�i����C�~�CCC�����T�~ǯ׈�\�rWRRRJRR�����ve��<�����H ���ji���*q�m;����X8��营!36�磣z�������s�����an�9�5K�����,R��|�ʞ��3ok�@Ґ�6��Ӽo�@l���].�d�V��1�'Ca}��gD�_�m=�]��-v�����}Sg�p�։'��䂫GZ`�@�Eh�,o �i�	2�a���/O�/�I���*8S�_.���b֚��J�s,q�����?9�=S3fm������40@?��	�e'|K�}�w� q���OM#KF�[k[�)9�S�QBw�W��3>}Dp�j����g�������Af��T��?PP�(�3-�dOav�Խ""�����-�H�����6��������I����h@}+_D�1<5/����e����Z]N!�.�/0i�N��u��I��L��!|vQ�}o%��3��_�E	�I&`���=0�hɒ��"�"���M'={�ғw�~[	YPdd:�B�x�DC��F�ְ��Iroޓ��8�� /��
�
N��0�)@.��^	@����Ȕg:�:PW�z��>od�k't�i\G��:P⢤���N�"�֡�k7����Ғ���ƻ�#8�9װ��)r"��	��<��Q���y�J:�c6X�%�E&��t���+���,f�ܷ�܀^�W�h~�׊vMd�O�Ҧ�=�L�dg��r��TI\��^�����\�^HKރ#���k�#�5n�/��J2��[��K�(ݒ""��y�&�a�I�}{LG����ߚ����;��:ۓ-SK�z�h��)�w���t�Q�)��"{��\�rC��M��`��ЕJ����,���l칡|Mv��6��������߿����ݻ�����%�_YE>)<i�hru��@C���9���W�˗/�,,m*:O+_\>1F�)~��J�h��� z�1�����������R�r�zp�t��DS�Lmc]]+����f�'��H�YBJ6�JGA��W#k��gG6�	m�B��<;Ƽ~����w{}�[d�LG�C��\�]�������"�E��A��G��_?Uu��^�	���D�u���0�V��eJ(�� !�:[����0�G��o��QIЌ{h��vGǐ!L�D��m2����!�~,����R���[(?Em�t�ҍ[����a�::��g���YT�����'�?}�B��O�r���8{H��K{�:�ŋb [�ȶ�v�- p�����7Z	����ʆ�����;z�;e� ��"��{r�Y�j=-���rZ�w��	II)`���h����%'WY��u$ܣ���7�J�T�J9!�g�9Xb#[es�t���d����A�<��FO��U Q{�4�_��^�[}��}7aL�c*O�\��w�w����8IFV��W�жA��m=�˔�o^=��G�>;,��6�wJ���FC��c�@�6קyRY|�!:�
��/�{���X��l>���Gx��X"E������Q�+.6r(q~�L�Yf���55����s�l
Kz�-�W����E�Cq0���$b`�P�=���!ܚ�<��1C��g���8p�Z� ���@�[��2�o߽k+vZ�����߰
�fҖ(���=61�"�%�Z�Ձ���qE,h�Zj�$jz��(�t��n���lR\�"�'�����klT���-X&�I�����77gg�OAye5�<����t��%�kW����͏អ���T�~�V�|�x��a� �Z?G�|mH-��&)P�~E�vvs�J`�U��>����!��"ӡ�g���B�C�]]������R��/����vR-�v�y�,��7ڀɰY��G�5q�='%-̓�\�!� "l��SV��9JL�@Y���C8����?gx�>x�P?~<Sz7J�=���LD�1F�>�R���2h�|"u����,��2�A�SϷ�aB�����������CY3/���6��`�@FG������'���9�C������XQII_j t%�GI;~a �rJ��d033K�N�a3�mld�����IMe}O+�=�;�p	�- ��7ys/1"�6f�E�g?���׺T&��\qo�P5�K�~LK�� $��en%Lj��d�qQ����hT�jd4|�,ʟ����5j�����	�o�,מk���Mf0����K\�2�8�%��Y�AvO@H�`du<uU���Tp%�k �"�~�]&@��z`+���x�J<�L�(��Bq!O���Wh�`v��@F6� ��P��v ����㜖^��e[�.��xz"8s��OU����s��
�~R��:�ߜdL�̞���삁U�ˀ�09�y��x�kp���e�Iz6�Ǐ�0
�A��^)0��ǎ}-$c�QN��x����#���� ����HA��=�B@x�_ݴ �J98D�f��p�L�Y�'>q�m��HTw��Nh+��ŋ2����������ڧ��!��X1��lmk�5i��'D�yd~�,X?����
��zv���&[��h�z��Qqy`~�+��5d=�Y�$Y�ǟ�Y(�Yt�? ��V~��O��g�ނ������s�v��H��)�9y��я����V�d;ʻ�A`�FO�x_���P�7w���7����I��
�������dK��������>�w2꫷!��3C�!�{��&׳y��;t��a#gh���d��� �T�
T�Ϋ���Vd���U�v�`��M���8�Oc�e�0���9F��H��~���p�|���_$ �cN\�t��u�MT��_,8\fa�"�h�3�M�)�= ��[��`RC�����,����FJ0�M���壶q����6�4�8:�[[[�c-t�e}��ҫ٪@sz��ؒ����k�«Sm�`�ύ����>�^f�u���{������J��q�0��������ߪ���I���f����G�y�=�iU V�uݰ�{phO��ޠn�P�;米�����ʨ����%U�+a��
jHk~:UI���P�I¦]��\���>H3�Q���-�G���k^��4�zpR�l���,��ϿM�C�j_˾G������1�e7�ͥ��^8yA�}w��2v���1��B�j�x��� �n�2W���`���	��w3���G�C@@r�h�l�2��<�_P�X��qo�#�5����-�b��	�Ǐ�-9Jמu+.��z��|Q�S���Dә�z�(��l:��e`8�H�_aJ��� �YX���͛dBBj���-J7�=�ՓR���G�gB3VZ$���7^��F�"Ga�O�ѥ���l?|��q����	>�=6:��14����g����X�Jݰ���Fý��oN&��eT���"���<����T��^������P�% <�o}}�2u+�!g�%X��L�Q˭
OR��%L��D���/ᖡ� ���Ǿ!A�!��]��.&����8C��"h� 4��K5ݛ����oy�ud�"L��&��b<XZ�I�(�3n���L��)z~ j��4�$�c0 53��M3���P���������P�:uJ��E���ϟ᳌S	w٠8`�g�Duc�jZD�����̱)@݅�޲��N'ğ!�.qFҜճ1C���B�
E��`���7翼��\��_���~y�?c���[��#G�(����$�RS3mI���@7�`^ �������t)��̯�g��_�-pJ�����b%�~�C�A;H�v�1��<<ɾ�t*��0c�],Im�v�c�Ev�C���rssMMM�oȿ��B�p�g��F�����N��� ;²� ��o�+\��w�_�4���?���3���}���w��%v������ٷ8��t,W��4-������ū������L}��(L�}�w�O�kega/�����Yq��DD�8�IFY$=(-*�HB�+ڡtH��.wP����hjbR73=-���A���I�%%EPQE�� "��Okjɱ�S�u���G�����P��mY�y���R��'�S�ґÇ+���>EGG���8AGC3k]��}N����}0�(�;̍Am\E�Ӏχ�?{�'��Wr����2]jz����Bv\a�V����df.ܶ��v���������>n�ޅѫ�e`�61_3}���ZhP�X+:�U����{��x��4�9,S�i��%�}�E��?�:9���#{w��m���w�h]b$~/�1hdmaP%2�cG͹�]�����W���K���FQǔ�[��ڴ�;��t��0n�^���q��X������?�����ѝ���F�o U�\��@#�L�.��M2��ȼ��sn�z���+ܱI]}�o8�Ӕ��P_��n�0����qs�%;��c~מ�[y��c��d�i��\�Jܾ�s��uw�}}l_H�\�d�t�Ѓ�'��W9C;��f����3���le��L2�,� ��;���ԧ�D�C�Â��2�x���w;2��d�[{��,F�����;���ܼ�yw�nTέ4�,`5!�^��Spp������)�� �B�t�@14�Mӡ�!H������-$s;D���b��ݷ:`�������,�F��m����{��X�^���� v�Xv���w�ky�穋�R))*��,��� ?J�4p7_ad���3�U���o�B���M��Oה�� ۽o�+��V�(vٷ��-A��_##e��^�Tժ� (����>IKN�R���������!Ӡ1�_���ST�c-���?΃�c�*Y����\Ft���c�o�!F�*�#.]�G:	�тদ��. ����6��(���n��1����wo��n�����%&%������z�U����ӮÔ�� l�
����A�cA�����stt���Y7g����b��cs���Q���֡��w��W8j�޲�.x�2�l��ژx��eMII��ty�+)��<������� ����uzxj�ӥJ�(�.�W�������v{�7���F�a�E&�"B���,%�_�~}"���/��8�mf�u�{:�ï���/��d�)����)����/�����w����Ą\�5��Էo��A\tq,X�4�39����������J��X<�V�Б�=W���PX�Aו��n�τ��Lw���ef�
��ʆ�Ye�T�-//��φzROqqz���!l���P�7�ͱ\���<�~���|��MZ���Z�I��U�ߙMK� ��7�tf9�D�PQQ��F�y5���5p�7�e	L���VŬ;s�F҆�1���D�6����J}@�%�(?2^΋�vjXpрN&�f��݁?6���3G;��j����
ZA	f�:1f]�������o5:v�����Ԕ��5;�����Ҡ����o��ٜB��+W�|�$�u���/e�U�%z��������uy�  @V�C��C�!�:���"���>���-JM5���LS�P��\����olYZ�j|<���%:�VH)���~ѿq�m���U%�>��4��9�W9
�۳�Y=g�y�>q9�4^_�FD����\�͛ϴ��.����P���r_c%'	Z�CסTY="/))9�4R}�p��>@�h�+c?)������q0����4���5ݻ�����*b�v�,��٪�ie.�B��+�3�vA�.�9.�S,c����z�������傘�1�߼ys�R�����������8w���K@k��>��������*[�0�)z�t�Dlssen(S�[�f(��q���L�H�'�jZ�Ipo?!��"�Uo��E.JĤ//:������z��T���#͑.��~wC��S�+KY]]=!..nm��|WN.g޵�P�\��E��r	�ݭ7Ër`��f���j4��[]̸͓�`Q����(�/p钞��٬p({J��٤�/h�me�Q�q1/u�`Ӌ��r��Z�jkkѱ� v-t��K!����&ehR\���
t�g]φ?�)S~�b�4��rɰ�9���փ��s
�Ωc�q����/����S*���u�ʕ׏q�bK�l֚>��7M�y&(ݕ�D�3C����	���6������;3t���pD�=�,D�:SH��������ѣG���v�<NL�
ڋ�Uh�,���KIY9��iWz 5�t�#�-;�|Ok��?��>��(�r/>op\B��?{�<��{��0�в������}%-��]�v3o��_, v�l�	���p������|y��]Ni9�z�??�hҕ��I�j�N@pp��놯��>7�(ZU���L?�G�#��m�f��A-]����N�`Q�3H�=�:��;�4��>8f����99��^���,���� ߃a�P�N@(j6\��8IC�V�t������e�6�fZd�	P0x��$o��'mT`����\���GF!캅2ڔ�;D,aV�cll����ԗ��E$3�E�G�^����D���TR0?+3�>[����[��פ�0[�͘yO�����'իX'��חB�ļl�^!�2/���]��O��δɉ�am�Z/U͕��
�X蟮�t�����S�/����3����qp�FP�����z�c]``^~ND���@~IIA�[^��P���� Ad��5�k<]����,��)@}��z��	����10e�9Œ���� &���/ {ĝ��X&'�� ڍrv�DO����nՔ�t�����;��� ����g��l�p��ú��j�.@���DS���0�I/ "�����1����ƺ(ZI���mc8~h7���A���!�"��r�����&�����y��H��b��V���L�^��5���.1�l*^�E�7��NC��z{����������uttD�ʲ�3������+;<w�f޿�@���
�d:�!8���F:��'z�������瑂(���@�S%���*زO�C/ȫ�u�����7���-x�;(�⪙!��|O+b0?�@�߾{'S+u�^>�7W6F|g@ yX��e�y*���g�(~����U�VR�0�ֶ�DS�\��r���k�dŭ ���J����3���JBCϤ��%��tN�%ɕ���P�WVW��{@��-|�E�KA�6Ʌo���a�C�Б���� W�����y��}YY(>�B������ֶ��ly{��-�1%����e��EkP�鎔`<�tI*�/�t�WfTc��e!n�@Nf�n.G�wөFB�pD9O��Z���Y�n����1��=I�v洶xD�o���c�
-%� �v�����p$~�<ɕ�]. >n��@����$ڞQQS������-��M�ݓ�����G���G�/|~m�dY�Ul'�%m/�3��P����g�^����e��������A�p��Z���fҷ~K\�[��t)Qi����1Y�Jq�!\��jjЋ\��j=��R�ٹО���,����t�^��O��S�G��	7�=�e/ѝo�knk):� B���<��ě�������;ZZ�a(�mp��;;;���MZ	D"���Z�911Q�H��G�T�u�8����$kZ~;�%eR���C�<�w� ��U���C+��+�I��6����}��'%9�W������#�^�|�$	��r�'$T~�E�b�n���g9�B��1k�Κ��@gy�ؠ��"��������^��4l7��OL���W,"��J]7?�7����-�&|�q�nZq�;��CЙADD�	��ݻ?e��{�^�g{l:��M�v����/���SNU�z2X�4j��h�$~tt�uI
�>g0�Y�cR�Esy}� �gڟy���\%�C����;2�@ȱaBNY�ߏ�R֍,���ݻ�A���ж=�"��\`Ɣ���� �M������Q�m�/a�U!�6D
k<x� G�w��+p�o��뛛�U��:�,���ղ�&�);�D�7ߠ�8n���(�'G r�d�����u�2XpV���������f�^g�Z�=o
��g���(�	}D���*�9o��į��͑��]i�,<<�7wM��P.|B��0���Z�i�7�A��EcQ��z���z�/�"�TR�xAD��{���P�������޳�w�^�I�q7�	B3T�_9��W���#U���`��*�?[�Q�B��H�L�󭬷�g��6
ϋy�@���:+R�3�iݦ���d��;e�^�LCVMY��龿'!( p�s��Y
�"��^&�W05�Smǯ�������<�|{2\�0͞<�q�6(M�믗������m��GO2�z�k\�|���R�kJ���^4���L�6�_nm9�噅���nT��%R��m��_�_(^�t횲`��[翤��+��V[�v�?[gg��hN����*���� U�o޼�&� p����1g2���� ����j�C�+�����x�1��~��붒�����6_>�ݮ ���:V��M �,�	Y�NH^�o�9s��LЀڢ�R�uyy�G�>��� {�� 2�~�����B@/!��Ͳ}�N�����C:l����?e_T�f�}�őڂ�H� Бg��њ�Wmƥ���4Rv���Z�7{��sB�d��5�u����0����$QDz3�ٗ.^�T��:U�c�����f���|��[��?/Vc��;���*W��\�5hǫF��-�x9۰9hu�v.�������1�Yp�`f�S`�r�F�t�d�w����4������n��<F@eY���{�nD2���P=:66f�=wut|\DM]��y�Xr�����z�`º<�OS"r� ҳר�J�X�`�7�rVNS��v�����q���ύx��v}�^�ݺ��#�޾=��Y�����#st/�wƯ�"��� �EDD����㱟U埊���f�%pp���4
�6�U�ް��EF÷���,�_�d���T\\�{/��V������\�-�G�bB�%�I
a0KF,��=S��Yщ"���LvE������l�N��}�D���?�����ã#Z2�᫾�N�����)��20o?�e}^���T��mwj�_.��q���ꙓ^↑N�$���q�<<<9� ��EQ��sYiZE��@�M���L������LI��T������x��w�@�́�RC4�x5��-1d��c�pc?M��5���0Ғp!=��A!���|��OMc#��E�����nO��..//���5\R�h࿿��pm��z�p~#�e=:�ʽ%�H�(��������a����Eyyy�ʐr�ED��m����)���e����[�VUpr*H��6e����)�p�>G����G����0��>�]澟fڙZPg�%�u�����iPL;�:kR����X�Ms `a�ԽG���\Gs�dۚ&)�ݸFtE%U�ꖮ�n�=���lR�}O��H���#+���jٗ����� �����!���m,�l'�߲�kn�b:��	�1L4ci�1?��`��TH�Q�|��X�~pŰj�as������\����C���\n�7��~W�f2]��ZZN���C4ő��ݠ��!�]��\�LA��5�h���z� ��+ͱ��)	��_Y;L����8wL��[����VɫBb��0����2��v�WR��~�ldkn>/;wz��ԩS����:�_��E�q��U����r�M��az�Q����4��$+-%|h�����-�ZE�_�PPR�K���xٿk�י��K�^6�D� n�3���+��c&���� ����p�Ϋp�@�`hjH���ѻVVK[^�﫪v'�mg:�d��V�����b����L���WW�*K��;3�9�s$JJJ��ܦm�2�N��߃ۦ\�@0��R��7D#�>�X�#�O��c����ģ�>��8��w���E F ���)�O�5�@k_����{P�V�r-�//߂�)�Lc�� �x*��*S q�N-�D�ů_��2}�ԛ���}$b �Lll��YY���9�8�����0-II�����`T� |��?��F[$�)��;����8&"]����Ҧk���cG^x�:�'�R�h�"�xT���r����VVV������0���<DW��N_L���1N�H�Х&ɗ�"ă��ٕ�����PbP��q���������Jl����J���j����:�N����L[���{WJ����YiN��.�\a��,��`$����/00!B�sU��Ý;��^K���-s������%��&N\m#箛��=�mkJ7�]����`����}ѹ��w���;��[���$Q&,񀧦Z~Y���vg�.�����!�OȻ���U��-1�	Y٠��O�l�/�LDL���z%-��aK��!*���.���G�9W+�a�y��^��j���
ڧҸ�~���ى2Kw�]4�5%$_��+�IT�?N��a��Ĳ���-Cv>�7 x�ȿ#��(�e�r�k���0�.HӺ�Q�G�L���ₕ�^���6�'i�$^��~2 ��%4�ŜK�յ8ܮS￥������i���96?X�^1\�fN��u|��bt��J��N��k_�.Yh����dN+��I���k3��X�?��)ם�j���xA.r����0�j��:���#������t�Y<�>�I�:9x���fQ���ߏ1~:C8��E��~/��f�-��6�ϸC$/A�'�X���020��=��`n���W���$؂���珐�[�9�������M�/�
=B��ڂ$&���S0ؔ���$h?������y��m.?44����8�(-��\n�w0��rj^� {����ز����b�r4<��L`��":_�hܣ�K#�^�N�0o�:D����h�̻���	��vqw����Z�R���1|�h�&��#F�k �nV��k7'8�g� -)�
D����[?���j���?�|��\N[7ɰ}�S"2�Oc�FX�@f
ػ�g��w�Ɇ�V�?~�02����{V�=_�����H�l��O�_\� \-�Z~MB'ԍ�e�sY&3{)v��R�:�\A)�j>��3��1��<�`t�;BW
5�MNT���5�C@R��O�r��2��� ~����P���8B�^�GM{��7��b�uMMA�(��?�h6<��\�v&K�ٹ�U5���s�MNO�U��0Ud@��)*Q8�+��������8�n����]�
ۍv������Y�ٹ�>�]3�ʊ���N+��wM}�zۼk�U������U�nN|B9��˛e��\�&�>:1Q�o5B�q�|��߿�ҫ���Spgels"*x�Wt �� �yy|�F?�w���67�Y�Z�1�`�����ҿ|aR��7���§�6�r�[?��<+E1Q͔����ׯ���}1(v���s+l��&��7Bb/Y���8G:���$H��*�QA �6�:h�Q���Z��DG��@�<��&l0��Nˣ��f_!_�M4E�`	u>���Z��,���v��I��N�XC��j&^���������c�s�#U��:�	�ppX��r>󰯓�`����Zp��dt�v�.---��׀���+8�G�}E��f��mms��gҲ��.���]E�h8�ϯ�W�vS�����>�n�f�II�Ů���"��[vW�Ο�)X�Ce�A�ߪ�ؐ&Z�$��q��k���	>EI�A����cQ8X.���d���k�7v7
�<�A����:r�Z��Rm�TUݍB�[?��i�r�����n�΄l�DBii���p�?�P��0g
$�k��v`��4�ƌ~TW�3%Y�yrpэ�]Y�s��)bI�`Mq�To��k�����≍��,��-9���S��ILJ���D�Cy���w*�Nw�_��蒑���n�[�#����K�m�m_%o)���Cf�s����g��={{{���l9�kkj~6q>�_���m�!�� #�đ9�r)�qwj1G�h�țVPY����^���k�9eTsR��^�咯���,�4	jL
���g+E�ϋ��'�i|�ar��
J```�k��{:O����;šJ��HH���H=y�䎸xUA/����J���АE=R����g�YV#�sX%Z>So�,��`B���U`�r۷DP�@)����b ea'�	͞�g/����ROSY�?FS~�<�j�ǋ��`��(�h`X�YYg-4�4�Յzٞ�]��u?�������Z������ 6Ts�#~BҎ^��k��`)
�d���-��S������w �܊ �D0�cxћ����~�«�;�F
����ͅ���#�frg��`�.��h����	�W�)�8kr�����Y�"��S�tŴ�e}}}���F�h����l�{��(�U%k�,鐫w�(�u����ga������@2u�%
���9#'g�|��G�5��>�H5���s��z��-����}�F(���K<�@3���V,��廇�|)����Eq��!�c3�^�	F+J�"h3҆�&,W���%_PPp�E��d���eIu�Ѓ	@R쁼|L�W���Uq�e}U����l�������O���Eh�"<�V✋--����� ,���#�'�:'��-�zyz[#4F��7��jj�3!k��q�w��t��ud�Q�%�Σ����,��mfh�ze���L�bL�u�H�x�`޽{�&{��H�o�iF��|�d��t��b�F�0�����7��կ��\i&?��ٴϟ����y��64�ǉC�ހن��u��r�\?� ���sk�j��|��*���U�鉋�F0�?��hn��|ę��-z���(W��������8���ۨ��
�xD�k��r�5��bI���p�VD��t��>�7��لp6u�󔭶���g���  ,?g(��5��k�9W��t���5 ��.�����h\��D]v�YIɕ�s#�x�Yo��۲z����㓓���"� ��?"�eO�Y}�t]��խ��[�P�n�C/S����ٰ���?ޜ�0��5��_l}w<�o�����Rf
ɦ����2����ݱGˈ�dš���ǱJȖ������s�_������s��u}���~_�W�C��T�����r����w@]]���jǫ��'�P�^�zU��RSmՈ`�����]5���bb����?:�{���:Q)�]x�ߤ`ύ'�ѷ��E����{���MQ��-3��R�˅h����ʚ�S�#��E{�|o##����*��	�j{LL�����/��8z��lYf�i�ؗ�LĖۉl&zzCu�����9�k��PE�3�ˏ�ě�����1�7�J�D�'���P1���Zr���q3K�_�l3{#ZL��5�#�U�7����p�I��P��s1��n�����r4&�`QҞ����}���J5�!�-:�2�8N���;Q������ډ���iz�@��;b�ѷ��ĵ�p �;�bK�VrV,s��RZ��\�2�&I���=�t3�R}�yu81�P�U��1a7���=KbA�����q�d"����!�Oğ'�Q����N�M)^�ǹ�����\�ݺ	~��l���2M������`�5���ϯ8==}�̙���0������,�R��8��ɑR��E�i����ɶq�퟇PU!�t�`0<\%|��f��뭷��/����Rn7PM}�L��$y4��~��8?�����)��Ӄ�QW	�<��~�q���F�Ѭ�Q��h�0?�1��G�;���������e�v6ܷ?9W���
�<M��D�x|\�[7
g�E9�'8e�AѻTg3��΋+�s]Wq-�s���_|̷�'5�o���4.�@�%܅�oWёE ��o��y��ُq�BS��zz187� .� �xt�fg��ɱy��n].K�ZU�3�0h�l�܂����{!��۶@�����v/~B�G$|��莓Ԓ�,O]��T��'�� UUU5	�(�Ք�ɿi�[USs�����~a4�ald��Y&mk����H�A�D/��� ΀�{�w���FG�#��j#�C{��]EE=��t�9�S|�?�T�`�d$%��\c��/�%K���g����jH�s���T��ʿ<�c
��o��<	J��#g�'1L���Ǘ@R<�+��ۣ�:�vR�.���9;0��Q�dPL�@������'CCOݹ݊���,7E�̓ 
�	�t�/��';���U�
�\+m����1��� 0�[I�^Vf�mtB��Q���fI���x\fp^�hҕ-�-�̣q��a��}	����ܾ$$�gt��B�+���}�~��&IjK��O���]DV��e+���T����|����R��V��dh����
@���̢�TU��Y�N�?��M�"v����.7�1�;ުNX��	�z�u���vh��MKX��zb��T�ѻyꝧܴ���0@�Im��������@s;O�@Yw˅	8�B��5-#H>�N���(=~�d��x�
7Z��Rq���W��ޓ�d��I�
�L�����6�ZZ��J����ж�i(�Ҳ�޸*׼�����`ͷ���3�Zl/��sa0}��':�����|�����<T'����Ƅ�H�fg�M�U��/�s�u�v�\��/%a2�h�wo!,U���K�����N�����d6^��Y����="�hQ�81))�u����Z�J+F�e��D��R��z[5C�b�q�	�ޔ�y�1P���4���V�<����j�gPFg�)�C��~12���w���g��`�ǡ@�-^�o<�Q���`��-Ӟ*�ڳ3:;{��߼���y%%��Ô�#��������y`)�9989�6��Ov��><<<�������6������7��&�ѣY�h9�յ3���-O�4CZS35l�9�~Ag{Z����ל/�t�*0�nDfA�Ɇ�\�k(Z(��D���%���
`��:@of�m��iiw��
�y�@���A�h��|J��(C /������.ްis��)��6��j�`���l�2 ��>��S��Y��	�O���Op�3%_����3ȃ6x��Š4Ի6ic����)��0cׂ"��H���|��H��6�ѕ��vsZ.o~��O�J�,&U̐��$76>��쥤 ��.0p�ΏB��9Z�,��
s,�_J^>h�nk��X�R�>J��v5kml�����"�Z�Kx�����V���{���U/x(�Z(H)�L���/g�)�V�9����}0rc5 �V����+�qÇ���vӕ��u�$KܸQ�զ�bI��W|:~�<��b���L��!��
��kK1��w�^4���e���2 F�[|�ٱ'�F�"�+f���8d)J�궑�Af��u��d(p2O���{�r,X��Ҍ+�,D�r������gYXn���?S��s�q%5���)A��4Mb.A�'~���l�aܬ���c�8"Q�G))��P�x�n����?����<~��h�͵(-������a'^���.RAW� ��0|�/o<���$��e��1Y�0YM��v�4��t �������j��G���X111�n7�����bH�%���m�`a��b��Z-��ZZZV��#' N4@i��s�$_���w/�Z:zv�R�<��;)����h����;m�in~�[>X���)�"Opz:ߦ���T��0�')""B1���o�+��@��,,,�q=�==���UQ9/�!��tt����䦿�f�l�%�P?F����`h8���μ���!tFP݆�����ÊI$��~�B��ь_�E�FW�.�����ՕcƐ��R�*O~���W����� �,>��Bk���	YX̬w�P>5����
D���Zե&af��GV���!5+kN)���`^�6�B����lkd�AL� �X"�4��3��6`T0��S
�Z��"�j�����>��ǈ'�k����̪�����]]eS2�̬����=Ӷ�;��m~��'�O�а{zzn���<zt����������k�U�vN.���b�����?~��=�V�����:cRvvK�4�g�+�B� T���%oc}e�����-{�"x2��Pc�3�\�鑥�6�������8�[�4dQ��y}P������y NG�xzy�|�rÙ�-��n��M#X�:�a�&I7�-"��)>�i{m�
��Ž�s��v�X���G{t���cbc��_2F�F,2����$����:��hY/��ˬ��{�yfb���kc�EY��z!|]q��6�Ho:��=RP��|�NLf�]��yj���_Y���T�dF��G�"�&\j�ꊮb� ~�b��d\aDK��8ղ�d��z.UA���=�A?�^��!�_&�Ro���UCc����w�2op���W���6���`��ƌ���hP�_2	��N����-[�+�ٽ1�G{!����B2��~H�܁6פ��}����F��F���� }Y��k���������I2�_՚��Ϡs�EǄfC�H�.]ZS �L5��i����N��΃y~�Լ^ohd�(�μ��8Z`��q��hk{�oS���蛗.^T'�k�t���ǃ�_B	 7@��XH�b3����
wq�!|
��w�]tl�zʆʓ\Qjʪ��ム��s�0�����-�6.OT�'�F�<Zܺ���FRe���t�ƫD�6��Q8�]�s���`O�7G.�D�����**(����Ԡ��h?�]+~XB|��W�+@>�^�zE�>�������ղ�hj���6jsԔԙT��+!��`��Zk),�斖J9A�9�	�!�g<ԁ/���j_�ٳh~PޓZNN�roSU�n�	8`��}sN�u�$���9/ ����a����S�~����e~��'O�@1}
\E��:��u�0�xv�ӧO?�\�<�q
�S36NЋHL�e! ����O�"1P���5x���l��a���C�
�.�%�h�ϛ�ƻy�ƈ]t�iOAa���	^,�#�����Pd9�F��d�sƸ	jpMs�VJY�w���w\&�D����܊C�Cf����i8��	1W=������J��2!*(ǩS�6���Ѯta[&��{�<z!�p}$�f�2�u2	���]-�d�Q�BM��ty���ƞ�d�Q�IG�tSm��/�uh����{���B�F�Rd;�D��g4��Cq����ۯ�~�زH=1]��܁̣���W*�d*��6�@�2��B��W?�ĔE**��Kwf���{JJF�� ����S�T�lޤ�H���a����2�3�ˌi�̯`�M.^�T���a�	�8R܋F���T~��ſ|�Eq�`gI��ϯ��w屩WlTV��SO�B�
�Ɔ�y	���۷����Q�`�\��(c�:>t� 3G2����nNt{���g�p>���ie��R��ٔ�����C�~hKRV[U\��W�w����ԲM~ʧ�����;p��)Q��+!6�>|K-��$�4���p�C��{E�����ԧ�+����A��3:��������	[)��@��q���C`!��JH�2���J��ϫ嘶��xC��o*(F@Wt
5ut�!�eJ@\8�
�I�Mic�#d|�e��
������1���jNj9�AW0"jo�B'~�o ��ε �+)+/���1�����JC�W�յ���ڡ�[��A sM��94Y��BT���{��;�'z
�@klN&�NCE3�S�����[R�- VjG�	<%�e*�4x0�s|�?��5Y�f� �&(%��[���mX_TŤ>���E;��~�����(B{����;R�rccc���+��s�q��\��˲ 6o3���h::��8���������F ]\y~��M��:;��]��~����a�f�	4��@t��<��]i���fV�ښ�U_��8�7�%�$ ����ٕ+�SC��M�6��~�C�
Z+o�5_:aK�@d�5���(n���J�; &��(D{fMgn��'??�	@Hoz�M�ҳ��Pu�`/�K����A�Z�,� ���V�K��ŉ��^߷W�?~� �Ҿw�t���y���1_�Hc+�4S84�w�<iApr�S|�-��Hi9�78�b�A�)��2(lh����S��П�U�?;;��}+t<�"���
6��&����znn�;⛑��՜�"��3��b\�ZڴOR�w�����94b�%2�O��T1��H�yR�����P{�;���Tm6;0��ou{� 8��B���ء����ϟ��\z���72ϓ"���e+�E����/z�E�S��Dݼ��X���K+游D��-��B���@{�{w�"ǹ��6fm�[�ܡ	imD�x	��\�$d;/�[�7o��̇^t�`��X}�b�W:T���&#�D5677���\Ϋ�����lӰ�ɡ��Na����ϋo,����w"�b0L7�/�6\�l��|F�;Ӫm�F�^P�~d4��<�t^�/��.�����y�;����� ��?���dd�t��z�8��/��"eL�vv�G�M����a.4���8��K�:{��h�2�E��a�y�8�OE`�d�C:�rP_ܠS��i�p���x�����t��DD˼N�0�v����`�����@\J������Kˣ�8�ص�y�	���Jw$������Q`��L@;�YT�Q�nV�S<���\BZ�A�5�����	Hױ}��J�.�v9Z��h�؝���eq$�"�M�4Z���H�C
����`��$1}e��YYYfO��Y��d����[�~"����70)�K��-��N9�-ii�X���[��V��*FR־3�P���c��8�0�8hҤa
2� ��vW�0it�Z�����b�P������l�����ݝI�����Fe�v��|4�{+�0�c�^���C�^���̌�`>!������b�!���=���eB��ݻ�#���M:��}i�<C����f����+��P3s�����)�oK��\���_�/.&�¿�OP��o�<y���8S���N��zS]���j}���ҹG[��MC$)�?�.Zm�-�5�~c�W��-��U6��ɓ���7���b��P�Z����;���F*廎��O:3Go@Ē��[m�W,E��:k�|��1b�W���B�E�f��^Nw�p^��]gA���4�oA�������Jܒ�?A�0?�e�&�������������n���̌��늁�h���˨����������� �9
�@ȼG!�$$�mR�G�~����H+ �<����+j�U�,��
�A*���׃y#��:S���M	$�[rr-�5( �6��8��HMʾ�x���`?�AG�43��l����T����[�0K��Uү}�wsske��er�!��n�zT~�����&MB�p����}	�Y�.��`٤e������TyII��4�|���gɇ��dx�L�?�����e�I_u�P���3O�>ʭqi�|�s��'�~�Z�2���z'�,C5ndfV�;2���ۛrs�N�enػZ� �1��tim]��j��E���o$�$˴�[���Q�^=d_a�c��Z� �	�VEi�bKP������S�F�F�eځ������ƚUTTcs���.7`��u�v������'(((.���۾��d�_�w���$5�b>�}��gGr��F{���(2�0�ٛ�@[��_�^:\&�0��P�g>���iI��f���]	�ޠ)�jttt��t*�m0M�͙�S����F�mi�U*�4:Yr�hdb�(t.`!�&? $�<:���^f��___d��Y��t� ��;q����M�L 4��'۪���I@��b�f���60��X?����Dl8�$��L�&��uP.���@o�<x�Gl����l[���(������<w|fzz�7d.�ilh����už��R��Y���u�������ŗ�#��[���G�"����۠�X�(c�Ƃ���r�?���I�D��(���h �������������P�V�I0�SjS��jhf�r�/|QPP<�?C��f$� �D���0�*&���>))��H�ڝnۋk*�ќD7�s��K�M �j��N��$m͝�X �eo�t����R��d]������ǿ~�3��nf����{��h�9�4��.�ۤ�S��w%�/�����M���MB�[���u��񺴭����pA�� Gh3Cggg�
ZW|᷂.z���!��?EBJ�X�i�J���˄3�ݤ����m��-.���S�,"b_�;u��,,�
�/�����Q�X�"�W��qe�
���l�8�u0̑#[s�\ڷ˒::�k�M=
	ğt����r�.]��HGhYs>p5&��� <~�y��^�2fN����mi����3�k-X���������hi^P��(���Ԑ���M	A� ����n��ډZ�@*Z����#�`�WK�^0��̸��63r�s�6��kK3;!��Eu0������9d�x��T��l��û���C����hi�@l�ˈ4��L7���&$o����ɟ�����4 z��� yk���8������Q�D��
�j�����r�ᇯ��Ê��4��@�N��J�|����F�prr� �iYYY��]WN4���R���ԏ
R�b�f�?C�>"kd�r�O��Bz5R��A�*S�5�CrK��/mi����W��:��x	�'��ހ@�}`���#�����ؾ'h�Κ)��i߄Oni��;ԩ��r�t��3t�n�J��h^[&��T�y:��d�ӧO�'��d��b5�Q�~����yJc��o���إ̬,�dbC T�M�Ep��5Y��%��UT�a��?A��vnm�C>T��ߊe�ֆ�ñ��I�$Xmmn��(���J������J���Zi��~d��W�@��JB��޳s=��5<��N����� �S�Vd(����}��ɜ)��[`�K�4��b���ğ�3�Tf�d\G�<�� Q*�m�N��[�nQ��%������==�*`��h�BMM-<P�ܳvR�d�P�FƁ�7]�""X���KX��r��֖��v�����C=H��$���r>q�p~�,�J�?Ґ�V���.jho{��_he�y�ٴl|�|x<#Ҧ�5d2ϊ_L�@�;ƾ���"ߚ!�h��3���u��߂$"��tV�����@�a(Hϐ�_r�j*��
���Cp��V����ȳ�0p�9��q==��p�1�{_]�X�Ǜ�2�_n����+���l{��9�m�	�P:�oE����YɃ�_U |`�:L�̪֘7�����c$r>}�-���up��k�r ���c]5�D�>> QQQe���摏�w/nv&d��:#�a��;F@��O�^N,�]YZ���e�z��$y����ܱ}N_����M1d���[��A}��Y��@���V0K��H/7�d11�����������C�,�������̐u��$�eR����ʲ������4��m���ў���m�I@�:���:�@
2�P�LKK�Y�T�4I�Ίz�f����W�[O[08:\�5�'[����B�Н'�I0��v%�e�+�:��Ob�322��_�!t}����u��FU�ƻ�A���l0���/�I�^j��{ޡX��¨��.��b��֬_���Ɖ�S=�`�x�:���\w�����Z�+V�&~�b(�C�<E�U*�+�~��>"q�=;�gW��P�l���.<�/���If��ϐ�D�;e����ͷ�f�D��߹�F1��ˋ�=��G��1yl7�`i�Y�w׷������Α�?��~jBF�m���qc4�^��O�y.T�>�SW����h������F�o��Ta�P����oo�}%�~>&��z�7e&d2X+oYZZ��E�zF&l~f?c/F���_=��6���S�<�G��
bBCC3�p+�]C�r���=����@��7$G/��`�8*)�k��ڶu�d�\�!;D�% ,8���g�*� �g:g�'a�NhY�X�l\S���)�,=�P�[G�P�6�PSq��F�����"�QJt>�|�ZLO�A�}�p<`Okl��Μ1ϖo^�N��y6�S��ꭷ{R ��k��S��k��g��kE�M����s�Dmu������Qki�K���N��3nڏj*;S�	��q��ʺ�&O�e�}FhI��5�:�)vSY>Ǻ6=:�}c"-,�Y;(c��gi_H#�qP�[�/���J|4Wx�%��F����NQ�-9�L��-gާ���^ յ2�@iU��}%��M�;��8������;�P��D���D��V��o�JT�o�F>��?���^m�p��G<O��Hm	]�!�\Scۑ���|u��<k":�c�i�+�i�PI䃵����ᬂ�釟[w6�>s8��x3R���D�0Y��m�꧘X�OY�*Fe��D�A�0�dU��ɗ]�:$4�b��h��f![�����=�M;��=����/��Թ�˹|xy��Y=L�����$�[���^c!�<�$F~?kn�z���~s!�e>�q�����:s��p�y��'s㩛qSLS{��Rm�p7t��y�߿�9p/�&S�l͜�Tz��<e�>��09u�+K��_����~������T7m���h��-t(SW���}�:/�!�$���i���B�Ģ6s!Z��-�8��˗���9�n!D{�I��-��mڲ���;&��6ފL/''G\��ئ�x��������!��CPe��
�nd�e�����?z#HC�[񳻻&���-4"BS�:������b��2P��mc֚�Q�����(B$�>n�+}}�̣=oK���������k�"e�0��k��?g���$ւ�D�|rK5y4W{��_%�,�������3_B��8����@��@N��SF������Ҿϭ�!oZl�S�J��n�
f����A[@���6�.��\��g�����^z���o�E֧��#޿�C3�-��W�q43�.۶y+�p���{��#|�m��yA��������83C���{�i�5T�����䝣;g�n[��؀c�B��3�1��-�\�T@h����4�Uj�"O=��>�#�T�r�p��M���sn*�eJ���Ȃ@�BZI\>nf�f����4)6..먾�ܳ�q(�v�2Ҧ?v�T�w����}KT�
������n2�mn~�?���lz=��mEEŒ��,�>��p<�������!�	'�L�Yo0*yINV��64x.�G�f���X�+d7f)u}j7\��\Ӵ u��g�]*N��8�1z�o�k3R
�%����4�=��_��j��<�����yV�����~�[3�ڂBQ�}X�G��	:��fQ�Cb�Hn�C��P��UO��WQ�m:`�4Y���G�.Mr��������Q��O	�V�����e�㮵�*�V��@�F�)�0��縩��A?����Yn�)!�l`���/��c���buԡŵ����_�GƦ����օ6��n&�9���\58��w��Yo��&b`+���������4	Z6Z�����+���� �w(���Wj��\�u��N�������C����{������sԹj/[��:��@��C��t��#��*���pm��1�-�C\��0���쑉�?KF�L4Q�0����>�������4% "re"���d�?����MC�D�A���H�v�#?߃&��{��o;���)�?�fq/���>{���)?a�P�*����Ä13T�^q5@�Og���H1 �zt
���9��MD�A�'C�x�%�mҺ1��ϟ?@��1%�h]�zUbO��g] �A۽"	<{eL�Fs0;������AA>�O@��652�W =�����ɐ�6�o�E8Q����!�mlj�;v�D��M����=��h�<�s7|���͔�����J��=Z�nV��/�h���AO�fgէ���=�����_|��8*���v�xf��`[J�3J��������������������Q)mo�n2$y����qS^%}���@�_[uX�'^>#�j׶]XGٛZy�t�VbkW�]�;EC�Tr��ٹ�� ��P�&��d@;y�OG��f�	����bZ�.	
:�&~lSS~QN�Hek�t����^�
�DV˄� wo�����N���xy�l�lFU}�!t��Yq		���:�,��7 Q�u[�Zr����{����Wr��@vO�m�NF�g�2�5�<� �74��s;w<�@�gn��݃):�GRB���P�9�4��$ pݪ�Ot���M�Q�����Dw���x�K*[�K�O@��S���HG{�m!�K��Ši�?e�xP;O��O�\\��z^�(:L:3ohkk+t�p�b�1,4��Kνw��3������'�?{FFz�����3*�ުyDS{{{��q�<�H~Jc�W���wYXY�/��Q�0�1�z��
fڃ�qD����+����u�*|�jب)MQx�?΂�X���o~$��C�}ra�"Y�it��ׇIDޓ��ah̏�~��ݻ���Û�)L�,��Ϧ�{�l���'x� Y��G�PG�V�CCNJ4`����L~���6��K�T�C:������T���q���	�m�O\�qM|(�yћ��@��̐�N��j�����Ӵ����5�1��f���a���������W��Τ�¯J����a�dW�Ж�Wsp��N� �����+����j���#�L�-,,��P LXOo��o�E>$@�@s]����'�Ḟ�7�����Lt�<K���~��z�ݽt�����r��x��ϺEm����ً��XHZ��ɐj(u�>>F�|�)TV�4&ߟ?~� z����0p�'��۠�����x�f����O�Ő*�t*L����E��k_SP��>���VG^OO�:�����6��v��B�\ �2O�^N�6��*ܮ�gH�682�a�Yd߾}�0�	��ૌғ�M�ǂ����_�45{6.Q^���˷J
+�~���'&N4��ƺ�v�f$���eGGG�C��ʖ����������ѺY8r�����솆�
�k$�l=І��[�B�G����b�q���ܖ�S�N�x��,��~hu||<�_\��:n�ʅ���~M�u/��<�r�R�������乍^�'l.T ���㾺����Rj�Sk� ��t]>6xN穙����պ��<����E��$����	����7B-���ihO;���.�j�	j,'��� �'�hN|��'X�ߌ��������u2�79�k{�p�44�����T�PV; �HB�C��@ͼ))	��!����8�n� %0�8�>7���mj��1wU-�'x�E�X�
3�g!>>���$��L���]p�"/.Ϲj3��ѩ����`�s���bl���5h�K0� ��2�D�L�ی�z����s���)9�%��ڃ��$˵p/Q�,�p��vG�H~`+����>}r@'�t��E����
K�f�M��8�&��8�Q`ٯm�NHB৥�o|-!R� �*�Ȩ�vtT%�rd�ύ}����|��X�����C�̓�P��u����g܄�Ms� ��G^�I?PSS#��	=}y팖�V�F�$&u���G��SS0�@`��lįcO���֨ݺu+ r�l�z���{@�)����:z�����6��eeeZP%Rs[��FйKr�pz�����5�$Ry��QbRSyڛ�gwA����\�S�L����o:��3Pv?���P-w����hhh��d��3۵�����[W�0�V���c��QOlA�8�K��g��FILФ���M(�'��E��*�rrr�����]#c��W�5j,�K|3`�B��ε��>J����̮��k(ml��+�
�����s�p���[��V"��ΡW�
l�b���q���v��,L-C_N,|,u�=�`�\�|<<������z��{7��UUU�:�f.]�́�V����.��R|'tx��dv� 5e>����+=�72�W��S�jfk�������i��x"�.���r��TCC��9�bRf��~��Ĵ���$���>���\��\XX�y����63;[�% �ONzz:w�jFyx�O��G��������h[p�x'��$����Ycff�j�Ę}����q�um��_���N��{vv�G�ٹ(�^��-���c�����~�|������;���ⓓ{����`TB  ��.N��n��yu�;���H�v��qt��=��*��
:����f��C"�2 �h�Li�(7���WTQYd�'7R���BCB��R�v�׌�����F�����07�g��u�0;Q ��5��V2��	t�lm�-��Bb��Ĥ��ʓ�mR��D�X�3�X6��t�u*~*9��.i$��M��,?RUU� �9Hy��+�稨�hN��@/�$��Q��\�,M��#!���yʀ��&L�~�3��?L���{����S<�bU���ʣb`s;�6����W��B�;]P�xKQ�)	���c�kv����m8�}������A�9�V��e� 5�%Tk�8���?ߑ���F{�V�q4s�z]j��!�!T��_.�����a�0�bg�ڷ�2bQĴ�������7y�sҮ����VŏY&ȱ
�U��T��pX������T�]K@ۘa�.`���`L�)�g���'1�����^s.VsO�f�_C��g343k�S91���5_C�m������u�`��Uz�HV�����z�x��+�$��x��w���?�,�#�X���ؖ�JȠtbu�~IHo��F\;s-"�ݻ���Zw30�&�t�O�K��ڼ���(ݹ��?���ջ�@:�a����nkhP�[��	�y�l����=�؛�v���kd%zG$�j����D�9���G���>_��q�
Ŏ��{�HH����;��c�	.��=Y�"�\N�8m�g��WR�A�Ӻ�0S��g@$6���w�X׋�k�#ebb�����痍����>z�}�;m���#��'�YM]�l����Y9�eHcJ����J)+7���Մ���A5f<	B6nx�n��7��ξQ'��v�~���h!нnF5���=��l��B���'�W��i�L�,��Y�ʜ��,��w�
&5]V��Igv�MT�\S�� ���˝챡���S����N1�Ǹ�wEr?�tz��2>�|��By�Wq�]J��MDp�ܪ�����~�����ѥ��dF��U���ӗ> �q���B*��ګ�β�\�;�n��޴�X��L��vG_���?�o�;����v��~���|�\���M.��<���A�����������J��ϿG���4alU�׵��v�O���906�R�&+��Vа�[��6�I2��/��^���^BBV1���n�F���e�AOI��{���:י.:Bp����6��ù���'Ũ���<kg����Ϡ����O
�Az����&{:p���L�7�ZX��rm�3��hC��A���6�7a-y_-Z��\�%&��T��J�֫��~�5�˃�k!`(��$a^}��@��lœ�<]�ݿiΞ�s����-NWgH�?�>�_8.�� �4&�o�� ��������$ r�Z�ʤ�<a�=t�hZl�0���Q4-��M%�(P��EG	�>R�	�m$mggg���f]�t�Q�IO��H�*A�#З�J���:L��P��I�T����bbu��
d�s���٭[0����d�T���Wɮ��1���־/u��a�R�Z;��rd#V-��%��*��Dg=�ͺ�U��'ƕ��D(���R� �),��W��X�&ί��w���
�����Xk"��f�4&,d�A�"r�5��9�H����ݛ<��t 6��.�n�땯���_��'I��H�jq����N�]諨�DGF���M[�����D��Iqt枮e�̲�+%1!A-���kX!ꀸ�{�	¼T����|S��Y*RS]z����M�J���6�:s!fu����ѩ��/��9v�)�]8�t���L���e���7��$��M�FV'��i)T��`���ӅJv�K�V玩�)rt�KA>��a ��r�Z;z�hZ7�Tx2�|�W%��E}#N���2���p;�&EHrZz</��J+5-��u�.:J5걱1�{��w~Z�IWA�"�ozR�W�%�ݻcRRn_�p!S�����ꪪ*taS0��Y�ȣz�/S���̧��QT5�wT��'�E��y���=���mb#%&�7��6�����d����w��s�b�Z49n<��X����(� �łW�'j��
�~��3��mȏ7�cu�Q�, �q�%���q�&r�=�d!Qg�
��&?i٪���F�,%2���#ɚt��D_���[A��PhN��Z�l$�+'�tmҩx�}C��X��@y9��h�(��;P��厪�]T������_�'Ȓ�p���?�~o���$G90;;{�y\�רycYĩ������J�+:OMn�2~��Կ/�� #��F�A��A�ɀ�y ��W9���.$��ʨĖh�!�;���f��K��0T�Y�{�O�[�{��K+��X������gF�o�}���/�Hv�a�.\w}�_G�s�`�:���1%Z�����?�dh@&T���5��H����C�������K���6;C=�*QMu^[�9}������;������x%��'��Wsg�祟>��U=oimM6j���0�t	G#`Ҏ.��z�uC�@��t7�Ws���!�./��t��bl��~8���Z�m2\LL���8\|�qd����{.I��S���tHA��_��ט&������oJ;�P?�0�d���;��B�C���6���N�8��7�b���P����t��NB���B���kM���Ҁ�!���Ǹ�����{q��Qa����e��bH���1	��Gxq�.�=9��} �ސJ���ŉx�V0Pۅo�S
[j���=깾��lC|����/�4�焄���|'�~����@(��@,~�.�����ꄸ�C9&��^ܾ�i|��I����ymW�j7{�n��]��Ŭ;1�y*�����"�]�������|��"3Ur��AV �P/��'����=�m_	C�^��
����3�h�ݐ�=s0N���)ce�$���]Lss�c�𷭭�+�3u:�t��Udee)?�	��-��{ŕ�V�T��Օ yi��<r��5n�wEh@�����a������Y�K�q>��S���@��pLW%�&��Y�H!�,�`�1��1�e+1�z������0W�����ٝ�ͤ�s�ٯ��yK���#.��(xx�`��tp�rU}�]���z��� Ө�Ǿ�N�n����C保Bd�T�v�3r� �^�<�*e�3�3��ֿ�#]�>�O$��@�srK�"��޾8X�г���yE�3Ӱ)8�C���"�GNq~������hw����Gt�C�y��}LLhߔM�E�i�A�.���H�"`� �G�_>n�ϝasY�c��s��ە�0�w���W���Y��;�[��͟����s�*�Wi���Lp���t�4(���i#ło��=
��v|���3 rj�r����"'��g�oW���p0�+Rk]����	u,�
��D諆� d@𲽃X�o��o�c��΂n�Ѻ~���4�+���N�R"�eݎDy��;�9&X��r��C�F����\�'���rRT��}���-=�z��������:�.	�|w�e^#�|�ki�^�_�+��}Ļ}�����:�0�U��n>b��%��~�'��8`�z��q�R�mieu�~k��p��ȩدGԷj�/�VE�Q�����^��z$H����~������\�)�"�Py�]0+^�	�{@)ESö����ǎ�OK=�nD9���Vf��М���X��E����l���u?��Ǣ�ƿ
���|�j�fVTTD7��\(3?$�D�K��SY�LK��H�G�OaѣqC-is]�\���%�{A�݂
񧡩1c\�.ҳ���.ں�A��߫��p�1��F.Kq|����4�^&�<j��&%0��Dı��S��Ggs�����؈/̥���_�v�����;�]�LX܄�>S(SJVgִ�Ǖ���Є�s��m6�x�Z��3ӿ|12��I�gJ�%`hl�T���AnSb�\>�� �F�\�d���K�oP�WݪŊU�Kc0�֖�Բ��zً������v(�Y+&��?��N����L۵�/��0�ݙ�����ycF��O�vz?���hn#�����>==a�m���~AÆ��Jؕ�Q�8����֦�D��R^Q1��D3�ܞ9�ৼ�L���^��g����b(��_w3��4%��MKK;O�i�V��P�s����3KK�.\��2��x�w'�X�*��V%�qb�<=:������~{[��u�+:��)n4ջ��ː�k���B�+������*R�X��\�e[[qa%0�vCKd�/eH1��c�����H	�>cl<Dΰ�
Ω�僱.w��V�;9]� ���,ME°�C�6ﮏ��'QއTU?G埐�/�Ȝ��+\��X��w2����5{����hH`'g\�E���zg��R�ʕ����������+�q����{�`���U��Ѡ���F�k��ms<ވ��a�C�o"�.�l�Aq�����,x������w�ZU��ɣD�b���Kqo�e�Fw�9�A�m.���0�N�e��*tBG��!F�2���c)�0�?�K:Q"��ã��p�8\Z.�XN�h�S�(ݍ���V󠳫��\}����d�5���i�^j0�tk��O�S�ŭ3�a���p����TK��;���|ͱ�P�2�\�̊kpW���U0�Ĳ2n]K�c/p�ى�ۣ����m��z��I���O�ѓ�4eZ{��=��f��"ܱJ��lz��(O����Zև�j]�G��v�mmB\���5>�2X�Uo�D��`5�� '���Ғ������Bw��� ���z����IA��s,������TC��o6R����ʆ+:��<��mY���2I� J���fV8Ǌc�a���}F���;��f���3Hg�]V�mw�[�3첏|��\l�t���w��߿Wo�Ud�������k��?[���Ww��o���G��!��e�ZS*�.�͚��T��	M��u��Hu!k�%F��,!z<fw�Y/��C�0N��imW�b���U��YvLI�~W����ꭣ���?Pi�	A�k(%����;F:D����nQ�;����y��w����r��3s���s���Juuu���  emNXbr�x��ߔY�&j8Z��/lmm��7�����$CI�2�A�|��h��]ώ�kr�Ôp�0�V7��v����c���Q����v�2���`����u{��_E�K��Z���-�}
�7��\>�ÿљ�s�Y4��{� ����!�6ݾ��x�m�2���H@����5�7thAE�c������!�<0�x�4r�2+���/~�|	�W���Cyטx��3���r/���$	�������`���wA�����.b���PX_��n`�!۴S�B��Y���)x��T�]�>���K��⤧����2]���f}��Ye=��Mt[����<-- ����![K!&� ��r���0,���[����W ���.h��M�F��Ѷ���Ty�"X���ҟN��-�*����������a�������sc�-�>�.
�F��[QK@�Ƞ�hŽ��c�Q,r�mu��X�}}]�cî]��8-�8��N��~���i0���L<'y��,��7��RR',����"</��^�S�U��3��uVPT4b�kE+����}��R�۾���O���D����{�AH��~��b
�d4�8�@2�p�!V'::ziQY�x=|�7+�Q�χmP���+�������}��"4cc"d����Z>k��Ge�L���N�n����r����^�z�&��#�\w=�6��a�8O�yĴBES�7U����l�}�"�!��0�W�1�����1�;����P��\��Ґ��򭍗�0�A�U=&���a����Ͱ��/�&��_���ʽy���%��a����
�>U;�d�v�{`��/-P_5uu,e����L>6_������Aae�j��r@e-����~����d5Wn��sc �b���t�b�W�
�c1'�,�ڡEЊm��43\�C�*�[�u�=� hҚ�=���qm/^�W���C��4I�Y��m���n~���<�$ro_�DB@��|I�T[r)w��ۣ������"u�P�X�ӯ�N�g��V�'0���{� ��[\\���l���:��i�E�յ���d�����7��myz��QkK-l�K�*�!����X��6.:�e9����.�G@2z�4�W:��:���ro�c�KY�QQ�u ��0����]�l�?)��r��cȴhUR��#�Ʀ����e�6�\7"�Z>����GZ}a?��o�n��[x�B'ݔ���b�[&/��q&#:J፾��/+��5j����C�?܇LUkO�*W3c?��T!h�P%�7nZ�ry�(\j�(ǣO�)�&��z��{�������s*I���AI�͒&u����Pe�i�m��&�*����<���ɘn�<�$?�
8\|lx�H�n���'2�:~��\�|W����A}��亁�Z�j5[N%�_¤�%���4�����S]dV��� �v����R���KN�W
��R�-qZ�Cݡ�h�8g[�G?ܰ�/���7/�ӑ� P(�M��-7pB�!�u�?>1!G�7�OLL<���os�����}ԁJ:�">?#��x���>᠍y?:9�3�X{!����laz�+P U��7�v�G��l�3��:�Bw��z u�V������I�� )�����T��u1��� ���2}F���4E��Q���Q���~����"ޛX���9H��6� i�<s���%�� ���s���Kh�'Қ�r��J���8|y�ݵ�Q?J��4$��3IѪ����!�6/_C���*sp�O�N�'$$<�e������uH��g�"&(�sP��WW�n����}�	Y4��
�s�0���;e��"���t1�9:��`�0|�֗㇮�Ӈ���;<N�2���m��i{�9�lP�s�Q�3(X��0b�ߵ�]V���P�tE�B~8V���[qFe�5�ѺCb�φ�O
��Z����D����дWgff��Z���;�|�O��شB.�:��=���xm���k9+ʁ3�Ѫ!�T>w�z=�����9�3�lp_�-�A�c[�Pd���79O����W�@W�f���q��0��/=��O�Ѫ[\�۩��GM<�^��F���.Q�G;�b�rY)�����ٌ�㦙I�~�3��U&����=���2��>4�
�}������|�1::j�5�%��c~s�w~~^������ܦ&]������������H��8KFv�pv�i$���MW�M͊��4�O�Rk���x��y(���&������q�����E����֦a|����I��0j�(O<\��^w�t+���l"�7�ݮ=vr�N�22(�{�"_а�?K�񥢴���P�-��0=��ď3߸���Ӈߚ ��~_�;FF���XUh����m\�ɊMA�Y����K��Ǌ�������f��i��4�$�(ʼ/�
��A�W��3����gY����nϾ�mk�'ə�H*0���@������S�?ikc�ڵ"�����Ke�c����� �hr
��߿��P�L��sz���t�{
���Hr�ʈ�T��~�#0&e\��Y��]^��;;���7��~�������_P��/�.:������A�'K-�c�d���AJ�E�Co+�7�y�&!h7�g�1�^Ն',C�u�~��_	��_ܚ��mO���]u�s��sH�����/��s���&�G/�x�՗!��'��R��eNN|O��$6��G�>�����IQ��Y�J	Sӵ����G�`	m��딓�1偭�|��g�h%�Z��)C���X����q�{`��į�.����/cO��գ���!�m�$�۷X�L_ME��HZ�Nn3������M;��(B֟��{u�+,�S�-9��b�~\b1���z����m��� .\�U�<�M�&r��M�w�m�ױ��	��: G ���]�xƘ����l/�揷l�U�]�G�>AXN���Q��Ѐ;9(b�&��-�m�htB��r3B�S�'�A���\�w�v���?0pʪ[�7�a����&TAʨ�(�F�듲F�ҽz�����
�UU!l�N����}���}�kԈ4��7���nk�t����}_7�j�;6;_��*����XX�[Z|q�f�@@�#G�$=S�>a3~��0����L�~�#K�� 	���;��6i��M:7'E�:�n�"HJv�2U�ZV�� -i͞�o��G8_�`�?���? �os)���.��m�W�ڬYka.::��g~�~�U��ǽP�xD��J�����~!������[ɟ|2�7=����ﾼ?9m�C���}�$̼�.fXv���������ս-r�J'����3rl���M��K*ey��X�#)ejR��cS��ί_�q_��7'���$��i�'�3l>Z�1��$Y�ͯ��������G�Ao���|����M_'��K�ʖ��̦����Ș�7���h������Ûc?AZCOO�K��̀ ��%a��6vvz-f�q��F��y1B���"hhF�@^W� �t���#~VH�w������oIU}ܸ�B	&6�퇢���,��Ć*I��.�L9k���Ё�� 
�_L��\�9Z��\�^0��0�3{����B��M�	53���]�v�'����{J_�����
�3$l&�d�γ�^5���;ԩ=yXه1g���.i�����W#��&ߺR�f
��=�#�����S��hS��:(�c�z����k|���p�$F[�\�8��7L��Zg$$��T%�;���!2��(m��a���iA����o�zqk:*�I3RQ�f�I�0�>䳆�zY�Ȱ��Y�C�O��>�]?= �[�3�ܐ�(rl;����~���z�n�A�n+|���`b�� � ��?M2Y�_"�7Ra3��&�dr٥a�]g��h�[znJJJ����7MO��TJm.����h�$������e��@H{��[S��\�\�8���l�̂��wl:]��Uu�__�9CJ\�}����.�9�)�f�ŏ.&&E�Z���]��]��?*�0AK��+\z\���E��a�0n��1�����X�ǖ� )7��rC��������(�fLH�'�-w�M2��
�,Ѩ�.뻬�'چ'�y��Xz±��L/>7��3�&ȷi�5����yʗ�4!����c�!4��z/7�O�V9��K�����߾�%�����2پQYI�ׂ�g+�b�lr��/�#K��v"~��*$���i%�3%�*t:�[���Y�\�݆U���ָJ�BrD�\b=N#��b|�Iz'�"�τl�I}vXfIm Qo�pL
ҡ��@BBC9Z[oC�u?��7/Ê}�~��~��v^�?��&��ς%�;�F����a���/޴-\ʇX�5��a���ӧʚ�߷��u:���ݝ�'���� 8���W�^��Mq�δ�	�NnN.0X�WOYr����d#q0q��'6��|-d.����>�U����8<L�E1�[_wFǔLjv�Js�Kܳ�w�����pn����<��V���7褓��F,������wl�sk��3��9��VT�\�u���smoQ%��W�~�;�v���ٳ}��u���hyغ�S�#��Ȑ,�8����F�[��.�jK][ډ�"��@�7��-f�ah�/%�h���斖������}�/���f�d	].�[�27Gb�8̡��I-���}�$��X���e�H'�2e�NY�m����1t����^IP�th��$[��~E��etzqw��RӿaMڸۜKJG�W��[�u����T"$����<z�V�)z�Ns@(�*�0Fr����f���s<AB��PQ|rr�t��f���+@�>��[�3)ʢ`�S�C�d��fOb������{�}}}���4ٺzo�����7�2��%�޷_�ɹd�����$��h��E��g�o�Q�/���?�X��H���u@)O�<���^m##cs��"ܶ���^�������]�-��w�8f7d$S�%J V+?��)}�vwۺ��V�,�Z�����G�~���>H�DS����زކ8H+�Y�!�r\�j�3� {�3@8�Gh�(m���m(p����Zʬ��ȩ�l�*�J?��Nac-Z/Ts�D<��s�=����0�\�۬Ө��ӯ3*��.��09�z$�\<|��0X�Ar�����\���z��t������*q����j�j8��� �D��s;a��C��S���\�����%����e�5i�5����h��ܱ���<^������E��.%�#m*��wɘ�0���p�-����f4���]m���*�HSj��k�����H��}��ZQa�v��%Q����*�k���=��d�)-��8�|xshI"c]kL�R4�0Q5��i��2�Wn�w��W0%kƦ��܂����sA���;������'�v��[���|�-�X��N#LRSAH�l� ӥ�VX�����7���Mޘ(�J�˪I<�=}:�5R���<��2�\Ğ�zU��V�<;�ڛ��4� C��uZ~�K���:4<��Ca
o� ��[Ty�6{�^�S��}�/��.*UW/�����0���Sew��~�D����/_^@z�)�Q#"#��_B�%:Q��p����_�nw���O�?.��&hr?�f����Ar?qa*0�Ї�|U���=M�"��?�E`N�����>�)�c��I\i_��V��oy���B͙['��_�T�#�G�+xM��g?�<eG*ϣy�5����e?��6���_t�݆���}�z�$�m�'���8���c�~��
}��n��#��q�z��ȅ��;{ꬭЍ/��WK�&�����(f�Pjd��ݣ��jk�l�
`'Ҝ�����J1z�K��x36r�/9k%l�ƅ	{��!5�Q���M!!a�V�Q�щR���V���1���d�E������%���Bf��$͢��K����F��5��������_�h5�,��Z]]嗕�

sp~��1�\���tИ"�n�=�Y{�!P�����&�OZ'���a�}\|� �@B���L��W��.���Ϊq�?1���c7]���LS6��,e��fMU={�L e��ڂ'��)���[p��#�hg9�h��z�0�W��ZWjL���`�����q�@���g+��V��5 �b��� �:�U� =�W�\��Od���Ba�h�ToǂD�IO�n�^�d�����{҉?b;�&O�	�3tz�uXh4����o�*9ss����� ؔ�������d��B3�T�6��-,��ѥ,��P`�+++_y��x����g�܈	[j�:>�I�}���)��������87'/��`ӭ���j Cǭy�z�EJ���2&,�"''>F�E�����}��m��R-���w��ӈA����ܕ
l����l�Fۖ�d�?�|�)C�_A�����?� v��ߢ�9Y
�����R�:���~�n۾Xl����gZ!՛��������e?Il/���i�����=
3�?}7���X�!F��b�ѥZ$4��Rk�OD=$�vи��U�}g��~����j��'���5B����V�b��h!]���򅅅2����R0�:�������F�J�nάp�y�@�7��̉���G���L];��/~�EײEu"Ve9�@C�!#'�3�E	�C�Z)A�d�����8���Mq�d�q�c&ܚ�#���a�����>�0�� |�x��4�o��a�A0`�eD������u�
�܌>.�ԉi~_o�����v�AL,	�'4��F�[���l�
Lj�X6E.�T�@h���� $
��n9��3����(���#Xy��I^(��,��������3�E��d����;6~�K�k��P&�����p�[� �J��m	�/E��NOk�n����
�c0S�i�m=�b(��!������t~ʶ.���eo�)��sj$���R�p���e}O��Q�����M?P%�ՎK����e�4lrx���N{ڀf��)����#�l���fY!���&���T$��X(��Jb���R�(F���yf��x�b?�غzZ'����F=d�=pi,}���@j^C�L})S,� ��5���bhG'<�u��Q��#��п������~R�-]ː�{�:��F��^��'C�B������ͦ�-J���y�,����&�6�D�����?�jc�΃�.�F�B�҂���^g�v��S
:��F���3Ј���"t�55�띌��<e@醆Ry廫�����f
j�Ʀҭ���-�T�{����#��WؠSjDDDeHHH꿡L���뻱�T����5f���-"w!��W�I@�J4`��O��Q=c�%D�k���WV��k�Bb�(����˃��=E�8�K
�f���
�S�q��-I*��l_����ȹ�t�![����q�~�P\_na\�Cqe
ԍ����! :�_?]M�ȭ?� ��n���?	D2w����l��,m���]JP���i]��2lC�
V�V�g���n}jr��]����"oh����Z�j�`�h"b�����f��Y��^a��i���͛7_E<�a��-�:�Կ���҅�x�u߶���-�������i۹DsWT���{Ci*���~3��U>x��" �2A�������V���7�R�.H��O�P�@�akx�F������ϼ/6¢��(�0�9�>�hx�?��ۃ��1絜t�����g>��_�ꗿ�?��!����@��i4���d|���lu��rRd�Y�uG�u�M�8À�ak���^Ӕ���_����]��M�;��p�A#PXj��xxZa#I���<�.������Ic��w��rr�i�G�v#|9�̜v*ފm5��L�*�׏�{f/�J !|����|�	��-�����>u��緉�22&���*E��%X^-����'�=�Ė�4��e����}�IIIi{����k�f>56BF����m����Af��kl����U��O���4����?�y���cIe%�\�ch��s`b���X�>����;�u�t<S��yg�TX�*e�-����1�(�Q�z�k5��l~ҲEQ�j}�,��GR��S���Rv���J�W{����J������Q�S}�S��쀈*��-[�x.%�Q �v ��;���/%s�����8�@[���:�M����"�Y��6�Mp�"^IG�V����k�n�'���t.�����%F���42P��KH<�M���`�$H�
l�����>��ҳ�H�qf�+#��Ֆ����@�:�����"���Pa> ��)�h44�\b��^qp�ZYկ��/HflV�R������`�#l���1@Q�ۜ���7c����L���9�&a��\���^�w���g��L{iQ�K��A]�E#��3ϼy��U�y�v���<=��:s�Qr�(
�6Zä�.�O�Z >V5̊������ ��}f��N�♏�"���k�)'���\��lH�R�!-ok��@t�����D�ݢ���D����eC�j,�<h
�)L���5\y)�Ho���b�\/	���Þ�e`c�
D�!J_qc��洣3�oA"c���@UZZڗ�����rI��Q��Ԛ�K���dx<CG��Ɵ����������}�b�� ����OKG�v^�7�ncgםĦ;<�GN�2���W@�z[�y�|:+[MZ���36�h��~�E�=rWE��c׶0�dS�NI7���qkrb�)~�BS���w���ޤ���0ӎi>�B��Q���0��1�;ie���2��S��Ӽ@�A�,F�Hz�ΠU���$5���gЌ�($&u�����^x���0�kNi�8�4%�05���s�/��1�����%��ߘ�9RzȖ��r��wf�dN`���A�$ � $����c����w�L�l����_�c��ǟ���ή�@麰/����z#���-:::�rYjF4�%c#f׻�dg?�B����&��J��)p ۰�:;T#�o�v5I�Z��hO܀���������'T���c[&������Is{����g���4�ǘ�7[]��EP����uj�|�E��K�}���U�3_����͠y$�Y(J&8<G�smpQ$8~��">Q�v�D�t(�g��11b�����'��G��� 1x]\�}����A�N�Y�fx8�`�Q
��������UG��tk�sh��P���L���I>zq������H�9�8#��: �b n�=��*u��ߣ��Y_2|���H�p�v ��WG� �Q �����_�i���B4�$��mfwoo[_V�#��Wu�B2�!=���S��Q��j��a�#���9\G�wYfH�����]������/�+��%��Z6Q'���S*l���I���h�V�[(�˻W��[H�H�_�ی��QkSyy9y(���"�]�Ӄ֯��ՑϞ�K�}W�&u/qQtvsg�분)�r ���F
�/@��9�P�&��L�Ǟ��`�[�s8@.۵�� y�tdJ��<e͊W4���:��-@���l����r��lM��q��]�ީ����� ~�.��b?c�յ���rJh:$	��'��y:�&"B���,"L�M�0��=��=�gl#^�(uv��XSQ�����X�s|��S[�	wo4���c��X/�*؇2Zbw��9�f�2B5���[�/E�}�8e���+���������}������E:���f���4��.��/Q[�4֭�����C�9E�����K�ab�2H#=H-⇨B�h ��	6�g��1V�V�['\@*4L]ӑ���r�7�j�\ՀT�NGj�O��&@���k����i�'?�Z���B�{��=e�|��YV�[�	П�`SF�GBqoò��i�jk/��*�����@��礤��zzzԉ�/!����j"�uo��#kO�����
������911�X\R���;{Dvи[�����2''��xa��.��EW������7�hx3%�����!x@(�r�j@���j��J��ZT]FG�Fi�t���/w�b�i~��O*�����Jw�=�hG{����Y�Ͻ�u/��u_	���"�L��ފ��oz���J����O�����:�<��{x����7�Sō�-���&
�Z�>���3d!.�\�&�5̯`���o�lS�6�E��0�PI�v/Id�D��4�cϗEId����u��sf�m�*&J�Z$�oP��k�|{NFv���'������ zn!���"vc��GK��,�s.`Lp�V��g��Mp'�hxy�ⷶ�� �яFH@�L��
3��H�=�� 7���e��dL��o-H���K�DIT�=k$h�h�L�������I�ys1J i�{��f�������8�������L�`d`iMxԗ�+-�����1���	�`ʴ8���.�T� -꯰r��Y�ܻ,4QN�_���=p"l�������z��8�E8�Z�,
�r~i���I�'�����;���ˁO��*;j�eї�^Z8���	���}�-�L�<�D����a#�f`oE�;�������GDȫ%p"���f�؛A�c��X���3����� Ӆ����	�AJ���h������"��ww߾|��9b<k���ߛ�� $\��2�5��I�T�&4�)��׸��/�ß��1�d�ќ���?3�n�fN��gU�<����_}A�*��y�3�<�	k۸�׋�첈���{�v�b��џ�Fw�"�EY[l20��t��.�Ms���N3���$���Գ���Y�/1U�1 }1�gl=	�汩�s_�EjKEF��H_�p].�k��_��/��VC��#9�G����?wbH���.G&���"[MD^_?=��p�+((hj�Ϸ.��Pr�P>��sP��@4\#�X�+(�fd`�v�@z��qfgfFh��w�&H��v����]���?sc���`���������NYi���*�J-Vx-���H�k�NF�]��E㈊�*L>u'/|ӟ����'�4Y�z��n�4ޚ$���I�����3偀�}Gʰ}.*  P��� �����+���p���|H<%Q���d��Ha5��"�s�C�F�fX�	��-ݓ�^�#*��=���m�jA{B���a���������MC�_mD��F�Ksma4$�k�Rnd���A�Ń%p�d���F�Gw�����q�Eq�?�_�Eu����hZ/F��W{��-*e׋=m33��q͛:Iz �츸�@[t)�"d�&)ݚ�=O���-�X�8���<���Z�F�MIM�0�����B��:k�l��'{��82�,�%��Ñ��Ri7���Ņ��+$��גr��ψ�/�'2>�/����VDQ�^���*b���
r�q|�6��![m� t�dhr�:��h���XKǏ ���B*��f� Δ:;<�͝�N�`
9�,�O�� ���N�?`��2zC��㊬Y�~�QȻ廙;}�?�$� .z�@,	��-��u䝆��$�w����"�i#9�Ej��888�J����8�-՟>=137w�g���
q?���1N�ߧv#www��Y�.[�V1��Bᇩ�$�o�������Y�����8]kO����P�[ʇ�Y�C\Pk�w��+�p�<�M��)��X�B�hv2M�l-m�7
�m���nnM4�9���X����^vC�v��o�VG��-�2=�:��	���K�_Ҿ$>�@*­��ÉY��ds�J{z�����5Е��v
(�f1r���?�<t;n���2Z�	���a��c�S��H��9*�8��_�v'�@���o1h+jh��� �ypL�PB���~�J~w���-2���D�s�k���>}j|wu��_�|QŌ���B��zY*w�=��S���Ժ�41x��� ��\��S򯮫��,
[2r_G؛�"P�#�m=�|�=�r �p��9Ą0�� ?:��5�'������m��cf���|�Ȟ٧���bGF��{K�
t'\���M$���23��2��H����2-4��(�9|�����|�F	`1���M���˼��~Wj[�W��k(A�f��f?[-!�a�bc�F�壸��?M��&�wO�+��\\.N�9��xT��_i�-���[��B����'8*LNZ�(� fӡı���OΞ !����
q������n�22��B��;�c��|��#��m��L�� �jj29��jjc�Ilk�3SF�F�����.QNd�\$����6<?`*l>�O&N�|͔`�+K����YH��p_�ݜ��ZddW1�M���$��~�猅��)[��y�����M�\�@1��� �: �9�O�wǓ�dCqM�A�h<nV�x� �x~����y��~e$�_�Ǔ�������ϼA��~�����]kl]�+ W9+��=���+���者��9�Q��i�,��h�w��ʾ<�����E¹&iu�������*ƛ�]ԧ�lV�rq*��KZ��ו��$��]�w�����y@ˆ]E�b��9mӬol��찺�
����A��n|jj�����F1�������)|�2��K;+��(��̄�5���O���%EhA�����s��l����;Y�+����lM��Ͷ�n�>fJ����|>ˁ|I2e����ݙ����3��?K��|߽����>[�O.o�k׎"�W�B��F'���0<9�*��)}����3�x�����-��i�'f�&1�sχFM[��������:��A���n��qx�)}�K�{�6���,�KE>����bps�kG�I���weҾy�?���($D���*�Xb����Y�?��Юc� �>�
�0D��GtJ.V���o��輷`��-�gA
�,�\7��ۀ2p�Q-���r�gd�����X�	��	RDs�j9����VY�%�9be����U<�}e}IrE���d��Ɛ�>�h*����:�/vB�z�����#�N�o���[Pr���OѳI��8RS�g����~{����A���G��G*/q��ُ�%�V ��=>�$w��8���_���\2�cO��G�:�q�Z��;�r�8�C+�����T^@��	�s�l�]I,����-R����_}���ܛ0�=9J��[��y��w)�N�f��L���3�M�=��F�r��d���8}����o+��Կ�i�M�Hb��M�c{���c .p������YYY��q~(�UZ�+��u��09<�*����϶�daS���CBB��������C�)�����.�����e���dQ^�_�����"  �g��m\D+��_�=���f��X���a��=��
/�,$����5��5��^�����^���ش�z�"����C	���2�Zj���7%�S�њ5x�BQ�vW,~Z쐍F)Y�՘���t��S!��d�{����]���e\Y�����D�B_n�����۠���+�]���U7�l�?U��%�{G12a7�������R�V��ϑ`���L�f�:�u1��&��o�94n3 ��FB�ѱC�P;�x�NSRRj�)��᧓fm���\gĳ�C��;�;99��{�J�ݞ��ߤ7���3[m�t�ď�?M��ШI8�V���uYY98�s����w�e��<��h��[�$�T�⭳��]yxxEz�/�ӧO�63s)c�R22(�-<T�{��^�Ō-#�ft-[�T�*L��ӂ��>環%�0�=�!�~]�~g�c�f���i�ܣbo��Hؕ���aiۛ��K�F~ k����G4ʲY-K�Rgvz�6�8��yN��	�+)us�͝�ö[�Ei�A_��>�Дh�q�1��r��[�S?wƩ(�.t�� �����]�^�8�'e���Č"j�I�uWLrD|�PÏ�D���$ �&8��B���৯~����oVI�K�j&ͱB��Ds7)�R� ~̸��ߟ"B¨��S�	�mXcB{{���$ߙ����<Z�t�1|�A���#��|,c�X�@9����od׆�H!x�r�.o���8W�[��J�	�> ��Ru�P+ޔE��R����u���m�`��h"B��-��R��� �%%k�D���&�Q�!j�3�����v�T���Pճ��l�$Ѽ�ZHL�h������.郾:�r.?��.�G��tw6��t"2_�B	��ow���ۜ�W~=�,�h��+���M�H������ĥ����`я�����p���i"���o�mo=���-�-�p�_�D�5j6�D5��f�})�,�} �Z��ߪԃ8�ی���2z�Ɵ����,Z@Ԫ���ҡ��Cn�tTb����8�G�H4~~~�@��.ќ�����8ۭ��Q�ۂhDdd�㒘 Es�aЎY���in��H��' ����4�P'0�!��Ws9��U�^q"A�����a�Â���"�B�U)Pg&@��D�W/|�(OX�Z@�ά�U&M�@Q�dR9o���K�8$eo��� �}��YK'���aP��U}�b�'y����L6������;!�v1�ݠC��t�^�R^����չ�JQi�g�:��=�'}�п��Pn�nB⧷����'���P����M��ʝ��Fy"g�De�9t��>�,� �I?��_��-���c�h�{�����-ܡ9A�kA�����l�E�U���Av�v(����� kp�/3?�A�`iaOѓ�����"�ǄK�d�"��&H���3��eϯ�+�U.�>�"�B�ܵ�t�J�.W�����C�b�WO���I�'�%��E;*Q2�?4�>�D눋�>�F���ES�G���H��*Ƀ�F���4�~&�(�.���;]�Hmǟ
�����,@�Ӹ>�Y�৻(9�.==�s��7�-%꽮%"�p"��ny��쏉��%��o�=�X�@�d�� �t�7ՠ�&�E�Tid���x��N�;dS�|;D)��8��9nf_%�'���7<�!:�/ �fp���2�0_�B/$�W�Y���مσz<�FK�'�B5�`�1�~�"Q �)�$a�8��Z��g��':%�0�X��;���+(H�`��F}�X����롗�����!z.<����Fp�,��w����jk��joA��za$6�^O��g�^�����G����ԦHhC�t�Q�'Y#���(.Zچ
>�/5Gﴣ��m�O��-6�q��W�E%�S�!�.s��Z(���N��?m��B�w��ڋ��%�j���/y%y��BTgH��ڶv���K�_�r�I����l5%�l��U��s���Jn��z�������6������{���#�ÿ�A>=C(,,TQSQʇ?��2�5�0�<Xt��^*�y�6�'�jE{��H������Y���\��T<�-�,c��zG�p����<�,D�x���ӎ��gu�R.���ٺ�$a����+��,�[�>H�,��<ӹ�`+�o�8�`(�	=Z�������4w�X��Z���B�ʨ��9u*���R�τ��4��<��5]KQ\������<�rQ����)؛������?�רp3.�Ӿk��=j6��t��j]U財��;�%l�u�t�w)�M�i��RS4/���$ɟ���X̶�Ø�J�$��O_�/�dA������T^�	���|�+\�����c9Bv?y�9��,�;�}�2-z���YxZ666 څ��~���r~m�ߒ��@��1�,S�#"�Y67~d�Ж���'�ߧ�:���0�L�d\�����iӖ�Z�ӹvtq����2�E������-��Ԥ�h�|Z �a'�3����Y�#+����*ֆg���B�G���*ݼ�,_Ms���u���n�5w�w}�tm|�����_D�kz�4\4=����JZ���`�_���C��$����$�P싃���K�����ފ�W��R�_#��z��nymln҉�REJ�Y[0cj_А���)���d0( 9������n%:H�o�~���3�>��x�륟���F3-��Ĵh�t�����/DXhI�29���l׾�cd &<�̱�3����P��W�Yﷰ�Ÿ��j�myu�Yr��Z\.��ĺ�Z~Uf%��D�T�����]o�����T�#}�����vH�|	���:u=��H��&�q��*���M�1�'tst���['�"<����я����x�]����qo���m4��`~��Zy����L�;�>����%�`�IPj�9n,N�ml��D:<�c��,��ڨ�>6�լ����y� *g� �,NQ�/���*Q���@m��R�N�M�8;J���m>��0}�W�3���!2nn������XT�F����sE���v0b�p�R�>���Κ�x(}�X���7�w��2��u��;��A鲰z;,F��F����j> n����%���o���}��N^��F��P�5��<]~{VG���kjF@i�1�ٍ?�bK��2���/*���A���$��@��	��Ѥ2J�?��#+޻����B�#s����JF{�<[�����]Z�p��qR�p�Y�p�3�dL'�G���^�m���7G��T2d*D8�"�~H���X��Mlֳ����_O��|�]s�ͨ]��V4������	�+�*Yn�!�q��`s�ѯ���h��ӭާTR��s*��>K	�k����p{y��?]��؟����|�a�/�@�uvJh�hv����p��J�ptZ��537?Fbǭ�q�bR�A����y�oT�ޙ &1�}�`?��M��W'��G:�ͬ��Ȉ6;��p#,"H��:{��O����Q-���<��!����8�8��^�ϻ��\��1�����<���V24V�bW�=^@���/9u���_	
�15:D^�,I�q�V0����ꨨ���AQ)I	�����T���DABZ�[@D$��n��x������t�q������8����,���VՓ�%>?#j���f�wW���gz�?���ܒ�Q�%)S����I4p���g���Y�8)���z��M�5�*��[1����t��ӕ<�qG����ɡ��Ɔ�����<ڛ7w#�Eԕ��A���B�8����N(�*��z����~��R�Yn6H����:��Ɗ�b�'�	fo@`���3�C�X�'ƀ�d�r�c��09{
���m�Ņ���g�L"5���4��F��\J������LcH�RD��<Jz��Y���+���a�Q�>Ɍ�s�v .��]F2�䔥���=�9�MLđn��[�W�Y��u�/IZ��7����ܝ)�$���g����V�q�C�w^�Ȕ����`ëB����&��)n�3A[�;a%qڈRΆ�����_R�3��ӏii}dc"�Ԓ����ev�bC��@�)(Ȗ���$���P<����M���0k�j_K(w���2�8�G O;�O��Ut8��U�|-b(���������]_��~s�����dm� �u�3�);���`�n��~����`����##GMMa����&�fP6ٴ�z���4>�C�6��o�q��Ȼ񒯗q,�@��Ri�q��"�s'�����l0d!��!沅��*;�T�ę�t�t��Zf��[p�3���P������b�xxw�%��7������e��@g�|=c府�@?�N�������}��*;�v*-5��Y�o�.�#Ra)���q�����у~mzb��|�8T�{����#��:)	��6{i�ƀ7� �#���(Bʱ[Uuik�3%ẍ́���c�)�q?��p�0�c-�a���!�3����g��k�P8C�B���eC��-���RE�58�����q��ʓ��c���'��(
>�̝A\"���@.��^�4bm͔6��nԎ-<��n�&�䟺��A�"�G/���.ICq=)ᙢЧT�M\;}E��x��+ؠ&L�|}u>�n���#���v<V*D�N	6_��?�i	K���"�1����5���J���'K~T]!�׾���[}�ر~yz>���8 ��8a��V+M���;Wơ�`�U*)�ZJ@v9�K���E/��(F����q��߷"[��/k�̲U<��k|`��س58ʕ���+o��>��\�@G�$��f�;^ցR���_r�}W�*�Q�K%��v�Fww�}<<?_X�h����.���T�I��3s�(Kt|dm��a=u�Q���x������L|����"�k3�&b���U�F󡷣l��î�2������",���3��ln^����K�/�Φ�,C
�`?8kwՉ����~�g�̽�Q"�^��%<&�d��u3-�L�h*���<��U��o�@���i�r�%���:� �^�����4���9�f5!�L�|Q��l�-�O�Zr�y]{+s�ߠ5��"Lj��a=I��<<O��/��T�� ���D"�65��JK;��?&$�I��y�R1n��������J쩣z�G����m1��r�I$0L����Y���̺�=���+��d$�A |у���-��*""�l?��`[��X0d��j?(iw^[yn'P����)u�_v��UX��u�����6O	�5�]�����������	��Esu����^q�2�'3O��+A~�*lGԳh�9%���4�?��R�$����FJ�#�a�>ߔ�U��L
��#/*�~�pn�3I|,,�2�--�G��9_�ES���ݷ)j��Ds���gTÍ�[��v��x��:���T�@�k6R�Xϣ�Q��%&����]�hʲ7�(�!N!���N�z��=�������x:!����v�Q��C֝m�<���|Th��l�wkw����;����n��G SA�]��}^�.Ш����-L�����A�0��!�ى��S�z�oEruT��;g��װ)�?��)f9Y}��e�C�)A��qbbb�ϵ7�*�N�Q�����������$�ת��k�H%]�F�j��&/Skk�7����X��PX��l�0(Ƹ��^���^�W��p�i)�ܢǖ˭;�2�&�vߘ2�K���9~�8h���JF؍�>N`gWV��['���6M p.ۨ�
�ZT�$l���q�멉dm�[�!5��s�vME��M���b��ɡ[�Tp������X�Wҹ,���,�i�;3���T�C����e�G�=���8~���HL�hA~~�H�6���_��Se���v;0^;r1SD�o�����f���K�n������NX��!,��UN��O�^{k��>�uT'��c��y��r�^d��w��;f/"�B�f�l)*�g��΂��[~�z��[_��Q�,F]��PԷ������5'=��e�N�M���y7�j�����p$zq��R�,�߲�iXG���	� ���/�ҡ�"�H��?(����Mt��*��/_:��߯U����A.�����Ee�g_a777	yyq'��5b���(���J��?V^r�u&���[7��m��o���Ӡ���`�{���~;�w��
S�r��ul�S�s����7+�÷�a�xt�t�n�(5��f�vx��.�{; ���*ϣ=G�}�~�#���&1-o�����o����9��x7���鷯e�p�_LceKQ��lw(�x/�Y�oߖ���`��1����5�z8�-6�Mߋ�$
��Xd�P��9u��hck8e-��n���ь��K#�w���G�ʧo�'h��{��%%�t�����Q`���*E���F�
f�Hrr@U�G�;��� _�b��֖�@+b�����p�>8Vi�+%%5���r�%��ʦmV��5e-�a�#a�p�lX/	%�ZT�������ie8m���ۼ5l��ƅ�d�[������o��	�ʘ��-���BTz�0���M_��f����if"]���h$p���oK]7y��*^D��ś�xE�E��x0���:����5��O�:"6>��6����߉,!	�n�D���`?6v�6�m,P�����Q^�'KS�����ЇJ���l���������[X��b�~�Z��E�D���y�����B]��m��9��/X�B��[���l����H���̢�
V�n{��R�R��̒j�1aI*1�<�d���ckw� �I�j�c"^�/�k����_JJ�ux���~�҈If��O���J�A� &�O9�<J2&�`�i�ܸ���-ѣ��U}r�w����Ty��<m��y-���]�gP&@6�>P'��劎�x2�^���C2���/��6M�ڏ��"��Ԁ�:f�%��p'�Z�@�Q�>#�u��#�Q����~!�i_��i�:C��E��51t3�2�o�/j�f�lx'�e�N�Y˒�}����i{���CSS�	K�|(O�3�w��*�
y�N��OM��k�~���z��a�ٓdJ+@_�0�ى =T�Z����tGd���ng#�LrVgA�����Wl��B�T�]�^;;s@]�=Q~�X~r��rX��I�zM��-��� (�uԄn�z�a����ù�MW�p��e'
w���ҽ)}LG'@���.�
 �2��\�=;h���)�U���?�z��"����i-)n<�=V5�%�a���ܐ?�'q{U>bVvh�H{�k���"�;�����W3���B"��t~��G���slg��{P��N�#  ���i�KLr#��䠤����S�۞�����P"�KbNNN`�+=I܎4���Ӿx���2�U9(��QPP�Q����`��R�5��i��\(yU��a����ߋ�w�6�����B���\������}~.��e�p�-�58x"&[1R�W��RPI���Ly�v�!2�nj�}�l�5F�07=J#T�\.Uכ��R��*���%=$���sM���iO8s>�Ѵ��������S#���F�6w���{��q�6(��@�X���k4MMM�*��ܖ����L

��"�����&�~>�
�1n�W�-s?2&%�͙�":b��_�r�L?�I}�b�>���~Q�3�v``���F�E��t&Y8��1^��	��D�!���g+2×�U�n]]M��j�A%X<�v��^{xEw��&>��5=��1��BLd��Y�O�[��@I��ӈ �C���fI��?~�n3��_5`��M����d�^#���vF$����!'V�[���쌸Zz���X&&qKw,CTJJ�e��T�===\j�Z�8-�B�DD����p5"����;	_�@�z�0z�~�`�A��)[X��?��$����^�bD��QѦ��X�\��J�TQ2[e��F滗�G�ܳ}Z����g�i6r{c;���\UG^�L�0:��IT��l��o� ���}�2������>S+�.ʲwE�$�!\@0o0����6/�v���)�'�c6�O�z��17��餅��L�ފm�%d����CEš�{��h�*��f����1]v"g��K��j�$r���/��e��"
z]6��&i��JCi}A�T�Z� �u�D�ah�}���|G1������%�vK�iߠr����cF��00r�8���M�Y�?_'*#�2_K�jG���S��&��q��[�DC�m6�U1��/�����JYo��w<���3� ��������J����u�v�C6�.�(k�6f�"����|�C�!g���ǰ��O8��W���3�qc$a�Q�<q�����0�N#�o�㙮��|6Q�}�k�b���f��Q�ר%ϻ�:�>�j(4`�[Xx=+>u�WH��d-Ȗ����K��������o��6P�?��PUR��:Hs?_�U��*�����=}p���u?$��e5�^C��~ ]�^D3�nDCt�ӱ�H�@���zY�J�o��0�����}���I�!�Ϭ�q�Zܦ
T�)���&5;֤�+������z�Nr����G擔�
�(=$l����7���VWQ!����ٲ)8��M����a\5�AUfV�co&�.-P��lQ�h�������X��w�,���������*�E���j-��7�V
iZZ����rY����6���ݻ��xߙϡF��E\x�Ul��D�`*�I���SrV���YVb��T�G=d���%��:��xÖ�F$�0���1mZ�u�v�8S�	�-[��c���ԝ�\��SЍ���U���J�X��|�DG��bS�k�u����P�\dǬ޳t}@Vg=f�7�Q�7�Ф���q�T���tzAȵ��g�Jh.�)Q��y?�"*ؓ?����n)�L��%%{���3�뵟?����Xm3˔��Q��C�1�f��N��o'�iboik�%����'�an>9s����n稈\��w<Y"���F��	!��l.��Wg�C(�򜒅ٶuK�:Jbh'�X�3�ޅ�$�+?Ϳ+64�͜8�G+U����x���i������Y7��EP*s9եz��M���l쪚n�\�o%��=�@Oy���Ҧ��EC'C�����RQ��xLRL�e�ӋL�!s0yD��*�\�\���-Ӷr�`�����u�aH���,ӧ��^U[��GUU#�lB��=|M6"U/��j��'�H~E���t�����[Io����� ��3e+(*zѽ}�����j���OUuu{Љ_g��{ނ'~�sIS��J�L������DfXEQ&v�-mA7Q�Y7�@Lگ���}��ݟ��'�e*�m"�� ��o�̊
���^G����_����7�����_T#и���k���kQ(��i��w�z:��$����]���hq�j�j~�C�(^N�!�7Í��vx�q`!��/��T��[%�_?T�����rP��r��q�E�l)`�ƍ�5)),���ЗA�)�o֫w�RRV��!w�r�NX�C9VP[AA���jltt4��oB�T^��2;�Ah��?����}��I�N�]#(KS�����X�/C�z�źd�e��P)��#�]��{V�_�`nƣ��u↤�ݙ�����u9���N^�wihZ}�����NӹreP��k�A�BE2�{e9��DkfB�7=�/�Ӿ
j(e�|/���l�v���2ő��KT8q���gS]kX�>3�����g�X9L#�/+��C_�\e�5��!��EH9WNUH�ω[AZ:���[�nu5���'�7t�%�_�]]]D�Բ�Y�J�.y������ T���XAg�����ݜW�U�i�coG�H67!_��v»?J�Q���hM�e~I������{�˂"��>�~�=g�H��j��Fas����1`a��,N�
T�7�P!	}3��]���b&1�Y���sם���]�Ɏ����8�����JCNIzr��ȕ��j_9Wf����������x��8#�C��tԮ�d��ǰo��Ǚ���2��$4�����
k�j�Ԣ���Y8%QD��I!<###s�e{.�[.��ӡ/gUQS����}y�A&дӺeo7����:1�5<2�����I���O�Jw
��3�[�Z�,M�)��=6ֶ]V!C���+��?��Ӟ[J�n�G>�gS�=6e�^w�=��͑��Gi!C�6�s�G��W4�6�J3��*�tF���d-F&}�����;%�U�J}�3XTiS��a@8y5V3<�cH�H��Uy����ƽz��j]#-���6�u2�FƂB���ק�j��چ9��d��jj�X���ӟ)~r����T�xO����˫��S���^`��M����h��r9g=?a����b����e���cP[㽮��~��$|���1��Hv�%LO?��}��A0T�Y��ьs�5�*y#�'�,����$�`��#�(}���gSV�z�ޙ��Y�n�H����on��7b�Tj��}��S���dy�t��9�g��`?m
�+�+�@u�S20��˩�Iސ�jaYޣZ�|�})ǃd}�B^gD����j��}4 č���1
�/Jq�;���o�^,��ri�'�
 b7�	�I���{�Y\,�W�~��=sSS0�wqM`0�-�+=vu��]0d<�<-Z>�wQ��.9�����y�=^��vC�0�zp�/�F�iφ>�V&s5���`m��V#��Qj��A����3��M�g��M8��_�Ṡ�9�PO���~��-�Ƹp1ʉ��ҍ$٧ �z�ۼA����7 ]]֨�i�?����SW���r=�Gn����<�d\�ڊ�1=;��c��r"������=V.lffFOO����u����yͤ	�u@�v�����R�Ƿo��9��x�i�\;:&5uFݙ��oo���! ���Gy�x(��Aj�`\r�g�bK�R�X%;��B�����=zgd��W��I� ����If�^��&����H�fw�xs��d�s�>8�����HOe>�^:)%!����0���l���IC�B�Þ�u�94*ʫɣ�ӌG�k�Z��i ,2"�o��&e���j�sw���ui�SM�9��T�^Yw8����F���n�V�xJw�\�#ia�!��֪**y�����c��GG����P�����{����k����{8'�`�I\RXXh�VO��K
Y���ZzZZ99���~L\��S�� Uhiie��=:��?Cy�~�4�Ӣ"Y�m��a=W�w�˥D%�Õt���3k�T|����_Y���ϊ��|����N��0���N�Ź>y��#��6��@L�f�s$!f��ݵ���/��U�s6gk�*Xs��i6��HyN�/�V�*?���|��J���s$o^�:�)�&б��kE������:y�]{��~��'=���\�Q|=��P*=�(ET�h9��z��/_A-��k�(Ű���MU��� +��srϮH�'�+Ԓ�'�|��w�����"���B��,����]IM-n`pp��i��p:����;��uuĎ|�a0�w;�'�@����V��#Ot����N~�:�co1�T ��v�y��6o#	��2�����Yh�>�HƤڸ��g��~ k�߭8���օ�h�y=ޥd襃��8q��@���*���)�gDuM�gǵu++4�GZ�f;�hhM�B]TX+����;�d\
�dʹk�6���nojv�R�v�O�S�?�3��QT�����h0''�|�dUUU�|���$A���ԁ(VTV^�;tu�iG޻y���F]\<HK[{@��6���+��;i0Ln��}�߆.��uv*�����~�
}-;;�j~~>p�/{��f�ߺ����\�بkee养
�[.�<ј=q�m���������/G�w%⭹�P��M�5Q�/l�X��#�J/�v���,=9R��ib��!�ŏ0�0�U��JY"�ԯW1y�d�>��r���~�A�}}� KQ����Y�'�Qf�*� ��`�U�LN{�i,TN�IkUH�2�����vzb�	&�D�ț�$'k囿u���M*��P�$�@�a-o�曌ʯ�:�̣�W�^�� 5���t�ӌsxuU������`+�����������ϕi�����џ>-;�_�U��"�/=0�]��(��HK6N�d��o��;�)AK�<��C?$�����J?���x��7�Y�9���`�7�2���k��T��:!���p!Q	I�U�h����~r��=ǵp�GJ���%��C��%TE�5�/S�=�|Z��e�s;Ҧ�Hr��̇-=�#�; ��T�=St;�Z5�w6���M�}ֻb/	p�=��1���FryA�eGr�b%�57`�������mq�����^�����h���I#ř�e�Z��J��YT���h�ݛ7�P܏�n���͚y��B����z	c��=r�z��	���������<a��'�;��?os�-Ey	��K>�o�L�K���K����}j����s����}jR�#��ӕ������7{��0!�|Y�����:,��8���!��0���$�)��'�2+7�V^��O�n��%If��� 3���,0j0TtlBƅ�c:ӷ}��?J�$��%���je����Plll(� ��:��.����:��������kЦ�u�U�k���-��ۓ�����C
 �Z��"ľn�O�s�~�^�2�pӼ
�O�L�ی�Ì�"����F�1�m9��洳�j��&�)��o����[3���D�[�gՒ�i��9|+�k�%�@l�OcM�j^۔n;����3 L��k��F"?U� �ί�@w���Zyv�L�蝖x��2�g`p��:�~(q@M=ë�Ǆ]��*�܅ׄ$S޾B��yC��o�`�)���`��Kr�ժ'��_�U"�ȅ�J{��;�����@��/%� "��X����߅~���1���C�hħ�{Tz��9p�ӳ��ԫ��v�E2�����^����O�E�T�1�g:�8P	:QQ��՝$�����χ���ᆒ휮�#����M|��4;�P��ql��� Jߊ�1����ŴK���Z��W�0�5�Q�A��U�YS��H/�(�?p,��8��;�c�95�u���4���0t����W��E3��Vc�1�Vw$�k>��6%�m�u�t�*@�h;�I襖ʮ�v��XdC�Y�� YlQRV7�W�Cw5u;9-�'�@u������+]F���T�]���.�g�/�9`{�][^.E�C'�֟n�`���eJ(x�5��my�K=��4�T���	G�k��Fi�QtX���nLttօ�7�q���s��ɼ�f��G�D�ꂅ��"��6~u/�忲�u~�|��������� ��'�5���K�F
�����F��S��)��5Yf�0�P�ȦQ[K�<���h��a��3���~@7�)hI�
j�DMq�����	�K#�(���^֖���R��{���I�Y���}K V��+7\��:cMe-��(�����p�N��Y~׈�d���$�E�a�*z0��SnFT���@¯܍J2��K-�O� Y,E�k�x���x&aK0���׃4Z|, �F���x#/��y�_.cʣ�:yc���zT.Y�����ʧ��+W�{��g?�Y�6�p����޺�%�X<]A察��gT�Q9���3�.��W=�6lI�<o��`�[qc����:��f�K\P�����#�S���ėYl�gF ��	nR��M���ɷ�m5Z�r�o��r�Ef�@�6�ֽ���Z{m��2r{�WV����ڊ��| "��o��e�K4#���6�V�˝�c�r����B&ԃ���vP�����@)�h�#���n�r� �p/��9��w����O.���Ύ�M��#/��r�d#�-����ΡB�L�}���D4� ����R ds�އ>�7Rz��03B���Z��U����3Sl���1�$ŊD<zhp{p&���\2���[�v�G*]�uϔZO��*}�Y�8NJ9H���ў��y
ľ�����{GE��S��k�~eL�̈���0�L��i�(��.�V�I��0���h���6� 	�����.V�⵭YܼR��=^�8`f�z;���\��N[���,��p�Ü����B�]�����2D�S_�E�?�6P/<npM��6/��a���zU0D`b�'vͦ`�Ѭ�3|~��U��T�������KM��C0��b��ݟ Ȁ�iU�+=�,l(�%�w�����d�Ms�rtl�4�Ga;i���#�R'�4yǉ��j�����ju@M~���H�֬��`�U�z�h�P��W#V��Wr����}�~"|��yA�-EŮj��S��oj����9�����i��M6d~K�6�g+��>}X��Ț�J�o�zw[���p�ЦHBP���68M�:�������dc0�뉳���;�7�f
���y�_3�6Z���;�xA�$�?�"W9�HB��廇��Zk��"�� �r"߅����AAK�vjQ:����?���/v�IJ�Q�����j���R��辕Pb�J�?X	�J�&&���k��q�6�3s��l���/�i�+«�.�{�x��b:��=���y�)[�J��n�%�@���Z��R�w�Ǯ7�7L_��I�+�9m*f��7nh�+Ι���d�Q��l��G�Fg./pE�����l?^f��$���M2���F��Gb�rIS�T��Z���� @y�{��mݐg^�h6���M�=�`����yI�u�h��n�4�l9��h�����V��x��ba��Z��:�V�f_�����c��p{�y�Z>�Z/���Uj�>�Q+=v?[�V}r\�@���"
�Ҵs?տ[$�,�	c��~�+��ٱ�|y�WD	������`����<��:)��f����?Y�>3�����S��9asuƄ�!j�s����`��m[�>$���ю��u/JV n|��p6?���j��0Q�8f_ߞT���2l��.�7�@9d�V\�>��g	�9! �-x�eo�Ւ��P��v�Ϥ�L��cu�����hH��x��7��J�Z�/�_�/��v��Kth�{�%�f�<�H8�4�zgů�H���T�3�J����I/7+@ 5� �b�t���y��4�p���R�pU�#����10xAt�pI��Ҧ� iB���F�x�$�n����H����&4��������Dg����E�f�l
.�:}��\yۖ0�F�e�>2�J_*5/FQ�@i�&�QX�[�沩��'�}5��U�I���![Gu{��������&��l�������V!�qu]c��A�3�\����LM�s��|�~毚��;װJ��LtT�����^ UQ
��Kv-N�kX�\����f�� CC���U�ݧ��=���tQ'IMr�P�;$��oE��!7��#�h4�kP!]�R�/��� �b�k���D	i�6^����9	u�r�ʜq2DLpz?�~% k���,��j�]�����utc�	.�x�[g�v�4z��w�ˬQ�t���5�t�$(FAk�׼����8�7���t���̘b魎�� ��,Op���IdmDtoO�9�����O�FJ��[��<I�T蜗�.b����5�S�Z3�C�C�>Zj$���H �Ԣ9��E�����O�J�K���ԭ�b9��=,-Y!R�v�V�*��yb�3#m��Pr~���E$�������
�ʗ0,Px�` ��q�S4���W����T���;;w��4Ζ�6)�vt��U�]"�W�S�U}���S8��t�K���GK���>! �?w�9��k�����*��7�k?T����kIv�NH��x���*i4���2�J��I���|4R�����SJ��k���v��nt�U][�g�07e��Z�U��^�x�J*2�+#֯;A�)&g֕��{$�@0���ô�Ù����{%
�hg��)�J��$!ܸ�V�n���NחKͳ,;7��Re��?u\6: �3���j.,��
����A��X�7)��#��g ��;v�p�3_&3n�`s��1�,�nn�D�K��|,��8X ��|r�8FY��aj���Hq�)�$ĺWmڳ�B��6�*�=�	؀�>�������9$7�X`.`1�5�Ux�Ԕ��M���o�:�}�2� v�R/T�r����۸g��h H+���zV������	���uk��F�^(����Y� �N4�?���=@<��l*�ɧq���4z��F,lu�&�������i�]� ��C&�F�pT]���W4s�zZ��׸��q��N�v�lú���F���ʅ�W<���<D족f��[t�҈z��1��W�����%�7�S^�]���y=Y�և�ZsX��gl�K�7�-�{��Lt�gZ5�E 򳍍����h��Ϡ-��L�:f��s"��_�<����Ll�����8�ׅ>=0�5��"U�r�@�7^���aC��(t�K*y�Q�x��.��N �����E���j�@j�N��5�)�M&�@J�M����<3m���~������bbh�q��dQl��J��厡8���%�)�<�I<HՏ��������$Y8ϱg��r-�/�(&�
��~�L��gS�O
*$�+���eAd�����gc�zݺeP5�����)G$!���~��M.5��&G�I�5��{n���{>�\E�G!���U�U
�&�`�AR��-JOd�a�jh�$T����ב��厙f��"�+M�a��.����� ��WK�/�&�3�?�l˴�KQ@��]�tzMI� Cg kX���$�8.g�؜�R���-����D)=%��H*�QQQ��-� ���*YKO�[E�N\߹ůF6b�A�7��豹<���E\���t�(���y�Y�)U��j4,�)Ԯ�݂'ʰf��ĐVy��a������GO1�SC�!F��"P�������~��î�����'�k�5���_8���V"�/��:��9	���7T+5�a�.��5�W�z���e�� X���:�K%S*��$7���"aAab�����<�%+��"���s���*���m�G�iw"?�,<Pj��~�W#X��g+�Hym�"��;�&;jl��F�(�\�ҥVw���
�乻�z���8�������dҺ��TW�y��I������=�7��-pA�a�� y|���
'���=�<�=��Ap��$?���������e�!N▜ץG��wb�T�z��35���	��c.s��^>�@3��avG�(_�:�(�J����H�ǋ"��3t����S䃀�����K��} �
̠�}?ac7j��Pw��/�t��1�u�Z�x�&�8�0	ƗF�/%������M��J�U��jñ�Q`��M����l���黷�vԬ��'�>;~g�h�˛:~?me|�˴���̞�لN������&��{����K-�p������q��E`�Mє�ab/ ���0k&���.���s�	�9ТK�ȍ�� �N��v�nQ(ȞB����S1꿒�yAH�/���N�!�C�U��E˃�`�>�Ai`ńDx���<J�/�ږ�^1�f�<)i�l��`���J�o3�T��j*�0�S�z����hv��)G>U�/OK�C��$4�ǂT����9e;|G�sY�b�MY�N��"�G�eY��@�#?�����3�╲�鉍��p>@;�>�?e�y�A(� 6�hr����)9z܌�V����c9�����R;W����i���p�@C����I4�b-;cW��M>_�y@c�g�H�x�b�4oP��#ߎ�����{��Cf����Փ��?»`܎M"-G@���kT�ƌ�"��� 6���K"��ι�����lKQ�$M��������������L�Z�
g�c��1bC�Xڈ�ΘB�:S-��"�}���y� X@K����y$����SX��@�ēu�A�X�	Z�B��)�\���?��l��S�������3e_����Ú_mx����H)]d�T.s��D4B��ɗc9��< 6)��?�,]�ZP��l�
�y߸�m����A�� ̀��Gr0�a5���#[���4�?����qH��I��L�-#��Z%�a2�w\�%��*ۊ_{�~�TQ�h���pDa{ �H�U�R L� ������꿲�jS�uxq�:�ul�3n\ž����Ti�
^�d�4���&��밼'e?齸lK��2��CL�׭��dڦp� )IɁ��������Z3PK����D�5��Ŧ{ip��7��S|Vd�0 ���'EPa�<�e��b�����A�0�Q�Z�������҇�r�`���������N�vf�6U!2��7Y����DJ[?�ww�2� �{#��)K׼V�&�o�0�S��D�g�Z�nc֩4�b����~N���_�J�~����ߔ��V���dZ�g���x��Af�Ў�;Ku�j���"���ګ�2��̳6g�Y4���S�P��s�0��Ŕ������WLH�`Jnʁè����#棯�`C�W�6Z�Εgп
����1�sЗ�%��In�y[�^ǹU��O��P���FJO�R�[��O~�U���p�A���P����#F�:�`��+5O��f��g�᧑I�i��� �cIu��ۢ��W�/�ð�c�.[]6b����>، r���*�l�S	�]�
�4�;����]S]��G�{�b�ޗk�O�	��>'`��+�L�T�d�
,&�&����`�q%����I�`�eY��V�������Sq8��t�n��wu�J�B6���Ө|+	:+'�}��o9C/�{�U��cA �]2e�!���d�宝�_���lIU)��ܓn�4�>��/k%yr�,�I ԍ]U�J��.OJ��O����7�2;$�����,�R���\c���{Ū�~�MH �+y^)���h��8�6.}�'�ݼ�,�����f�i�����#��G����;�Hʦ�6����B��w�{8�q�Z+�(W�ڷ,�ð}Gas��t���(��
6D+o�㳢Ξ�-5p��o	�#� mܔX�.z�6Gh}Ʃ?���F�߽ٶ_�aن��O)�W���%�̈́���M�H�.I�'Oa��ɭ���߃)�q�֣�8�ttϧ_ ��R�3��C ���+b���zj���u/�A@���џ�y���ҡ�u��>�,!��X�b0��>j�q>�����';�q��{� �a�
L���W����D+ye��J�^�%�&dԲ����pE4R�#�l��L^�FE��	C��vg��O	����o�(���P������p������ �N�S���w�랇�)B����{�,����}[�4Ö>��y�]>��1�����=��K۟qd�Y2��R���i&㤅!���yǻj�ŏ5Mp͆�D��Ͽu�|���sL�Lβ*-����΃l����!)P?����<�O�kn���3>xL�)W�ɖy%-B�0�	��wF�H���2�3�.'�=���q@ގ�d��l���[${����h3G =Y�a����0�\�`�d��e����wMy[���(��k>�(r�|�J9&�����k%���S���/�]t/N�
�����ax$��X�[b/�E@x��q��y~�x���)k~l��K�H�j�IXϫ!k�Ay��_�b#R�B����嬡3'�`Δ$rO��� n	2�Սf��T7|Rp_�^�ț9�j����e	�)1�d�|���m� f�������7gI�K6��%��jC[&�|��[!/q�� �JC��+�M��mu����+��&���أG	��Yz����fɏQb����.|�M̬��}��6�R�͖�uڸ5��8�Xed��l�UKRҲ#�$�@� �<��h�fS;<�����	
^�j��L�Z.Br����#�U��;����5�XT�ޛP�)r�	��y�;qC0��e��̪6_G���[G�ǀ���Ӽ��VJv���U�s�j�^N�h~��u �V��{�>E�؞�{@]�g
�2�^���bN5��q)A��� �v(n�(�U���wO�I�sɸ',h�<_Yy9�e�^�`��h��r�.5k�g'!��i���#�xƈau����w���]#^�mI�9�Ȓ�}lZQ>�B�tu����H��H�_݇��ә�L��x����s��!$���X�|݆�Q��^�q�&��9QD���]0/��ff�<N��D�Y%� �'�W(2�#��^�b�>�����fh���ȗr�Z��ޓ�nu=k�߫����s����siP��|�/�˥��9���G�RȚ0���ѾL �s��=���eS����ۿ���>��|�D]�d+cy232�2�6�BV�^�Ql�[L���X�>N�C\*IV�<�@�_Gn�$�\�Ǥ������� �o�٧�����1������I�x�
�t�k��`ro�L[ʩR��C�)3��Su3zp6n�@G��$H)��U6x該Y:,gR���W���`�����@��G����).�����A$Qq1φ�J���B�A�keV��� �a��+���h4��Ie��9j��j��[r�}u����\+�D�x���>qFnO�J	@�s=�� ��x|[RNI-gu����wcw<~�iJ��Y4�?�4�`��dV<N���Ɗ�pw��&��Q-�y��i�x���q���������G%ݛd�fO��Z��zi9�z`�Wo���� �(�� �W�4�V��;���T���[D�����AAa��{��{���f�]K��g��~���w�K�L�5����k��g9* ..�Q-�즞'o ��2��>0�F5'��9��Y�.���������]��7_����?Xv�ށ��`hY�_��{�?�J�,���rL���y&t��s
�3��j��I�\iu��B�����2��Z9bBuk��G}3�L�a	=�Lـ���G�p���jo\��$|�>H�� o爩��� �����sH=T%��X��כ�w��z�01�>���{��<�j��!k�Lc?L1�.L�ʝ�J�)�<���zG�#�b��,{T �ssG���#�`^�sz��ҭ���{��-%�B���z�^3s��w/UzWpp�Ԇ����]�BpH���A�3q7���}S,E����q/zR���Qb�;Y����%oI���C����փǎI\"��j�{Tn�q�@	�ͳ��\K�m�T5�D'���Y���C�0���h��cU���^TF��i�[M��x&���a�����Ý�>�׬X�:nH�N�瞎����M��Q.����KV�{PdŃ/Ӹ	�5T��nߛ
��d#w�����������u�P�:@��b�6C^�-����;��?SJ9��_��M$�	1�5O«Ȝ!�I��ř�"w��6 �����6�>���*� X�,�hs%�� U�$��$���E] P:Ճ��T�FZ��+����4�,���>*�a�s���!4e�}'��ԿJ��Q`�A*�y>�6���%��7�"_@-�:�cJ
��f���1)�Y
#��������>��<�+3{y�o;�2>&����i���ս=
P`�-�3�qh�P� �i�R�V���Ǎ�:��wD��v�9��2���#wd���ڒ=���h&�b��Ёg�=�L�k'O��Z�)�� K�Y�dWxI�M!$_��x���c̔��_��Kc2�a���lˡ�?�ڒbԂ�u3\�X�M�j&[����+��S��ގl{�����u��骧��!N�-㷙���sN�{e��� �ڢ��7�dV��/Y����!'G �=��m?��V�<�J��Ӵ
<m���ω=�������!Eg�:v->}O�u��	2`�����ďI�5��u\�U���"���H��2�7[�A9�:�U���+�|�u�6�cVmb��o'j؞;�K��5����:S��ȃ�/�����^լ-�~z[Y�k�I��gV��} �{��8O� ��`?;�cI�9G1�����/&?�`�l4���W��f�-)��ZMf��^e�!�y�58DC�'q^S'��T\v3�0���B�Z�k;���x�y5�韼�DY}�V��2�j|�+�?�Z�:փ�?& �	@s��s����Ȍ Ypg ���,�f-$1aXaWs��1>�݄�$�-�����Lk9��r] |�#�f��sM�:gUo;\�
��3�0��������5�kҿœ8�� ��A���Mc��e'KdOFB�/���s�U��Ђ�v��j�	��ǾS;��?&��xཀྵ���#�x��[W���\�r��#���~a����贑gl�
��~#���
���r]�[Pt2b��57�F�W�fs��t��X������FR=~�n9rc��N�0��Z��]]/��S믤�u���㷭�jmltl{$��śH�m�����8�9g̃.P�N��>�ܓ3O� P��F��x� Ӣ뛐\Zrq�K����]^�lDP�ڹܨ���Y�Q��I��3lh6/��׼��	*��SV�%���S���t��1ۥoa����Izp#��^���M�RHV�l§S��hHxc�ໟW^v;�0��D?y�Q��m6�2�kf�Q��{$�/�!��0��(��Z�k?�m��;�p�V�=�x����% E�g�DP�S�fo$�)���b�}܀�ۨ��u����Y���x�Zj�4uAj�������d���Y��#'�6h�,�cݜ���$DU�/݁�>F�����R�q�����][��KW��s�5����$�VI���Уm[i���
XCa�/��U�mRL�&%�^�N��'�(;��>߅�#�d���j��v��_랻ל��P\zBjx%��=��a̹�;n
2�x��/t�A�Ң��z��̿}� �� �'r[ȸ"-��j��%+�TW�6B�׌�an�W�ٗ���'�x����e��M�/�p�N2u�&���) �3q�Z�!-/v��b9q)nxXW���Վ�s��X� ���������dT�Y��?��� ��¢��5�!�R����M�J�X>�
 �x=�Z;c�f�䍙�j��-��
�E3��Bm����S�!����ͧj��߰��.�zj�'�V���z{�#^&�b��d�>qȋ��㊩��L�ΛS>]�}�F�	� X�u��i�x*���VL��������-�`���4Ot�*.S�޹�,�@�eL���V��Q���v`����E���o��7)���!.�n`�� �5�Vw/Tb��m%�����S��u6{�
��k��2�~_鄏U�x�C��=��C������D3.Y����|q�p����E$y7?�C�d�F��W�����b�?��E9�BG�l�wJ|:M�����yT��[6̫C=�o޶,�����D��s���w.L��l Owٓ�Q�`��V�7E�}��_�DO�|��j��$JJ�Bh"��_?B�����؍��[+)���KR�60e�ڙ1r��)a������⧳���R�b�˸r�3�������Qm��CO
 �rk���F{�1�V�M]_go:����������������� 2l��Hy�e�\�9���|��H�X|!c�<kV��VN<��B�p�5��MpQC�e-ҽI]� C��.70 ���_���i?+6�����-���<��j�־�\G�;���Z'xgF�Ԣ��IK�����[}���F��ڐ".����r�A졉���h�}bYX�w���p�p]f��w$[}����1	��vWߣ��;ր*��k��+�����d(�w���V��ئ�X��Uq��i��8)b�}k�BY�L"��@38��0�3t(9��1<.e�u��ʛ�0��T^V�J��,I���v�����S��H����H
k��޵D�k�#Eǐ�Do8!<p�ũ���ٵT��/I,s#_&s���<����I�.l1��� �j/Cq�ֈ���-�/t�I��?�Xm/-^릭r�Koٮ���-C��W)�)�6�H�_l���hnq�=||���Ǘ�2S����,�e�J��-p���O����\��8US��Sv�_;���O,(^Z=i�=�}��b�����".d�jt�٪�[� ��	���������y����z�J��\���'Sa������;��\7��Ȱ_%!�t�w�B���O4SM�N�� �\��9��W�HV���OM���K�\��a��ė���x��pʆ![�%�:����?d����1< T��T4��3�)ۡn�P���>5�|^�p��@⬨�4������4�3�2�~��_�˯ztn��b�n�X�F��g�����K�<�8e�F򵓚<��b��鸿��*��9��5���+���M�L���l���ݖG��G,�h�������7��#��Pw;Q9��
:Z(k��ͻ()z��c�y���䝩�T� 7y,�_x�|J��קѺ�H�ݸ����6)	����hi�2b	�,,��Fԭ�NWx�^IwV�&����*��I�֐��V��DE�����ǒ�O�^�ޭ��i���Vɗ���L_��j��oy��׌�8�����k�K���JJЙuc�j� 9Q�O�V��0B��x,����lt(��j4�$���B@]�JԞ�v���y^�EW#S[�.uW�j�%\����p��\l՚/2.|��V�wf=֚� �eG��Aǖ����6�1x��ML��u%*Ѷ�)geVe�eQ�XF�%r0��K���zi��a7~��Ϫ����6̞���w� i�Frw�L~���(e�q�7|n_��[���ɡ���e���a�Hš��,]�Æpe��kjVT ��ӈ�Ǵ�Jd���x��|֊��uUuF�v�3���c���^N�Io��S3����=�G�����C� �����t������-�X�a�"�����B�������[<g˔F�Z�%�"��/	W�e��<�g=���O���)�˗bG��DL7V�i���G8���3�h&�����}*ɞӧs�]�ItA���,�����he�3~�r�>7����Z7��.o��Pm��j��UҪ�*Zp����O�Ӿ���y�v��cI64H�g�e`����F�LC�Փ
Êн"_]�W���I�j��4��j5(���}��S{��̙Tsl�����r�$�C=���+4�,RF%~�g����:,�uR�MHjҖL$�ڐOV��G�Z�76J���-�l�[e�c�l��f�j�����5ˉ\�[4<���y�t]��Ë5!�$r��ߥqw�
$��щ��]� �!y&�����Xl����V�B�ن�����;�B��\����yA����i��v�T��xGz�:�$@�(3�,���GV>w�FXk��� �瑮Y�-ѻ�B����ڶ�J���]F��k[��K��a%�t܍�B��D��,4"�r5��K�G�:k�P�cU������X:.�;O�ט
ڒ���a�����~<fbA��X[�w4��`���&Q�O���l����H.g��^5��?p�w=)��vU������}��*]t���_O�I����d7���VK�q��	G&�}�����eJ�3N�x[�Ζ�A�<fe��R�2���r�5�s�����d�-��DI�T6P袣JYբ��fIz�����r�rz(?�wE�������C�W v����l�W� �n��M&
����҅���Y%��>9�)��㮪�wx;g����ȷ��}�����a��M���ಊq/�����8���o�ļ�g��q5������^W�i�T�̆ њ*Y�Mp�?�x�aXb�3�ho:ju�=�C�ʲ}߬k�e�"7g��t�C�3�4��'Μ�)���Mo�鴡��7�@٭��u������l�f�C���mr��ӥeÚ���w&+��k;�7�yM6fn�O�_�4�i�/��_�1G����/�@w�xa�7���)�u��f��|G��y�%U�np�L�k+���~/ؿ���=3�8.;����+qI��a	ʻ��KQ��$��Z�1YM��}��×N2�u5O�L�_�ļ�J�w����-_�ua��$�\l(+�LT������+�cmQ�"�M0��ђ�1)��h;7�o���$�?�@�E@�4)����?	Ku�ϖ��Q��;�Z\ibW���sV{�)�C��`�X��M\	���zM���r^`��;Pkȴ'�r#W���).������5�'�T��\�7_��Wh�J7OGdK�Y�ȮᕨY��X9����	I�Z�aiSF�Rړ���]��s�F�&��B#t������k+xj�A\(l��>�JEe>K�w�DQ�����M�yo�������/Lk�֌���?����ؑM�Ԙ:]sӏۖ��Y�ܽN�E�����C���]�����G����\�
7�MǇ��,�8�ȟa���a�ݬrt�j�rJ�/�8)M5����C�=V�0�(��X���ߞ�.U"/V��tV�C��=��H׊�0�N"Bdsja0�+ETX���.�Q5i��°�v�ˋ��ߒSe_�\�g]Y妛M93��9��់`�B1Ӎ/])��|�+LT)�m����E(F�X�<f�B�c��KB����(���n>,!Ry��P�
�
dH���f�i�~R����d9X��A!'��*vR&д(&�Q��U�to*D�<+�<�W���)%�h%,����ܻ��}F#;���Ĥ� 	Uc���Y��Q�����@��Zv����usb���cw�b5�PW�Tz]X@#� ���r����T=��Z�,��j�9MF�}�+�xe��ӵc��/J��\�QW/�2_�l�c����U�+jXh �i�ݵ�����%l�vW5VN�zg��	���1��N6�? �
����P��dǲ���c�62���Q�F�X]B�|�F�G\-W�5�`�V��a5X�p�p'J�~�*�bإX�֔M	���{*D�-�Lߗ���5���i6��e������g��q��0%ɡ#\�����ٓj���F�Zl���U��f (y3�2'��Պ����_6\}�#�Nѡ�ϙy�F	Q4.t�Ӧ��Fp����c_bɗ��3K��k�ZЂ��o@�
s��^ۖb����e�K��H�0(��;�8������T�u�#/��޾HS��[�f���0��'բ\̓Sǿ:��ػ�M[��X/�O�Y}d�ٓ~��̕y?���C�bV�@>x�ι ���%��c�z�~A�>>O���Қ1�.忒�o����P}��Jl�{}ե�jp-����D Sx�C����>�t�U��`���z�Z�_�+��� �󪳩Be4��\��ol�|Oʞ�ܧz���/#f����K58��!Z��^ᤑ������~��h���K�@��υ���!�������˧��E$&}��FM��y�\�x3jnݲf~ej�V汀t-��>�}����P��M�77�S_7}�3* �ؕ�����7�q���v�/��H��%~7���ԅ�90�.n�:c�ds	VAM�L>Ɓ��Ŵ3����sunof}x=��J���1I)����+l0���"�O�P��/.�$�^5����<� ��ȳ���`��Ԧ./6��eL���i����ơ��.͔8�f!���x�Y�a�n�>�SFy�����N�������L�|��&��'���c_�6 �&�k1�pև���a�KⒶ��+�kr 8�*9t$�BP��^"@�)<�{>�������Q@Gɗ/�D����a�$ �y�Bs�A����ᯟ�-K�}&_E���������Hχ	_�n�q�'�B���B������濾]�\S���7v��(6,o�H-X�{�	t���͵�ؔ�t���d&���c�A� Jiͨ�ɗ*^�>��[yI1���4�D E'�����ڔ2Ta+�R�L���Kf����̣�4�1����nh?���a	\wF,v���8Bd�ˁq�y~׋�/ {�7�M!M�	,lJ�Ǽq����s��H�g����C�yx}1tMS@�.��!U��/W�ڃ"SR+hqh^;���/����ӕP�5GgE=���Ի`ݒ��v��t��"�c"�51OB�&`��/������йu����L�rxWΑ��/CgӄC����MX��i�%�?Xw��xj�w�j�t�-n��.	̒+/�Q.�'瑌E����o�
�Yq#�B��xy~�0�� yn�g΀�PQ���X�{��L7XT]R�e� ]:�E� ���ڞ�&�+���H3kVX����/�
��iBO �oS>&��><�rL%g�-�{�݄m
�n�7ۼ�4VK|&v�W������3��;0}����V�F��^����ӛ��i���7}0F0d�=_E&@��7ł�,]�]��lH��\Ј��(b��b��f�+��;w�Z��J�D��i�m$=��s̑Q�C���yh�}N��'�����c���C� | �	eA�����ε���tǖ���"�ڴ{]��V}��O#>Ȉ A*��x�U\Q�q���+������J�a�-����nғXuZf���스1Cmxh9�����jL@*�)�����&�(o^���5��4�U�:��DKu�g��`3{�Hf���q ~��B����|��P��*�rW��R�S>��O�k?���D�1~�v�������<!;�f�9x�^�nG��c��)�C�Q��e�P���|����T ?��m�h��$�|��s�ϒVkމ4�,�]�Eс_2=߷B�~뫄N熫~�c��*Jv;6E�;�Q��9ru�c�.i��DG�>�oJ�_	V�FҚ�3y �:�p�>�-��G�80X��)�>�\}}��r����jw�|����K ��7:'B�4�N��0��b���C��2�Es_$��Ze�
cO�f�:�;���Nl;9?K�1���Fs�l��>V-�!����L�a��,@,�vN���ɝ-�N���mcGF�\��r*X���n�[�<F�'�%-P�9��[[��[�@5Y��d�Ł]f���>ǵ���оB�����؇�%F^�t�&�)1]ܐM�*4Rw���X��t���S���S�#����?�o
����{����^��k���`�m-'�d��_
md�`RJ1�.<�<^���R@�Vm�vБ�1�!�F�#���M���uYN �E�����	����tj_1�:f�KS��iW�Α����_�BXN���A^1)+�ޅ-�?d��<����i�2T���)اί�����6��yR��7��3Z
�9�	�5x9i�J�8.@�d�L���|rʐ%�G����O��iZ���^a�0i�:|ްt��/*�;c��[�"tT ���/J�����Y�@H���+=�<ŨMm�@75aͅ��
�i
��M.`�SjSٚ�q��8�n����Zz����y�Ou�t�H��'�&�B��a���d%��A�5 E򿩿	1�N�Q]��ҕ�dͲ��<���{FV����22<("�\�hH��_�ȋ�L���.���,撿=d;�.U�&N�I�	��R���eTw������D��M�,���w��ĵp��[���/� ��-@Ҝ,���(d�r��>���mc;Kv�Q��3=�J�)@B�h6>��C�/l�a�OC�jpv_�J�A���?S��C�YC�:JP@���T;���2�~����s�0�S�+J�����֥�.wVU)�q�=���7w�1�Ώ7[��1a�Γ׎=a�<���g��!�V3k�c[��c�7�Y�;Ĩʦ�偩%̏�,����$���ԇ^FQ�$)yV���e�����g.��\h�V�߾���d�KS�.�i��w �X�lb!U�R�1l#��ݺQ�ݬ���=%����s�F��ܣ����s�F�P˔�k��=֬��ϭ6�G��4
�h��5��B���� ߔ.w�!�[X���MN�S���iG:�I�p��`�cn�݂$g0
���������5�$���E�$�&���D%��К拿s�& w���5*��j�-�K��J����G�RҒx���O���H�!$X�I��t��h/����}���k�fژ����)����Cc�i²���� �߯f�!ȵ���ݱ����]����Gj%�5:�ix�������gC����6.�dZ��~�x�2E.�T,��Uep���/7oH�!�tf��T9z�N�=/.L-���F��|x�he�i�ӎ�T��\rK��L�狳�5�M_ą�^$ؓ�.Gy���=/�W.,������w�������b�K�:�Ug&k�ok�Xfn�Y(��Ӳa����
��+c�X��:�6:w���p�E�b̢��w��Lŷq-fZ�vn�>J@��2@}�	�4m�Η�@�����;oD)�1Ԏ�O�P��?�ک�5Zd`�Y�-�K��������*a)RA١������:�o��=�O�3n��5�&�vh�ٕ<��-o��G#L��8 %sљT�Ցu*���z��O��+��(�r��Vq%�i��#p��f�_4�wn��� ��p�c�c&��:� AP( K9p�����a]�	�1a9#�ze&s�
!S��}��eP�����4T\\�jťƤ�>�Ǳ�b�,/-Hp@Z*�$�;�m$�����՗����j5�};�������u�F���[��4�lz�O��e�c����	�D � �^�l���jG?���!��+ݼ�z�R4���|$E*��@��W$U5*|󿭺�Ӣ�V��;/�NN��y")P�����dCԄ�*bF�����j��,-���8_�������^Yf�O����!��1�rX.�xo��'(Z��Bi��Z;�G"'޵R㺋&|��m,�I|QO�f2i(}쏕b<�oy_� ��@���i/��IPL�̥r��x%�)��k��U��R�]Ԝ��i4���b�e�@�ha(�}P%���CH,�\����J*v�.�
����4�j��Ƽ���4۳ϳWͨ�UĨ)Y��r�[W����0p�*���*��6be���@k��Ƌ��G��t��(8s�kզN6ן	��rW���jX�j������@�r+�^�qu��$y�����������i�UNm�GN�ú�E����F�ԕ�ǦC�T�v	Y�	�}�ݢ�і=�7F��?t���l�pk�g��<F��]O���v��> �N���@�-��|,T���:Ƀ-�4��w��a���/�v���J5����y�Lg���_?�,_d�d�VP�ü����ĮM-��LW!E����)B��#�Up�M�i9t����lI,-��k��T��t\92�g	0�i��*�dÃ�-ZU������FW{�;�%sX9j�腺����YR�>	o��m�9ɬ���E`�4e���(�x��%地`���G�!	\T9yv����!?�M]�������\{f�*Yj1�Ez���r���h[��&�$^��fG۱�y�Q���ǫ���xh��U1����X�Α�wm���7	�w,���ܧN�|E��Gy�s�2j�V6���/��kk��t�;C�6S�]���3G뺼i՝�T�j�.)����0�5�|B����Q)��y��V۫��H��ȾUZh+{]Z�Hǣ�T�R�\F<��t�I��M�흥��Y�;��XY�5��ۮ������yq��c���ZkX�K��<�5�]�n��� �$�`�G���Q	'�ms�=���H�S��*��p�!���c �Q��h��j���f���y�U�ֱ�;C��ڍm���V��jW�+����'ᵛL9�ڧQ���ŀpY?��[��
�o>>��un��7�c��>�]2/���LǗ��re��R�iRD��uk&���%��qY�s�&Y�����������%�<�����$�T��XM���l ��ګ	vړ⺸o���{T5�\.�6g�-�A�_��|��B� ش�h�'�Y��O�� SZƨ�@�M��f-.��[W����O���a�����2_F)�~}�����ܹĺ�b Yv������k�0���r��c;�vm�$��)������hn:E���xT�y� e,��?�[W�H��:M'����a�B������SH�{�.s�fEީ�IA�<�`z����ax��d\��%m[�KA_��m �pQ�>ƺ䓈H�D�:���R�|k�j)���YKk�ݨ�Z�Z F�+QpfGX��7�X�6v�9o�hP汍W�Vx&^�%}�f��-�<��>p���B.��?}pQ (B��kP��m^����B��x��!0�ѫ6�x��_�h�w��L��f����a<Jfl�~���w��ٲ@�1��z�!A��A��O�y��!��v(�"<�� �����c�̗�b�(��	:�c����}4��:u�Vĭ{O�%.PW�o����Xb
$:8t9,r5�;�L���P?��H��c��Ee��{c���T����"ڜq�,����敐���s�0�Bn����)��'����2�gk��>oV����B6��"?K�8�7�AY���Cא���S�nG�඘���V���^ѷXϴ��\Oq��RSb6��X���������)\�
}�Έ��r�����X1��/�����G��4w5�v8���k̜�`婛�Ƥ�����2��⼹$t1;�B8)T᪷�]��6gE|F�� ͂���G�k �$D�TE���X�N���#�ׅ������F�C���_��,_��2zi�#�Sh�?)����a�&b���Z��sU�ێ�a�d6G��0�|��J8	hG��Pu.<Џ~Q���"�u��TpW�L�x��Ȃ
�i�`�-8/�}s>_�^��U�i	��6*uNYi�-����\����w+�Yw PT\�������|���]��l�߅�hi�&�Ŧ;�ݟ3�\\�3�{W��C���m�ѩ�wD���"_P�)l��T?/uT	�"Bvj��"V��pv���ts�vk�#��C�����b��ܹ��z�����܄m��яg1�?#Lrd����Q>�Ypw�r6'�5D��w��Җ����
�,�;i���O�3qԤZ�ᓦZ#�C�q������:����/�n������Ғ-��7"��� ��t�D�q3�o���	���[uoP�]��E~�����z5ռ٭g嶓(��k�^&%��VG;i��p�8�ؿ�k#M���N%���㦲�'� J2�Xa��Hn��[V���J��搣*�����!�\��`\���:Y����5�
�����t#�%��J@e��r��d��}���]7���YiU�	d+��0i1V���\����s*��5�O�?��p�B�\۴q�jWV�����j��3���?�սC�o�_����'�[��؉$�ܖb!#�����顰^�<-L�s�Nʎm��m��ݵ�T��ǲ�''�;g�4x�ۡ�L�l�"�:@�J����6�N��@��P�������<O�Bk��gm�tm�a�Kn�f�m���r���>}GVC�}�JD�f�d�P��$g��\����+o#��<x\?0���|6�vј���ުަmb�$�)Γ���Z�vJ����]�Y� ^v�,�2R����q�"k�E���I��P���>����0����9[�lH|z-�
̬��@^�	��r=���K�Ŝ%3��\���*����@���+6=br�3�W�k��%�������L��`ak2ׄ��!�	�-���lHQ<?�Ɋ�o6��� p@Gu���_��B������#�W�U�:�YG�خ}���|2km6u~ۛ��ܟrR6�N6��SL�!�r��t�8�AN�����=�g�8��h� �ɾc����9
)�C��§��l���'��ە����PÃqV�o�E����ݧ}	$�&�>���o�<��]�dP�V�!Q�!`���*�Y�l�uɀ�I�uq�nn����5���w�K��I˨C�]?��`�%�G�6����!D�E��t^�z_�=Vɘ�m�3��g&�3�f���������������C��Sg���t���0��1}QG��0c��XX���d��� ��Ѣm_��ˑ����'�u�i���&`~��=D�?���涋�� y��ohgQ,ԡ��g��������}
m<~��.R�n�Ԓܒ�n�2�6�_��6�m�����h��X���QG��}&v{�^7���浓�T�L��K.�VL�ݹ����
E�!��k}�s��o�b�Xb��	~�ɨqk�b1ц��7�ɓ"^e��H��ƶ1�-�Ҥ�SE�a����< �%�LW�Qk1�D±XRP�{Y2�����~E����D(I`oi�����)]"���Z^c����_nF�����r������/������T��v�#�aʁ��ҷ��UwsG'��eT���<g�at�.��5���HxN���,L�d�
*�� �.v5�>����K֛I����m�R��
 �72��l�D��	6vSGe�f9����W�*S1�X��Z���q�oV.V˖�?�&�q��b��+:^��Q9�(D�[���Ϳ�r�;,e��%vh����RM�^�i����l�:��*�0"q�RX�	�zp�N?d0�e&mxG�a�۬��>�o�#�F��a�q�CZ6��t�h�m<�︋�d%_���&P���}���k�.�s�_A��?���ݱI�"N���'�?�	�tx1)+;)k33='�UG=�܆�c	����pnx !4�F���bg�Y�/�V�6�U��u�?7��lcG�*O(!k.5&�q�����9�\ZLI��N&�.�	�89�L6V>�˖���䨩(X�H�C���O���rɣkWd�X��i+M�K��N�f����ʩ�hw~Vo�kh<�(�����'s�GMea�nP�.^[[�$i�o�Ts�������.��m���_�Q�&��z|h@�%�c�v����0�5>��s=�!�⹡X*�$Ӡ���Q���e�v:������۱���BO��|>�~/���1�������(5{��g�l�_l���?�WB�n���9�5Pe�C�ǒ�}%���=��"C�(UzU[!�C��g\�t���f�d>oж+��Œ��&sl��:
{�]�,�W��f{�V=I`��3�` �l���-���j���h�2l�n76�ߧ��:p���d�υ�s6�q�Y��p��<�g䚕鵼7{|���MX@f��6��qr�����`�|?���>����Ә�?�O���)�E�"[��Dɧ�<�$�\��>� ��"�J9���.�o��)oZ���;PyЄ�F�7Zn~s���>��;��8Yf���;��uO��}o� 
&�q�ޑi�kO"�� |�SR�M��i;k/u9�.Z�
�+S���� ����r���~}��2Ci0���
����e��f��Nq$�pf�$�J�!ҳ\N�6���Ra�5���|S�U$�~�� 1�C)�����2|��]�%���R9SU���?ơ����lxr\�7�d��]/��_�����38�6*?6��P���8�xE�f�8w	��Rt_��\O�o�`H��x%D�b�p��7H�}V���R�p�C�r?-��[��.p�M?�)�Kr���d.[#5RnLԃ-v��8l��?\v�}Ab��B��k�כF����wG�"���4�TU(d�]&÷Q��WV> �,AT�;?{����\#3T������*nGa�4�L��UĚ8��E��bu��dՕ�4q}��*�W����[��
w�3$9I Pw*l3&$Db�д��YQ������PUM'M�	>�d�T��N������ڍ家�m�vZU|��h��k��������s6�@�0�v�k�(�� y�c����/X��mS�T`��O����~�כX�K��H<��H��i�*��i�(�i����M��'UnJv���#w e�{�Y�5�|j�����n�2��efL��ܟ_�]��o��N�q��H��u��IuH�_��|�݁�*�1n��iI��q!hu��ct��W�l[�s`��������[�гJ�=\�4�T�-AA�G�I`�[�����~�2`�"��N	�F5+b#`]>`�+��(^4;�Y�d���b��ee�v/'�3n�gms5���B����l����qN��lﯲ\��wUsu��@�K���	}9�Q���(�X���1�s�3�޾:����,㟿}Q�XE�w�^i�������6[���<�6�|sl��UCn�+t�����y�(w͙ctP����������?�F�Fw�"��Ϩ�?� %�
FWs���z��Y��[��:��/ʵf<8�ϱaկ!C�h>�4��T����*��N�1�U�J�c%�8T*w&b?~�����?�@݂O|�r�V��h�qNO�x���v�����朰}\�J)��Pܥ�e��Y�I��|�����B�i�x"d�z�w�gb�QN���q�5�4D����	�M�um>��~gTQ$ӆ�L�K }�,�=�5̏�UM�~�;�7ͳH�[2���U�S�3�}gݒre?�O+����aH2��-E���@¿y?_e!����~$,��5);�7w'�4X�\��:�t�S��(}���"e;I�,�t����咵�/��XzU.y�n:8�V�6�۳��V)0�6���K\�μ�H<��P��#A�PT��v�0�����s��c�^�@����_j��{��{��P��}�<���x�ap�>�ff�ӏA��4��Eë9=��;��Z�@��a�@���U����/xBy�T�f�������	? ���H.�_�u�[Z�ǜ�'\�V��:o)�WEW��uD�wi����΍&͂�v�ro�bP�G�)`�Ԯj|kc��svDu�u�<E��K5'lE�OՓ�T�����F�g��@�(�p��/�C����ԏ���]�Ӳ�	e����g�i�2p�|�"Vᓂ^��t���b�]��D�)1w�h�U?;�?�Y��VJ$`�v��}�U�����7WUe�dm�R�%�秂T��w�ԙ!�z�1or�����-��0�lC� 9�UW�|6��ǚ��@��DF��Y4��6���WQ����>0k^�5hK.J�>jw�]B�Nю�>�f?���z����<zG�5�F��M���4�߈}�_���ztz5~���+��CF��� e\z0�}�\�m\��e,��$9̏�s��_ۍ�h���=y-7�h߶��9w.��d�f��v,g�����;>����;��w~@�|���eo��+�sgq�9���*��&K${���e�4��C��������[�~�s�l�h�1����i6�#�o�:����.�{!�����`�[�!��xc�	�>��׳�	T+2}�1i<j>[z>�(I,������<
����Z�����79˟-��pw���/�p5_���ӆ�-���P�}�_k��Q��j5xЍ_"��T�1�T�b����*ϑhX�"����W-��{�ݿ�%Z� �41��;A�� �Pa[1Mw�DN��Ơ��i:�ru�%�}��<�a��<홇	���.̔���s%���������P� �My�����3�0�,��&s>��s�D�y�[��o V�����0���]����O��H��
��~gwf���4�dB�7�zq���@6�CY��]�#	{J���Yު��gO�k���;��O��{P�_	yj�E�ݩ8iT����{4���y����whg�XAR�s��s�@�˧�ssC��:���k��āF|�������
�(CT��HC_J����缇�^��k� ��;�7�o[,n�詘�ǈt?�aq�n"V�74C��*m`���a�������̰���0�m��9�q��?��;��r��'��y8j�X$^��@��b�9*��k.�f�3,��۵+>>SH���_l Rt�9w\�%rl�p�ju���Q�Y����g��j×�i����Y����p�ƴ[�Y1w����v1um.�pI���Eԫ�2�o��q�E3ī��D   5>���rl ��brY����Kt����ϥ���(U_R�rc��w�;<	e`�#�����3�E>����5�*�M6i�n���t�d����O�Nq�غ�@��3�&.��U�6��3�����x�.���� 9�E�^|Y�9^�>׺:�_�#��&b:˥����S�QByu�C�R�*B�����ziۄt.)� ���K���  ��t��tI# 
,JI)!�" ]"ݱ4�����y���qTv������ra
R���z}�/Tӑe��N�#�[o�ֿ||����١���?��z�zWd1b�Ջ�@�wK�t=�Ë���%ڃ�i�f	d����UN;���׼���.¬.V|>
v�;���~�>~�6-^��۪�0�,��޷���T��E4��}־<���6l�,��M�d�\�����W΂��29ml�[�g7fO�v��
*�N麭e2O}���_\��:��Ѻ�a��
=��7 ����`�|i�Q̶�+��`����ۻbf����{�~����"�{� ���K�$�.B����jXw4�:YY��)�tͲ��z3�Uj,��m��qz�%"�֗��x�V9&��"�To2� ;���d�YB"��PV���ɠU�h�=�F�lim���0])\�u�� �gZz�J�X����������n��^
���g�?kZץvͬ������
՛��<~F��^_�g�͟��[~�n��lQ�%u�������,��N��VE����w��˽������??�5�z�X�BK���w`�ef�g[���G���S�O�T��n]�F��h���ZMa����8���b�*=���r )��Qs��ec}ƾ�O�0���J�����2��)�`7�obg�W�Λܞ�~�I�O ����gn��r�x�ԡgg��CZ��*�o1˸|�+�V�XN8s�歘��7�S�E7H>Ov8Ϡ8�qHJ���5���Cv�8J=.��b˔1�fE�H��v�k/w��>,���Ŧ�8Q���0�F��Z�:��t=n�^7^��o.,F1�g ��y~�m���Bj.'g�|��>�+wR%8R��Ij0I�1�_np ��2��{4@����+
�	ؿ5�F�����[?�Ia�"��{TS4��fi���ٌ�ź@�j�ﲖ�݃󲻔t�U��NuIW�����C��$�/6F=c<��H0L��9+�1Ҫ�M��e�*��Z��.�d��O�RV�|�'|~�)�S����X�+���	�A�@�7t�h�g�G�團�����d� �t��^�nx3_�׽ay���е6����̴�����n�@���������,܅��,�r��%��� �a�6e7������s�#����Q�������=��7�hhU-�/z0���1����t*�y��7"�?rdU�
6%lʰ�I��㺎���]�e<p�¬T塾�����<ݮ
l�3?����yt��B���{�zoͮ�s��b�HDW�A�t��"�G˼���^^�hZR���5���/!����R���&��tF�v� ��d�%��?��u�T��R�s�g���WA#����~1P� K�h�����SB�xt���s)p#��"\���[�ܺ_u8F+ȁ����W���������vy����Xp4���lQR�����g�}/2�^9k�b�7�5���y� ��TR���~�oט���E�V��%���О���S߯�����o��o(.��P�:��L~�ӣ}���{Ճ`~v�_�S�O��\׮��Y�屼�qxa�q!���Q��ηッ�S�'�����ϐ7����{��)ݼ����)��*/��}A 5�###yi"���O�444�w�il10�K�J�G�G.�tl�I޿%$iH�A��$a�w�I�gB�M�e�9Z+T�X�ⅱ
Sf�x���~�=j��.s�U�����t�������㷪㈴��{�t�!��R�t�So/�O�Tp$w']N�|�G�1����W#���$C����ŀ����ME�WS����G�|�Y�[�<��}������FG�vww[��+���:G�z�A�°�T���=�����,��`�q)�u���U�t&����ۇ�(ޒ? ����&����4��#2*Wm��j
�WW�pt���)ьx�w^��W�&��o>��*��W��7�1�#�AlY��_0����&'��+J�[[O;:X�M���e�,֘[��n��se�Q	b(�
G����Ì�V��U��ߊk�g�A=�[Ε�1���ѺS4���p�0���K<N�������;��ۿ�ONm���\�jE���O�X2޸�B��@y�hz[|������f-G�^\\�����>���䖐��*Mnmi�655�'"�9��)����h��U���$$"�����{�X���M܄��N�J���l6�}	������y㱆�m��7^޵�M.z=W�^���^]�ϋ�[�%F�B��&��ţ���YG�2Ҋ�R>���;���J/��e�~\6���.�?'�-ύ��8��f��~b*��)vt��9�+Y��6�@��B�9��c���KH0455���I3G�LK�LJ�00�j��R���aT44�-�0M�����\�������Jh+*_��_�3V� ��e�S޺X{ځ��] �[#ܜ
��� ��q��*d!$(<��{v����G����v>4$&�㠎�݈�ř6b�K��y�R�e��Ku"G�'�4/[�m�e[���x7+�)���������?⇇݉5*RD"O��B
�	��d��o<��CYW�?�������F�Y�BfV�tth���g77�H�^�����o��E�B
;�m�����ĞO4�4�n�گ��nѧs���X��>VbR~Zy�'�w�A��%�46]1��W��JKgk��i�XX����|��qyz�:��Bj;���{��b��&��R�#-�aq���w}�=K۫?�W���-��q�C�-C8cdFG���(�^��������Y����*VNN���öJ������Ӏ����tq{�fw�;a\b�`���1#Af��8K�����ȯwX�[���8I��c*XM���R�g�1��ѝ�P�c��
fI#Vm����Y��-�F>B�k/E��ju`�c2�7���7�Kte������Ӈ��6�8�ﱮ3I5��H=�&���@tgq�3J	�������F}V��h|^�")ɨk���z���g�acoo�g�ںI���g�d�$Ȩ��Y��VV�)��k�C�&�AR�6�������:Z�->��SG/&�dD'�
�������X}�`e$A5"�oh�y�~�|�Bi��e�K��9+��uLp�e^��ܗ�/�H&�xܵy1��MS�Kn5������/Ok:Q�2�Cvv~�]
*��|(t�����H�_�k̎e����C."m�0Jw�33@M"v'��X�s�#�nh׾�#+\X���l�l��}��r�3}�N�:���sN����܍/���sh�fvUE�k@{(�
�y{e#q��9(Y�7~`��e�ⓐȃ>���1royt|��KGDD�&'��a��w�?�1��u��vT@CC��3x^J�G�(�єOC�_O�M�����^O�9��P�"��(Φ,��7�>m1�&�T�2�H�-1���R�K����D�z��z�;�����ֿ�^��#q3�S�,nC��(:���Ë�`��B.���F�o���Q*y+�0���~%U��)))HX'��1�2Vlc�j�}X ������x%{��ܢttg��ӄ�W�]�.a:
�C�<.)���ǳ9���o��}�~\�;���{���U�)�or�O±��z'���Z-A�Ji֛ݨ�-)`V_>�L�qy�ĥB11��$�����E�q�`��a��QE�	������xx�u|����꺀9�����}��o�V$��a���u5����e=O`���	�^�oa�V��+�HY��,��p��%=�p��O2^�ޠԂ`Fs�ʸ �|d��2�bϟ�H��-q��e��*�?[u��ݡ��KSR1��"��� �?w�8Q��`q
N��0�d��9j���C�{��DFFF`��T����]w�u��n��rYI����wж�� �&��f
9���~-U�������Mj����D����̙MF��}2F��1���z)��ܻ'3Kn�t`<'����f�]�@�Ysu�DH�}3�b2����O��/_�̸��{^ߐ�0��:�Dx;	��ݕtOI]}�����Ų���/�{C�V����m
����}���i�-b�q�^5~ZnS��Û0�:���ӝZY�&K VԒ�����@��b�w��S.�6�~��ш>UW��x� }�@X.�H����u���t�S�H��b��z�7��ha41";:�����"	k��<:� h	�oj4��"&F���`��0}ą,9n>MZ�/�=�ߺ%���,�	� ڣ��V���O���&�1�(~s����)��m?���R���X߸{�g?���������ނv�H\�>� }A�D���iP��6�Yמ�uX"��[muz�pE86�F����
(?���`b�BLxq~�28��o���:ܼ.�)$���۰���n�ET|O��mŻ.jh��y3,�[o�V��N�J��x.��X��a�x$���y����a��ک��F8�,3 8��zkvnQ���SjbJm!�+=CB	����|�ԇ����@qc�t�+Q3hf���V��Xؓ�����!ܴ%��y��r�������Ջ��sݶ ��&U_��"����������t��q��%�k��d'N㞱7e)�Y&���_t����t���X�7�LN*>����� u� �U�~��$K(<S�c��[�@ x� (�nU��&4�&L��4q��5{[g�����G�SI�1<�Jʸ��T8<<<W;=7W9�~Ǵ=����ݿ��N�06Q�E>���&��ѝ�`�=� _p4j�I�7���瘘��Ƒ�q�M��B�&��¶ߏ�V��;h�~K9�W�,�Ķ��N��BhȿdL�tk��$�X�%������P.[���B�>u?�o{�/*u�0��R�+���+~�jOA,��	�5�0������򚱩�Q��
������0%m�߷�V��)u(7E�S�W� 	��$�rq#�f6�cꋯ-R��mG?�Wz� >9O[���6q�A�s;R_q��CѠU��2��Kė-�-�G�m���R����6�,��0m���z���*�j>��nl �,�@�:�����D���deeĆHqR�2�Eީ�gbbHcgYXBfv���\{�~��3��1�ʧ$V��H���9j���!�+|������v��G'������bᐄ��|U��u��Qc|ͅ��>�(M��=<?�C�tG��!���_QۛI��ԏ�L�k����Z7����Rl��*XAz�r*))�.�|���2�3��.ls
s�N4������6g�f�c}�P\��F���G�1�o�����/��<�|!)���3��� r����佤�G�8|�!9��'��$&j��qdqN��rX8<V+�Bʀ��q�#	���v!���H��&���϶��LO�C�U�Ԙ�4�wu7�����Y��	��S����]�/l��ߖ%�$���-�.�Z���ub�W6��9�; ����d���p��uG4�z�Y��T�8�]���hۘ�����I���xxnx�_�Z�5.�o̎��5��J?�(4b�Y�4�Og�����=�"��_�g�G��}k�bYNNNץ�E��_����r��f���±uR%J4�h�<L3*
j(
E���M<�k3�����>�{�	-Y!؝wz���f�M�����j�%^�<��j���I�oe���o�K�vxԶ��(�,K@C�ihhڳ[��n�e	��'��#��m��qP��/�@?�JA��u^P�(����<_�KWRSKP;.�!�#�潎%Nod�;J���a�%s[Cπ����Ų��<���l��P��A�oA�hR1>.��>�{a���9�Ϙ�7Ȥ�OE�0�2��蠩�#HyZ�).Ge�f���W���<Ze���c�L�~9��x����nj߰�G J���TY�?��ͷ�?�EX��c��0�q��*-���"����kC����/�:��D�B�7Q�u� �"L��ʦ�R�<����:�k��躒ٙ�'Km���?����g͇q�a-�F���?}^C����9K����ab�'o���Ĺ1 �k84�̩MnW�Y�-d����f��֔ɨ޻�����f����+}�-�d�?~D�4kV�}W�7�,��9��j���S�0N7X�t�+��;9�5L�<8���$A���u�����ҙ�SF�t�A�x�����:u%��-��&wȡE�$T3�H���-T��6�as&�=��� �[�[�>n��,ȣ'�nm���X�p}�k���Z�b���ТSv�bK� �5��S{�|`�P�e<�^d����w�0A�/
$�m`г�����#Ҹ��4ג��`"&H�|���g&��YZ����JTn�g̫�i��X��2i���(졜ު	�i�ml/A� N<b�x�p�I+c�bB6F�UB�,9`������E��M�m||�VXؘAscCc� �]`���9� #��ѧ�����6+uڊ'��|���W^������%g�]41�q�q䡲�}$�H��:i�9�yG}`��2T�=z�So��?�}��qJ�6�L	�*kJ�p�[y�&Z�q
�d�UZ��r�J��(	���hR����$�ޞG7!'葏T�W4�Lm����E�U�g&�pX�V\��X��� ��Zi��3H*bQ������8b�v��0^��;�je0Pj�Eo{�kc�N�q�4>�I�K�y�>?y𦝰��笿�V��N2����<gc3������]Bs]Y2�(�MD�~DƧg�+#E�Hx�A�;�g��uXn7�st���.�� wqJ��]����R�1Ӳ1ǌ/:p��߶Q��n����v��B�"��y�j��x<�ʥ<�{�t|*	�5�g-֡T��{�g7����yF��C������_N��ҐZ���7r��&�Q��Z�t����z���	�d>|X��5I(V��bI�$q��~B��y��\^���Bb��z�n(��)̇ZF����}�I���>	�'��hC~�lA�i���Dw�1���WUŖ:����Z�4���h�M)�w�J93�2�!O\�'u�]Ƶ�{5z;�#��2=� �w���8SipS�]$��p8���ӧ����0"[�Z��s@�X�Qܩ��gv�~t�Q����1%����a]:��V�hZ���H�W��gv,�*�"&�F(tH&�)��ҼܝH�6k�$H���1��%ht���^b'�ثX �6#���=���ܷZɺ�2U�����z�pe&i1��S�Ŭ��"Urb�v�ٙi
�Ew��9�A� .�ؤ�P��܋��1r��Dh�N$�|�H��:
���=������� �j�/��Ic{00l'<��0���D�8�q��ﮬ�v�:��I�I�ɻZ�Ab\Lˊi���i�G�p���<)�oę?�Ԛ-�Lt��J����AM,D��}�j�"84����~k,���p�|3,�Ml�"|@����}"2��� /��IH����je�=�;�' X�l�V��3�Sr��H^���=H4�m����S�8�,mx�~ t
.b��g^��	Z��s�hth�¬�p�c��B��������4�v�ʮ��<��gl8�?�a��}O�|��j��K�MAx-���@�Ϟeְ6
�E}���6�\���]Dһ��N��|�#K��u�?�H3��?��G�<B��e���R����*N�B�b)�E���I9�x[jH�,������'E9�Gl��1|"�q�zI��o���F�&�ȟ<͏�ؿ���۫�� >4f}�� ����ײA�M��/f��~�Ԣ+)��?z(��K��ZZsb��C�C��諓��]M����|.^���.�e�s�x�~�/��� I����F�"��?�*%ǉf �Qi�+s�`EΜ�w2ӂ{>���9�Ւ�&��C
��-�Q9��*_����]`_�{!s�5����ك�0|4U���T���N�5�Z��ftaf���V�K�p �@�ĉ�U#�)�ںM�`���r�{2#�Աhnf�=�K$70�������A�ժiu�Z>G��W��'�������F�%+���������J�eJ��{�0��yH��(7^ML�W�ePh�'7H�q63��pM*l\b�/����V����/f������*�� ��t�u�����Me����8�ړ�\v]�^�-�zc�͇A9�,�D�����9y<'@��V��7ExPO �}�~���4���Z����	p��Eq'������7����S�[KAg�,5���^3�gn+��_<X�Y��#z�0$a�p�a�����e^XX���@ �^��i�T�g>�"i_mA�����ģ�~fc���/���JZp�j`�������Ц��=R�.g��ۻ�!�ܸ���-��,32����E���� �=2�<D�!T(&CI��4�[�1	fsC��yv���û���[~�f	�5i��DQ�ښ�;a=|7o^;?=\&y��̻�Ăd<uGGi�l+%�ĳ IXFi�4B���x�RW
�u7�����}fD�7�Y�F������	�棔R�W��׭4���e�)>&�<���aG9G y�`Q�ƖQ�H;���B�"��ZQۓç�,OR�־�SB.Hy�8Y��t�U�#�[��a���NO�|��}�/WW�����o�������'2uFdAM�3��S{�/i��&&'q.��Tlmo�����n\M��J�Zu��;�B6�u�^��;H
Du��s�S⑽�$@MU5�ZrF�(	���l�<��� ����}e�/��T���m�F�x��e���3�h��칬��xhFT�e`u�Q�Rx������3�m4==j���7[�	l�G� ò5��8oϔJ+[��|�����<�2> �]]���D)�!ss�SE�2�E߾�;���V8:9i��%����><T41a!ƽ��/4�������sR;���Nm�N���߁�a�;����$�c�����Z���~��=0܄ǡ���rN*����U1}Ђ�� ��Bj�i:<��HR�O�M#��ъ9F�ddF��`3���V����{59ƧD��=�����7uw���#�b������53|�T�ם~]y�/�6�K�2.u���=�E�����9���|�Eޤ��B �zd�G���4}d��x����]��#'**�O��G�T��� ����yO�X�5ɯ_��K��u��`�J�OD`��iFF΀A��.��6�o:,]ԝ�F�ZT_qCV_��:�U=f�ɞo=�;̈́zf�)T���k�+��Q��4�Խ����&���w���I��}y83�_)G0/��Me��q��8��uͭ��`����Z�*�������X�7i�鮿~#3=�j��J���8�F�<�yڪ�LG����%��<3_��H;5���F��h
����h6g�:&�����`�ZZA�^&��$)8�Q���'�k2d���}Efn.~��F���Ν���Pf��7�����c�q�Yɻ��]���O��A9�0V���+~"m�=��JeS�2䃔���ʵ��7�4�	T��F�)9P�����`! %CN�`����8$�����9��u?A�������5����1�tD:��8.���k����Ɨ��۾�����y=�)�f��:TЈ]��}��
�`�,�N��~���N��cL�y��|[ɫ]�4I�ݥ���'��dc�/�g����k8ҹ�s?�yؼ�0��d,�XG���c��3�M��o��[�{DU��Ə�Y���/�]�h6�8rD=k��#%l�7x�D�}��Hm�gӸh��KUrR��eԡ��v��'�p���'1k[I��b�ج���:�20tI���ol͈"ox6\]B�0H+)5ŕ���
D����bXSn�{~�3_<>�j�ɡ��\U�,D$}q�������1CGǻ����u��] X1N�-+h>@�c�
�j�����Ī�St�l&?~:�z�=c⚌Å�m����y��Y%Ay�+_&��6~-c�b�����ϣ�����WX\���u�t�b�����pٟPy�.`	
����m���+{����s�`k(~Lh��Y&I�fJ��x (G�1�"�=���ذ�am�����c��S@�u�ٚ*�r���{}�Fw?e��/���?%fz%�q�{RÍ}�q\]]�n���ѕ�@��>KQ�yɉrJ��������yW9[+��ë�i�4zfp˭�����Y`�e�2��3��`��y�p�Hd@�AG�N���*�p¨!	~��.�J�wee�0��}ʗ�e��pzG���S(�bb`��@Ӗ�A)�76\�2VN����������y�z���Б8����ŕ���&C�L�t�-����\]����0�j+��4�}莵�u��N��T1ʵ�"�'O�#נ�+�kkk�	�-׻^��e��Q�8�?��U�j��:4��<Cy�lI?�ƻ��ƛa*A,"�-1ǚ$k~��~d߯FZ%Nu������K\�]��ԟ"��oq�o�!#���f����NK�E�3]��~"�E����b^:_��#F�z#.����y�~��wa����[a��U!!��J�K-zl���oݠ�/�:����f�P^U5�8����t�&��[�_�#��`��"Eĺj'd1n�d!C�̶|��c����3�Vx_��m�����"�M�PJ���k�y�*��!�;���`#�?�c	��O��~���ǀ�*�,-�̥s6g;x��ރ�����h�wa�g�Dx�����2��ҙ� �ŋ�$�1����Q ���R�U���++H������U�����K�)�����,B��s�+K�M"�H�j$4Is��j"�lk�)�@�dh�iz�w�2����I�|�ꥤ�ڗ:ҝ�����c��c`����(E	h�<��~�g�r>@g��rT�A5�'�y��^���~�L�I����<�%�\�ϗ0���R�57���
�`;ZP����c�1%�O*1�/Fy��A�@
ZpLKK[̉A*����zP���"��?vK�����[����G�h�;��H��+�-�����$o�8�����*$K�5�DC'Pa1�Ç�7P��%�	_{��&�r�g�ܷ0��/HV��!��:�~I�������r�������g�~��!a����5?����.�q�2ջ>�¨�V��D�����m�~����y�:�T�n�ޓ�U�Pנ	���G)��5S?g~AA����[O�][\\K� ���@Ǵ?C���/�Ǌ2"�q�oߚX�"����^��d>Jta�;�/#m�(�K��i� �Sw"������"`�O�����嚹�4��Z�_z#5���T�ZA��FW�l��U��������Ar�|�8���ct��~��e��gk�)��:�n���dA9� ��
?W�GG�sO�ٜs++E

�����mMAx;��ӳ۳-�Hm���S�����z��ŵ��;��W3:����9@��c����xk��r��������Ѹv�žZ�N�8Imsh�w��V�槃!��Χ�Ls{�(( ��7J�_m~t�������w:(��� �#7u%񀢢�
��V�=��S�g�'u�����8���r'���˨��-���]�Ȩ.K����g\��;����A�Q�V�;���ώw��~�B��������VQȤ�)��;b������.Y��㧇� �O_2�ޏ��ZlfHV.J�OŒ���~3��ƚ,�$���Q�#JXo���
��۴���/9���4i�,�Lf@���b닔���	��l�6��l�|�4E�k�EFF>4���.��o�ݼ,P����AZ@"u�r�7��VR=�ӀN��c31�쳮���%���y� Ɔ��VVQ)1i�Z���w�1���R��N���s�� zZf���x뫾��+L�K���\��c^�7�&��aL�4
�$ο,W��]m���x�Xx��-�B��x�@�uǯ���7��]����_{d��Ccy�W�U>�:��72�ԯ�B��!^�TO���j���9��8��@gd=&!�y���t!p��~W���q�З.�"j���W8���+}��S[a��_��.v&��x�^�k��=As	

*-�>I�_c�5>�9Y�P&����{������4,4U5���)6&��A6>Z�$�|��X��e$R�u$�;�m*�2��	ȟO����o��3M)����v���2�y��.��0<��K��L R8[7�s�w=�P�ZZB�&�� x��Z�ȺZ�Z���zx^��>�zw�ek��q��+�䘔�|��w|���85'�PR���W��������5�?X%ٜ���y�����*��>�"��٫���XuY��Ae�"*fd��6��\k9O6b�?m���!rW��#Ğŕ��o��_�R��ն�UR4j�g��{(�����88��b����>S��9��G��׽�Fڻ��|���߶�e����� �2U�ϵ9��[W	a��JD	������h�Pn^ޫ����Qs�yyy����!��!5���H-T��폽*���_|��������MWW1���!
��<�ƣq�Ν�g�`�Z��1M%�Ji�${���T|r��j��9��Id�땃�C�&�a��Tk�􁴴�2 �}�.�it�n~�����J�C�@��	T�����8h�l��I[֩�ڧ &	E�7�����	� �NGۦЁ
	�߁�rg"��dM�C�Y�|bb	ΕC��Ɓ��:�z3���L~w2�࢞���GЅ<�00ں�ad�-xު����z�B����<�]3
����=nh{����w�5��������$~�4�����[k�#"���M�Dt�ӡ"� ���Z��*m��_C��8����-���+�g��+4��1i��rt��K7�q3=��X����m_av~����{ݭك�I�S���8��;���Mk��f���m��by��^�������~����Q�'��i�4���h3T�Ԕ+�[\U�gY�7=�M�lo��������4i[ND���`��z�Ff:�:����K��8�3I5�W�}�Kt��~�^�{�OZ�
s5ş���U�$Q|�`��(�~�ao����n������4r��&|>�n���7�QhXS�o�}�!88��N7(�}V�^Ó���|��
lh��.!A�= 6�迗���]�{��Z�)sL7�$��\�62������������Y�U�S����Y��+-S֩	�i����A�g|S�/�z��ê�\��w#��1���m�H�u$&:���E&��S��뿄��Ctq�-�ۄqW�Κʴ�[S��)_��'#@�-��Dy�W�[	`�<��Y���:j��������?��(�DXu4t>M�ʿz�:Q5�����Y>��� `��0Z�����0�Q� ��(�����-0�	�X(G��H̪�Q^iGL$$���Pk��B^��:؎�Pc�y|XY�$i�~?|��}��K&��ۢ�v����=������hk�C���tb/wX��v��E�K8E�=|vvFNْ3Bd8�\�
<�(0l'ܨ�}����`H�]�;KʧN1�&��.
!��<T�y�{��P� �h��|?4�j�����h����#�U�l'�ǉ��$v�f><1����P��.,X_�Z�����"�]��jq��/�:�0|)/�i1}���6��'�c�M�@	3$W#%�,�[�|�WN%�M[���K_�	��W>v�ѿ�ee�'�da*՝i��v�gD0�����*9}b�����K͒	��nsh��lG�:wux4@/�;_#A��B�V/\�]�h�~�{��v��t�u�|�5GK��/��g#bG�������Oi��XP�D��}���lh*6��y��׽:G�J+�ʥ����P�|X�~�9�X�����fm���#I_��*��m���999A����s��R��P/��+�.eTN�W�+ڧ�;�ƺo�L�#E.�t��{AR�,�þ蟄.ܵۺ;��"�D����Z���V���JK�J�a����`���C��β#���a�.�;5��&���{����@�Q��s�ďꌽ#V dpo���ԩ ���x��Wc��"h���}�I�|��������n�3������A�����Uϟ���<�ĜB�������_��Ӽ�,&v�%�UZ���)��*so>3�$���U�eP�`�`o���9E`������F�ۖ������G`����p��" ��|�~=��_��
�DBo�PY"�,f��0�N��tCq޴�$�e�gD-�����?����q��J����?dV#�X�9��ߠ{�(�����ⓑ%�X��Ru��I4�m�8_e~���Xp�Ǖ-�(�{��(�	�|�tg,(}�'�jH��p���z��O�S@���z|c���1KH�%ũ���aa�J�y�2���}�b�(�Sf��H��������� ��n��TˋM���W��Yc����|���ry��S��Q���_�@[�3�]�>�b͈_]��qT�
y�ܯ6�z�h.��V�.��=<R���U�B2��o߾��=DMM�W����S�$4Ĩ�|Sf32w�dǀyh�ó��G�LrΜ1X���2�Y��Y��~
��<@-��oZ �SqeuwCȰyߥA4��EfƷ��)-��7��IE�Dr����r��p�S;7�ӥޣ�=Օ~�k�u��������C��HO̭FJ�ۃ?�!#�q�<��0��v�	B��!F���Z,��.ǥ�F�q��XL[.�pjȽ��3��Wc��u��.���g�� ���hllm|{٩MQ����?o%�֭8gy�����-h�U�ͽr� ���c8pz�S�����KK˙ GkS��wj�h�-�1�笡Q�ѥ	�w��Z9�����!*H�L�_7l� �|Q����q��%���'WR�`�-����=ci�4j��V&&j��N�f�ȡ�V�*��Ӽ��y��4����m}k?�k����fH�
�r��͂#�7�kCy�H�F�������t2eeez��U�"s>V�"�����(�)*�@�Q���[F�i��fB��B��Ӻ�J\;W�eת���GV�j�>8m*��~#K�A���>C4��J��SA��]v��g�<&T`����@4�����H�x+J52�ii����o\	wh����N�κ�'�a�S\�R�uOu
Q[�E���U�U�:�n�a�2��|�8�:��?�t��D����Ƣ2����,*���Ɔ�Є�̘\�v��VX�H��d��m�`����^���e^z�Ե�p�j/H��ǪY�m`j{9���jYY��G�W"��޿���-Z��5f� �0��Td��; ��;�Ξv|��&I/��b���㣳�����T���Y��=�qߤ紁*	Jf	��8Τ��儘{ҷ`���l��>o(�o`do�>5��j�M�{��K<AH��������2�ӧ8�>�*hR]��a�������	��Z�������.113+����1�eI333�
�����C\��ݟ�	)((��1`��A���j����q���
�T�<��Pd�mߞ4�+�6�x���г�ӗ��7/N-��Ð��P9߯�f������5�㇞H��OP�����5�b�c<��]Jr0.=�E��mYt��,W����)+7^�� �#oz�@th�
A���Xo�(�2�N|�U�  ��$x�懡Эɰk]I�1Rנ�����(�d]_�����;�5X�14�[\� ��S@��pK�յ�����B�0I�U8���`�u����~{{�?#��yb���KШ����ݹ���*�����T��ڍ�e��)�N���hmm���Ȉ�!sۚ"����z�$t��2�}W_}�� =��_o�"V��ĺ�]X}��%kB�Eæi)x���f
Yq�H�g�h�ּw'�*�V:�����W|����߭��:���(�U�:c��ܴ�l%�@��O%�7�H��l�s�Tc�/��Yg��g�Z���炌L�] Ș(a�%8�4���<[�� �H����n/ǘ~9������������ܜ��X����ˇ-��7B�df�'r+����L2�e�����_Ŝ� �"!������~�@-��>�1���ɐ�����������uMgaiI��{r���5�w@�0�C��uS������?~<3?���3tk�0�����+Jʘ��R0������Xu�BO������TV�S��	�f��P����5}?�m
��QuUֶ�р		;�	�O�=��:�[D��+�탶��<���|�Ǵl���Ry =�C���^��3m�:G��$��@Y���Rk
�6&|Ym�4�j����P.#��i��jO�����K\$�N17z+��;)����T�ޅ��Z~�K���ᣔ:l##�=%�y���@N�Q��/��|O��y�6�(^�,n��APX߽{��ty�N�eY�s�ã���Ƥ{f��Ʉd1�C�F�`��1|��XO�>��ݵ,�!e��R�w����<pHOvO��l��]��[�@>$v���������-L�u��կ������f�M�/O�R��0� �T�@LD^vDS��K�a�m�od�F�t����4?Zz$�m�U�8�0����G�U�ׯjy�s�L�j1�k֍�o��G���q#4Oʖ'����G�E�=��p�2H���-?���Z�L�~�ז>���̳";(\��O���"��L�^hi��0�xˑ���
&�I�% ��*��T�/��Ķؤ$�ɨ�����iy���-��A���3���?~�7n� �>�1H�LH����K��_Dn���2��k��TpUTnе6��}�M6OS@SYsJ�_;��|�E�^{>���͆�����E*5N^�t �wwX��p�3hS�Q��9 �/��n?6�҅Ylv��N�5�G�uW>Ҋ���B+��[�����|�9I�);�r�-bq�5w�T���_{�Q�����;�&έU5�����x{@�f�Οvly�T��S��ĻE몕!�b�j#�D ��'f��TLL�����(��2Z�TQVT? Q�['�[�^_�	����s^P
~�:�����*����-@�,��:��I�RC��c�+��캶AJ�.	i�.鮡T@D�)Ii%�a��R��;���A���?7O|�����d-\é}���u�s�3D.)�t�ʷ����5;�(I���OF��z��%�������<��s��b�HƙR��W�o��1���9��'��8���P�F�&&���`7�M���h��Y��j��F����衖︍&�/���ǥ�����y�x�-g�Ҋ�ޓ�FF?������0~��0:���D'�]����@w�uLs�!��z4P�Z�tm����5ϧ@�����;C����?s���
�3[ZZ*�T�����=2ؖ��Ҋ@���*�-MT���ݣ�������-M���d�r�p��|�%>�^�u:]>�t�FKs�,zW���	7�h�l,B��;�8�9'���PC���1�3o�,C����󽎀fT�c�ЩO7��Չ�a�΂���i��!�|ɰSu����9��v�o��q9��U?�Ed�D����cX�ϳ��X��#���ȯ2|j�{�VI`���f�z���R�F��"<h�>���lEz�g��ذRRR�F$�wO�q?�l�~)-���Qu\�:��P��3^�����m�����4����ZO?@�݅o(%�Ջ3��\"h��H��~�괫p�����ZM�X}%��/��\x� &-w��S��){rM�W�1����������Z������sx^�D����u�v�?!�v�!�W����p �w4�cA���~���h9ٝ8��ԃ�����q�[�i*m�͆�����:�xӫ�7�u�����G}Q�{��c��O����Ĉ�Ӄ⃂���w��Ξ6p+��+m��՛B���O���z�J\�6M�G
4��X���kn���"S�&1�9H����?عI�ft�0���Ɔ#`5��dJ��r�����Z)	����3/���������44H�h߰j���Q�|�7޳�Ҽ.���k�n��������ۭm�3"��v���_�a�/r�ѷ����<b�H.h�N�2��DUͷ9�B����@87�I:a���d�b�>2�}:q8s�Ւg�_[���RI3{� �f�sI2OzĦϺ��	3[-qw6=I�T�`@@SU�#��NdoH���G��9�n���{̝�0Xc>9�T�4xcqpn��||�܆�zv����	=��[Њ,��;�� ..���
^��TQE�7((�J[q�?��!������o�IF����Q��mYߠ[�����'2�������OJMݵ��{��5m�{���|<i���t�9��_������i�H��$;{$9aюl%��v>����"��}�	O����f�g�߮q�X�k۶��ck�'O��w{$�2ǭ$��}[G����ڥin&���x\�~��I�t��9�`<��כ9����#Tt剴�l>�,j��9=����Iӯ���1��sf�M֫�4�6��{:�o�5���9·�rs�����o��zE��AA�(��]v��3/��sto}������x9֛�@8VN{�l�R���6}�3����a7Q�����WOܵ�ʺiT8��l�v���ʟ	��̓���8ը�Q�_��J"�INƕ��!.�G����]�+�y��o�}����b�(-g�������g#m?�dv��AfG�je�a��������c�Vt:��ʮ�CݘN1��5s�n}��2{�|���;�眮h����ͦ�� ,�Dߘ���ҍ��o�گ��dVX�ڛ�.�ѷ��d�@[����v�Z�nfaR������4�S�99evc�}��l��-��rrOܯ�ű��H�??jeeu�A'��4P0]�̕	�T5i�kWv���&��Yt�ft�0N���w|���&��
�P7��T���yO�u�F@<$���������4�K�C��6m t����)���{��'��ħ�qBc��빯��G���f�4&+�.JL�PZ�ܽw����=+���A�uoѮuӁ����i^nN�����B���0s�-�ev�(\��X���t􉾁l��T���9��a��7�]S��׷�2��FϽ�v�Z����\��C�B�	����uY��=��k��/�^��J�Q#ф��g�^�L�4��]0U�۱�Ap���)�]��*�����*O����n(k�:�E/G�K�1�v�ew�!�����u�-��˙��
�����8����dH�GW0���|F�χ�����QU���f�;e?�b�9����"��z89�^�kt���\�y'�Ī��aa��Z�pۨ���ZxD0���& M���?���8�Ag�;ts��rqc^�8}�v�����?3O3f�]~CM�IЄ̈��/�=�8��{l�!0Y��EJ�x��r��	=4�73=i��G����B��;��Ѵe����C�}<����޻��t?l��PSu"��n����V1$�S)k���=���G���{����hs�>�0�χ��2{�o��w2���6a�|5��Ľ�(��{�SqH��H� �%����U��~ɔg����:>9)��x�BRw7>���x��X�VʃxvL**����Qk+����`ʽݞ���~j�s<�Y��]\i��dOiA9��[�c�b��fsy��׭���fL�%�C�]mY�q�m��Q��k;�-(>�����ɈSɨ�5��n��(��ʶ,Z��ڽQ\���/�	[���߲pcj� �(�h�?B��)(�����20#41W�E�K���B��py,��6.���P�t�H�=v|�M�sM�P���T�D8c���1�7�Ǝ<�T�Rr��`�Y\�	$��q ��	���}�Ŕ���y��Sĉ�w�8=�%��[��gL{�o��'�����&��!����̇.|���8�c������H�����4�{�\]]��yQ��J�z����--O�?�5= :�sq;�^ҳ������?2]�Ԍ�C�UV�����J:u҃�ڦ}�6��� ��+W�U���m^���y.�=��=����H*��6p,R��Y �У��Iߴ\��Jj%���v��/П�&GZl�U _�|���S�c�C�ӕ����O7����q�tE�1��
*a�O��c��<؈X"�+ҳ*��J���I�ɴn���m���Ht����(��'�N��Y*�0�5������>�C���B8N�E���@�~[�§ ��RPP@��l����	bV�ٲ�9�=���"�1��^�L0��q
�F��^b��:�(j,&�ԛD���R�A��l9��퍤{�F������`yY/���Ni��(nMU�Y:��5L
���w8��(5_�j~w�q���h��p�6D�8�a+�&q;cH���)�3�� ���Ha+�����K��Ԏ�P4?Vг\	��Rw����%k=gs^Tkb��ϥ��^� x�Qf�Ǳ���FæWB�������q:��V��i0��qԬ�F��)(���\!0-"&����J�����:	�Xw���y���}�c%_�� ����M����)ǰ�eN9]׎L��+�V�~F�0��,���W��~G�|[��ɗ�r��G��1N07x'\r�:��1���-q�YCS ������.B�ӷS ��B�ÞEsݢݮ,UV[V$�L5���F­�(�5��R�.A_ `�9S�v9v�WZ��,*G�} �28�zh�L�����}7���4�x�c���5뼽��b���W(����
q@���� �(�T3ߺ8t�����O�doZ �C%���HA�#�B�vVx���ٍ�F�=��RI|F��wnJYM�<�.ծ�N 3�䓲0���miad�>��b^���^��g��<R�'�z�¡I�}!�'���B񎾿L���?��D�.Ui�yٖ���w�Q�|����aVZM�C�k��3����6?@`}�c�ӯ��4�3Jx�:�|����߭�%��j�K������lp��G��޳Ñ�ΰ��X:<��&"P�E��6�`�x��̚�֥ͪ��p�pޫ����;�sʟ?����E��nZ��&"9)���s�V:ך��gR�V� ����SD�u����2و�(3�IǳJ��u3+;�x�S��ϟ,���Kr@����z�_�Ƃ32A~FhѾ�qT��ф���w�Tю�������:N����"s����}�.#�.G�X�SI��hA�$�3���-� ԃ�k���r٠o��cA�-�9����tv�LY�,�Zv-�}��4to�b�ܐ�����Y+��e-߀A�̩D8�����O�ωOQ5Ǖe���%��!���U�E!w~�1 �u:0��%���`A�wO��Y>��u��O�OW>(�(K5�/�/z�N��!Be�|�t��h,���:3�}��f뇎�5�8^G
f{{6n��� �-,�b�� ���g����Z��/^��D� �K��Ug��T���j���CL�H��c��m�~��T��;�S�5M �x�K�E��[�3GWI�����3�oi�]k�����(��K�)��}�+�}Uo��ܽ)0IX�Ǡ�q|w&{/֋���G����c�ښ=��&V�0�)��m��0tά��ߣo�>�A$(A�T$
�Cы����x��M4������$���]�:^��̈́)=�*Bf���2�	���� hv�?�2X(����)�|��_Wz�=����cI	5R��
��0@�w���]a��<���=�<H�a��s��zo�۲м���+��NL? ���n^��]�	�Bk�� ��c�~���gG�H��F-K��p��Zم:����N<q�/@sNŜ,��Zf��z>���?��KY��ڷc�}�6=}�$�F&�d+��V1���,����U5a��I�����B�/5�0�*2��������uc�U�{�[e�^Ă�}5�e�|�L��FN_��2&XlF�t��u������>���*�}�'@�Gٲ	+�9Y�]%nȓ2(�>���؈|n��pp��Ѹٱy\�̌���x�D.
!l=��mk��]��Gj䢲���L�('/y�����y;��	Q\*6��M���t[ �O�t�z3$C��H�d�p���_!��ll�6��I1V-$"���s���0��e׋r���%��0�z�ذ�G��-x(@	�W�αJ^��O���n
lF��n`�<.�E $�^���-l�]���y6��[}d2ez�j2}�\�\�s�
Ec���;����W�4%��_����b��&���G?�k45'�j^��D�����g���V���R���ϗ!u��/���.a�,�WM8��.�	[�0	^��R�>je��z��T���I���bqq1���|����:)�%h�.����xz����ެ�P�:R#����]]��Xd8l����i[X��jZ����FRYl ����H���qh��s�4�ʡxb��xba���u�;J��Ⱦ�m��G�_!�"]qc�KN��E��{#1���#E�o(�.�n��3����yY����%�R�)"fV��۟S|��>��Қk�^<�R����υ܌\=��X�K���$��(���ˌ]�F���|j��Sb?��ݎ�أl=��Μ�o��5ۑ�fEJ�9������ܲ&��4 �� ��llHAȃ���Ζ7K|���nei	x�cKKv��%���8�{j�]���Ҍ`�i����I$�?��t1�V���>���T�6_��ݜ�����۳�k.��0� ��ƭ�	���Q�������|�z�[�cE.��Є}5U{��N���)�!�~}:�����nq\R]#�����e��S)������a����-1���p�y�
a�R�r���;,��|U3l r�9���*�O�Ý�~ݛnb�Iz���z���e/�sz��%�-���j6,�w�u���!ֆ��fE���"��A���`:����',��!�εX��*y���7}�<vE��S���8L@5�Ʃ�9�����%˞p�4�,;z�y�8�v��t��
�����H��֦����x"�Ŀ�Z��%/�����ss:��l�v��_ۚ��a��d�����e*DƸUJ�W7���.������[�����P���˫nپ����ܳZl I�~��-�ϲ���~�Y9��3Hs���	��'i�����;4�ӻ�2�ڄ<z��{bZTpii�u�&�b�\� ����kՀ2�S%�����E3��%�А �NAA���Mߊu�#���%w�0k@�>���p���Iq!f^į4�ù����]~�xu��ub�@|��k�E�W�hÿ�Fv�җ]8�uZ��?���4s(�.0�-X$��Vo�}�H�^Z-턘�����o�?e���;ψ�B�+2L%�6��{��|~�ӶMX ��S�6w��5I2+����L���5O��S�g���gt��9����>��r�Q���c�ҙz��?�X\���v/-N�Vʞ[K'q�,�R/|Q[}�[ɧ	UJ���Z~����66>���>�H����噰�A���u�����z*$u<g/�a����9U��ڶ�[��3��4�Kj��!�r$�e�� �de�I�3�~.�;ZCCVK��`ʖ`�4:`7��~^��Ҁ:�W��Խ����){�JR���S�������0�K�z�ėr
�+�p���Rp�8ѿ�ym���&���O�7�I��^�h�V�������&��}��?<��:<����8�Ժ=�����gwJ� ���[�^Vx�,�������?-	�,ŇZK���}�Qh:(Dc/���n��8"��5�;��5N0".�U�#?TWSyyy�l)BGu�A�S6���ԋj���-����/J>��W�PMP�w��4���
w����!�7!a��EL<;���]��O�G���M��D�-��dFOci�p#�7�t~'>-�3��iW����c�'��H�R���t���M�a��W┐�I� *���VU�q)l恚�V���/�:�N��y�S{R���}&��#90�E%����Ԉ_޵7e�.%&)ġ�R1����t\+�^&Y��Q����M����6�m��)e����CK�4�I:�~p5�Pt���w�æz��)���%����*�ҧ��d���1�k��u�c�{p�ڌ�H��&�׀�����*T��d�T��ƥRrI9)�а��S���a+'�P�C=��*�w���m��3��
ӡa~�.��}�H-H������������nSw��k��3,z�B�7��k�Vq��:�t�H4;m,��0���MJ����uy��O�q�H�����1kuX��x�70okt�,�ǧ���ʖ���ͥ<pVR?��~{��pw�(L����ăɲZ˝2޷��w'���T��9R�?*D-�ϰ��c����]"|g�A̭��I��Q�/�	d�A�:���ul.���\/�)y5v8;4�����_�\���;1d�C�m&�I٣��Q�F[�+����."�<����?�a�d�U���I塜ݱ�N�oR�s�O&]��%�E��j��k�(F3�M���mL?�O�^ܑm�u��:�b׌�}���k��R�%J <����KŴ5�,�Χ��HǞ���U�Ũk�򻛻��\����9پW`�E\�)�1�uNk-3~x���|�����	���0��}g`�-τfM�[��&�լ�F�-/���	���/��DE�o��WKlw�t����TU�E;>��a�NսC��Č����^a]�,�es[���:������5{�!۬�}��L4� �(���́��#;���ΌJ��'�B�ڭ��d�|�( >![�o���!��5M��ׅL�
3� P/z�bnA
$���I�p	wn	W��y��@9V�K�-�d��k�B'.55�QMkJ-ʙJ�L�uf�(�k5�A����)���ӭ�t���Ũ��h2d�'H���1�T
�^���)��3~(J@�22��`�h���������,��k��I6׽ﳙ;�%���z<�r��F��{r��P�#��7+m�>��$�|R6�܄D<k���bvO��e�Tt��2l{Ε_H����v?"�H������bg:ɣF����(wW<��]6����ZJ2^7�TzmZcbp���K�c^�y��1G�m�Wt�^�]�yߐx�J���/���h�����)��� �my�b���?c弡,i
.�@�����"�G�#I�e�:�y���A���r��!�����O�7$�#��H�L��������Ԑ�9���+�@TM�/��Ě
Gd��k�Vr,�w�%��V�Z���G�RH46kΖ�E>�=�V�i��+]���Ӂ�ܲp��_#_�M"$���*��T	+F,y��p�veoi��#BnY�h?.��!�K�g��i��QUs�SQs-�����l��T~�W�Q�|���u�,=���0}$A�m�52i{��5W�C3p2ᾢ{36_鏘����{~�L�;r#�DC�U+ӷS�K^ߐ��\��x2�����l}��+���G܇��"J��l�b��e�������<�|1��<�E��T�r�+/YM�Ƒ�
�kF�]��0@Μq�8u��K��Gܞs��E��S�	������5m��*ߓ z�����J~uv�7MD�7<�*�* �!RZh[�z}�$�}J{�N�G�����JĞ;ȏ�!��R�~� BQ�����=F���{D��]�:������L�i��鼛�Tq1[��#ED�L�;?{����^���v���<��onKS�FʥG̾UujO7z��Ҕ�l�v��x�'��=��io*:;�X�X ��w�%�)5_͗�������u�$\�-��[4�"�h�A�\8�r�����whep��ܷ@�T�������}1EM
�V;"�#_?)��K�������*�(��'D����r�#���u$�W�ݬ���xS{)����mv��w8L������H��cg�YGN���qG]g��	
H�uA���@>&$��N��
��uJ$e?c���p ȮO��+x�̈́ٸ���a�o�I��uӐQ<�j(���]����FGk��utJø߹I���J��!B��6���թq��(Uu?=>��y�Åm��)Q�jq�Io�ב���o'�#*r� ��3�W���qun���&�6�G�A"5�9?vҩ>�:��v�	Ju�yd2�����3h�юV�C9��t'��[��ʦ/������9MXˉ����=Bn��د�}�c��7hP(�e0`���#�� rs<�|@==:u~9��#[:$/u}�T���h��>)�H;���+&�Z�S5>\���u`��'�։������sxz<"z0�tJZ�fm7+���"��9,�̾��O���/�"�"� ��V���Yg����Y��]<-B	��I�w[m�����4�6eY�~����A�w���ԍۀ��=�v��p�����B�v���
��a�A�CE�P���V_9S��EB��E:�!�,���s�4�E�>] U��tD�2S`Aq�(@�W Ջ�P�|��%�|(�]�OW(_ݐ��+�z}����Ӻ	�8�v�����_���b�W�>���;F}����'I�:�?�VR~smO����>� 0���Ǔ�MI4�5��s�H�����q�0�]�J>+���~y�|��k��/���'Q�V|���R���߻���c�(#����A���j�ܐ`H�[�������鱌2�%Qΐ0v�|ޅ���	}�w�I:Dt̕�S�LǾw�%$
��E�e\g{@����ɦ�G�In�q3d�z�)�e�H��4���p�-֜�g�=�Ҍ��#,Ι}ݺԡp-��L	7"���ܱ�1��f�z��$�y�T���٥+�}O��aa��Ӆ��`H� �C�z<���ʅ�u���N�]�~WMf�l6�Y��[G��-�����Ƶ.�!��������di��^Ak�m��~�hf��:Yr6C������a�����_��c�a�@���C�B���2���F`_���{�~�4[�Lf:a0���Z(��d��fωMɸb�Y$A_9\Ti�4<��D7rN���MqIq9x6��z�9<��^�+�j>�:�R}H�^qb�(+�ݾ��O$����bO�s��^H ���tW�)�z���4�p� �?�:	����Bc�38?>^�Cpw+���j�þG�v��pH�qڨ�R��Q�3���n��8v�0���>�����_�ޅ��AVI�I�v3��W�:�A8��hWZ�z@�{�
̮��J�8��F�Z� 4��UywZ(b$�ާ��=�st�<��}m/\��o��xv�������>���#8�n�K�T�kY|tㇵ)�z�%-���;��W�畞�O~�#C�(o����Xl�Lc���;*@���_D�ʕ890���f%�� ��	��ٗ�ެW.Y�gƂ�������5�5ȯ�x�#����@���������y�׸8�A���6>y"�M���s�`j.��}U�<3db�0��T������$&y�/a����;y��E֓���r�K�Jf��aX���x���aJ��J1=���lc�l�Ӄ�s��+����άC��t�V�)��6��^������R�w�G�G5$��-��%�<{��L(ɚ:�1+٨��7Jn/�ۏ_�EO��Em�ʢ�6���>��9��(��pg���j~;���Q=�_|n���6�&�N��@P1�È���0v�lcT�Co zAL+GH��@{�X�B9�	�߾�vT�HV^��8�+y_	:T�e�b?����iP�Р\]LJ\�8���w��*E���w$ɗ2��&hMԔ�M����`���`Z	��j���տ%�.$Q�qW���̺��i���~�4ZˌK��m��W����B7�R��������<?<��X��֮Y,��z���DTl�2�|B�Q�h�P=�H�w|����7`� =�ܾ"HO���S���2|��~��ҷ�I�w@s��T�nNn��"����|wV'ȶxZPc�|����IpJ�B��0��~����Z����`׀h��7aJ�E���ޖ%�"_��!ucQ��d��L���pr��
`���Ԩ�0-.���%j-h��i��ʺ��k���WFo�L�LW5O�M҉m�/�3�T(��a�>��h�ف�Ehe��,a(0��z�携o�z��K���#�eP����o��S@PB�ʎ��)\%�>�		�(e��	�gKu�S�Tݧ��5x��(����7w�gYr�k7��`�$�-6��j4%7��M�ě��G�r�0���h�_�\��($$��*ʮ:��giǥP�L�S��=j����;ymk$�78�⟜�8	'���Et����<����zR���M�`�Ě��NŚ�D�z0��Q-�e���_#{���Ʋ����G޿�M Z�ޭ~ 5U��Xl$i�h��(v�ss)t�l4�N$����Ƀz�Y���3>��,j�n"�{��9ݝ'?�<PV�I�3��j5t�˔�����3��TLj3��;���T��b��������a4ߥ*�ޱW��fP�k��%��q�2x��?&%����
���u� t� k���\�Zx�iil�
rۈСh-@Y�>��B�O	����!A�����y�<$j�:���p��zV �}93��vH|�����$��_�t�[�� Uo��g�-O��T�ri {!���A^���9�D��C1�s�a�`'��*٠;�ldW��0M����,�}��Ǵ��+�p+y��O�,ioW�����fx@�I�}bt3���V����8l�W�eϠ�O��>n�Bt�@E�S?�fj��y�ة�+}Ι2��"�!4�囙��b�S���j�t�qj�y�I'QY�v�⮸�%S,��;P#X`���w|� F�tG��'��6w�륻�j�&R���ɚ Dp��
]�r�+Ԛ�p7;��̫�ꟕ�Dj�P���Ϧ��z|drd��A���=�O�p`���s��D}�^�=Qx<��A5_=R7t��qm|gI�s����d�$_S��B�S*%��B��>�k��g��~F�Հ�~&����`�H̋����v;�̴:��5��,"� @��pD�0� V��_X�#E��)8�h3�#�pW�P�2�X�^�p_ma���~b@�-�I��F�bA$���ֻ��/����7A?]ې��|���Qq@C��q��Z]������go�o�mV��䀹U+��9����q.��.$ CC&y����-pC�JU:��M�x��F��\��D �'+����!�s�K�6�l���l^n��2�<���^�_�I��d2D!�`��z{�&�z.ʊ������!��ˇ���]�c0�f3�s^*�N�B�qE����h�̊���	JǋtO����h��NeE�t��T������"IY��2�P"B�[�Ow��r�v��2�"�����??q���s?.1��M+yiڬ����uEz<Ж͐_�w\\ м�	622��ی�<��=~���hS�-&��V�H�T�ID|3�k���gO+^M�p�w� �tn2(M�7�H�c�9�A��1���Plb��b�q�!��w��j$�~o8~PXK1����C���my�`T�&Wြ�'kM2`h���Հ,��� ��\8�IT������X�z��u�H�[nK����I9�s����x�R�\��wX�㎱�]V̩�g�r�B�	����PK�#�^��YE+S�w)����JNtfTߨ0������i���a"zӆ~�9��QǝQ��� �7}��A��2%J(�c

b�N\�6��0@����6�����L�XlC�؁X�z)(*_:
Ln(u�v� y�.�r�l�I�
���_��� ��5�B�k�	������/��"IW��аTj8���B0u��&�Թ���^l����^v:��A��)�f�L:^���;�	�7�F,VO�x�*�u�ޕ/x?~���[��8���3tB)a�e:m>N��m,�$� ���&�q��U�� ��fv{�]2����lQ�KA�����^	�^��������F��<�G����\�z���WI��n�U+u:�ª,^:��ן�x�~�DI���� �3'�ȕbh����1��uV�ꫨ*2�.	X��K���tw��sZ
,
�X���W�y���H�Ǣ���&��"��n���x2�.�����M��a�����Ah��{Q&>�#���=a���q���Avᾄa��*����H��A�ֻ~�B���N1{.�	��"r�
D���vd4���N������v7���,��<�PmO\д.gI�]0�$c}C ����ɋy��yw)�H.nn�j�'��A���s.�tC�"]:k�r{���ӽ��F�	��֥���F+o�¬ÂE����9��� My���@Ǭ�3��\Yd/T���� �..#��u����}t��)&pP�x��[�[X	й���E�q�l@qaaK٩i�q)j�q�����irG1R��b}����Q�6R2)��+�
ʩ�/^�p��_����Ύ�����`�y9t�C��
Y�+@M�����v�J�vk2B� ��(K��/9�IX4�F��)��{�봈{�DH���P���8��)�}���"e�=������1�ӄ�"�/]����>d��{�E�{�-���!���7u��sm���c���]祐�Wq&pc"ҾD���Mͷ���UY�)E���0+�����p�&''g��a����GcC$e��%�x�����>c��Rc��@7<7��m�C����8)�E��R)F��^�M�i�֏(���4;M�U� s�%�8�`�;�F�D�a�ʵ�k�?�}�A���4��Z�p/B*��_D�J{��D��kӏ�䧛sm:+`p��1���e���
Ea=�4ȫo���V�W�Q� �2���ep����Lz�lt����P�U
�Cq���Jh�����ާS�m=������!�6j��Ar� �"3m�&��L�v�b.��Ez���Tu�:�����׹a�ʈ�:��(��I47��a�yi��ì��Q�Z|�G���Y
���kW�|�F�*�P�h�go{{��ox���i[�HD7n�W2��D)�b�
��rt� �G�M�Pa��[��wN�Bg�83����#WQ\����,�LM3є�����M��c�v�����|��6b �6�X�X[=�*g8z��Ά7����� �1���X""i[a�����4�J5��W�g����x@��+��f��aD:�}H��]={%j�J�$������;��2���ip��Hп�`M���}�x��Q��蟧��+͖�J�	��me@ ��:�.ht���	�9�	�.�.�Q��/�7�^uӚ�պ-�.����G�o�Z�Z���3&'i%�c�\��`J�&J�q�W6U��ɪ%����Թ���p���!m�� {��m�4&3��`:RQ�ǱV94l��m�r t�D�ldѸ�S��Su��i���?i�_�ZF[�׷�Ps3��}�
g&D�M��^��|z�f$���?QBW-��$y�~��%v_&���R÷*�`)[^!��{v��'�:!ۂ/0�0h�I��7'����M��ֲà8�������Z�xK�GvH��s�K\���.$g``P�ԤB
�$$P׍Zݽ{ȗ�1�NM�_��k�D��dv�x�����Fw���><T@r�w��
&P��霻CSR��d-��1��"yq���
D�kᎤ0~ݬ|%Lnh��7���dCk�3}�pj���z�����y��
)��8C�����&Į���E��~�yF��Õ`_������8ǫ���U������@��ih@�����;����}:.M�i}}=G���z>%:�q����ɱ������w��	{'���sg�9�=T���i=Q",H�Ю.����֖�piHa��!�����d�(-�+P�����I�xN�gW�F8/��X�zR��k�|Q##�+�A��"�J`#��_���#�׃D&�������[h<	�4˔7	>���������QB+;�v+.W2�F��Ϡ."""h���� �[.ήe�&%Q��<��PQ����w�.�]�}''��㿞h>7y�k4V����"��?����^)���G	-4Ao��䏲�^�WR�bna�b}E.����Q��R���~��)>)�Y>��c;� ���xw�#'".qy���y`Cؘlgo�:�����V4��A,��ob(�7#�À�\~���y�ɠ!Z|���)h[i=�����Y���W��?�|O���6�zc�p*��f��9���R�����o~�A�^����]�X\B�VRR�̰f�R�xH"�ul���S����V�y���M)�K���`��X�������H!��]��.��w�F���̀���޼�⎋OJA8=m:,&"t�&9쿟p�Hh�p��
��8���$0�h�5��#"X4��	�EEAC+�׿���'
�8S�%Z��8�`�Ä�����ݫБ��$Ѥ���˩������e�Z������~h�͗4qm�����3^�3{�V.���f��^��%�I��َ�t#>�Y|l��Ի�t���׭瓼�'��<K��L���Oњtx~덂��:!�/�������V^o�4K66c�d��~���-n�o����r�~�M'%%���߅�b��XF�1Ա��߅w�ͼ>Y��EWY߇QQQ�L�x�|�:n�����D[!����7�=��#B�`v]V���o��	T\׊k{�\�O�xpٚo����A�[���<8)�{�l�h�lG�w����P$��/c.���ZeM�mc�1��V|��ߒ�W<��d<���G3��F\��t��N6{lb�7��4����~��M>��LZ	�JO�_�-���^�͗��:>��k�0��If��%z8���I�?���@;�����4)�[TQq{�q��F���.MП?���_D2�J�s=��Ƥ�oa�{uXX#33'���G��TӪ�S��ϟ��\덧_�َ���7N\�Q322����Q�6���?�qC+�.��<[̀o��v��1��[���%ݞM�L��f�[#�����R���,r?�p|x��P�8�������n�	�7������K�����-�|E�=�up������6�6�|֍���M�s5EC�tG�>�LMa�Sp� X�pdl�����xO�z��'��˶���\��[|�x*�׹]���@���^��q�[9[Cc#�gNa��H�F��R�h\�H�l���դ.n������R{��]5ϧ��?�����4��@@Um��׸N4[<D�c��?��iV`��2Dz�4Sn�d�����~�0��ZȻ~�3�/)��=n�˶�'e!���9`;�ޕ,da�>Y-d�9�*?RLl�g����\�{w�|�
#��_ZЦ7�)&W-�,�������Ao�ͻ#�s@J���{���. ��UZk�����a�}���]�9��fg}��]a�o��9Q�� e?=^OO����@̣B=�L����v����2�)����%��+�q�Q��&\5��P&�|j����'[m.`�˾�M�f�'�֧j�2dR�	���$P����D[[P��7�ige0�U+	A��ׯ]�4=�3���lqi����������sv�嶶ʯs�q��D��}�c4�')Y����[HuCCC��,|q�)������릑��me7�����ǩK��ܙ�ii��=�)��s�� ����
�
K���@�WǻU+��@�A�|��>if�;N�<�����T~��^ȋ�y�I�Зe�W���⫝&�����Ew�Hƿ1�љA?�ߵ�s�y~�9�/�g�Ew8U������Vw&�n�v�l6����ߑr�$(}v����������[��n�x��� ���:U���nH���K���ե�y\��Sj-��l�t4�t��'��,����)��I�~/��������fY�M)���AFV�vz�=�&��N|G�`�o���=��l�>eȰz�����P�S3�3���s�O �T� Jɝ]M���&�X��X��<1���bO��_���z��M���c�+O���9�ק���T��ku�H�_i��\��bhh��qqn.[ƫ���M���c�v���|��j�'��F3�`�OMѯ�G�����W����V L[[{Rw>�� �s�~%��Zt��߿�?@<V�� ��E���;ou��w�nmBB�B��dm!e/���%ٳ���N��Qdٍe�2f��Ԍ}c���>S�u����9�9�y��9��\��z�_������md��h��:� �E��^ա����/.�!�!���3�A�ف8�p�:i����lomZ6ň�	X�������7-���)��$.�:v��9z���@���Md�|��dd2�趻AY$ '���#`Q�����H�HHL$Lg���(��7\���;UH@�_bs�) ��J�Y�o�~��D���K'e��9\����
�Z�������;�w-.�����/���^�k��u�Vb��C�%|���b���Ì�k�AN���JOp�l��t�Z y1�j6�
B5xR���a��F���&�-�NBB�A0%4<<�$S���"y������������Hf]U{{����J��׭{w9���R9�� ��!��5r�s�����)�q����\�
.�r())�V:uq1�Ʃz��+ܛ���i��'�՟���Bv��-�ZZ^���|v�]�����������?��Q�-�_� "����$��=`�IcQ���nH�ڞX�$O��`�Dr���@���+�Ỳ�mu�Z��� ݮ�i��AL�cQ���4�u��rJ��q�5(�߁9�
���xLmD�{uO�ٴ&�������o��Ehá9���eȌ�)m80$*i�ML&��(��;6��
���H/|ОZ?�j����$��!��<	(x�o4�{�'@�O=ĥ�V�{�p!��{����8�U�����J��e{��K�������@��K� ak�H�&j~/����o������n6�rO8U���J\�ʥ�H7K�* '����]	]XX�"ձZ��|]�[d�/_�<Uq��ѱ$�;;�?�MO0%���1,�HX@��+v���T�E� $����AX����NK�Z$+������C1���*$1GIZj?�`�-�7���IK��/_ު�r�JQV���w�[F��\�G�P�m����q���	��!���⎄�s������@�睙��&q4�����ÿ�{̨������ $f
}7׼j9F�@
�_�Mt��ý���'2��%���- �d��8ށ�Ds<3$smk�hjj�W��Vd^���J����Ar���,d )�6�D�,�^ɱx��� ���� 6���.P^,��������lI��lu������PB��~�H��k�pK?�W~G]kZa��xKH(̗�B�]�,��^@�7�~z�����ђ�Һ���u""�A���Z������7�^ѳ�2 ���Q$^�-��4^����柡�vn��K�}�	P�G�u���]����?�?Q��� �����?�i����=�:������Zɋ��T��M��}�}�ξ�u����+��8� Jκ���I�.�N���ځ����c�bΌu3�SJ�_���d!+a��������8��Ͱ��?6���'���mn^^X�m�ۿW��~�b"+��(��|�ĵ��z�۫r~T�?�"ۥݰ+ՠ�S��S��^	0�����X��xS'�"��r��߻��\H�Ǌv��w������7��5�>f�7�	�LX�OW���3���Ԝ/FWis}ȹ���B'{���<��ia�F���Aq.����s�Zp�v3v��d�p�^"����k�y�L�ut��I���V�(}�c?��IG�U�Km�;�ַ��_J�~� ��ȱG8�i�r]x43+�oS>++�G�7O�n�BD�]����#��M/Po��F]�<��`�P7i��!vk�1"+�޳q�dϫC<H،8f^ű��e�����M�Փ�z�,��4YX�U9'�]�6v8��Ү�r��ҜL�N�;�J;�_yyЭW+���%=����J8]�t�c^��x��>��_D�?ےrIǧV�3�r��@WS~M�&�D�V��F^��@���%o�G�f�p�(�6��o��>J��:�ٺ�mR��K���G�^���=:��#rS]u�B�fQW�O}l.�f6F�ȫ�*�{����]2��V�:W#s����9�H�.�1<IH�<����#����W����,V_��=2��[{�������nt��N���ȭ���t��C7r(Q� ]�Շ%&S"�h��K���2�%��P���M�	1Y���/��#l'bq#�<��eE&���c�V^no��*�190�aD�辰�o��	V�;�ؑ�)���!���|��1ޞ!9e�G��X�v�hIA�U�B�j�׃���]�q��Ѝ�8�2^���� Ka�ۡ�B��֑�ٙb����Ɓ��m��V��+�/P�f�,E�ڇS�){ߺ�%��#�g�t;A�0���~t&Qv#�\�2CQy+�6iv�����@{����|� �z���j��^{�3��88�)����a��iᤗ��*+�y���9ƶ��3Tu�Orw%��{��#��t�}�{�R%H�Nl�%\�Ԫɭ��Y�c���3rxY�X�ꊼ=
�G��$�����8a�HхK� c�;y#�11t�u�����#��pmS��D�{~^����G�m�������Ǆ0�!�Fn�d�-�m}|V�;��	�`~׽�#��{#Y�Դo�������>F��U���)���&񗌔KMw��f�����fFҝ:���C} �CyLS�6C+�&�.�Ӽ�).�1􆄵����KC�ڊ����n����]X�2 ;�K%V���8��U��O����T��`{��U�f~�V�zd�(|����s[n�A���RH��b�������o��Y��#�-�JA�"+�TVF����5vy�b�r�,F~��GW!W�J��cs8�bp�sM��7M��
&L���-�~ߴ����!-��ɢ|ٜ��'a|]l/��n^Ш��
>`�.g{x����
e0g�����LR��4�	^��&;��@Y'yw���������K�?�����!��]����t ��^��H�:hJ=���o����=v��7/��<���ЅF'c9?brqje��(��0s�ied�&6�{Oɍh�����HԾ��Z7i������9�,��OO��P�I\2��Q�m��B/7I�U��/�f���t�)n�P�'D2���ߖF>`жjY��Ab��!ޒ�hlҐ��wU�7r�����Ϭ萕�[��ަ�9"Q����I�7�Lc���������)��R�f��M����2Y+H��Ss,Q��,���
@��υVB���4s�<*-b�U�6��&�)�qlާ(힏!u٠s"�����vxh��Μ)kG7�1A�����T��,<��I��K��W?��a� �X���O�u�ǃ`=���^锔�p^E�둝i�δ��;�
.�q2�P ��=��7k�4���_���L��%%�婝O��W�\�i�|��U���hIY��<-���ڊ�����ɱ
ۅ)L���8F�'%h�����8[���\d�Cu�$l�
���/��0Y���i����D'(���?��ھye[���H��In�a.����$E���K��(Q�hk�4�5~,B��653b�^����XO�!frTVvDNp=@s��5��Mcg�+�������A.mP�N��s��Ϯ`��Л�|H$`����VS3E���ńJ���ۅ^N+�|�2�T��
Ё�!�}JJ��'w�6~�. vFxnp6AĲ����9KokV��q��T�S�c)޽(C��ut�+�tA��ܻv�P��ϱ�$0�2��xM���pz�VĨ����T)x!�X���,��; ���䢽}��#c󓼨��i
��0����D�%7�����,3�
��S%D�Oq~{v�.��.u�J��^{���R�ڹ�.������sAYHy�k�-:c"��}K��gU.�ɜ��p�0\��wmR�+�B��l���2�>�Z�.bP�}��9؆-L���T��qjn�J�]D^� ���%qfnlhHU�
� ;zI��`m�IW�qO����fk�.��J��r�τ�W9�YL�N 	��8�\���.7B��W��Fq�B�|5_W�^cr���q��ٱ�Y_�c�Y�:W�vt� �z'1N���ஃ6 ��m�(�!��(�\������+�k4Ϣ����5T+-��!�cTr�Ā
*Y,V7�A6�S,r��iJ�-S}C}+���
L;m;�GU��MVV�l�,m����%��&�I80j\�Y�Vx�(��G�@8#�_��">��d��Z]��v����Z>*#Y��Q7����%��$�e��/�'��{9�wj;Is�n�=�7�����U,�(���(~t�T�� $Q)�>Y<"�s��^$@���>lXN�Fe�iX�_��-&09������Ҵ�ŸCN/Ç>�5 >�� �V��zu�dS[Rxİ�h�+|R{m�x.H�d��B������<�=:*����ZkjY7xP�T`��Xl������c�Y�nV~q	C0���)��^��t��*%͒e1|<�T���an�}D���cB�� �mu�jb~C����xx��P�sp� ��G�����RW�[��{��ʄ�F	��X�vP�Fs�-��ѤT�|f����C��d7��U�V-�}��I��\!k�>��Q�0ny�.��O/��<5��抣�QE�ؼP��n�c�68��;�N�R�us�G���_�r��|{� p�Ip�a&tg�+�3��Y���a󾺯�s٪xU+��o����P$���u-� ��v�0bF�:g���s�[��PCFta�E~��1^�hA�1���ګ�qG��K<r�`*�g[��?�f7b)���r)��3yke<�M{Фf(`nmA.i�#w����Q�o��,�#(�hN]�\�2;� ;2�j*�U�aoXX�����D`�B9&�u�{��x���Ģ��>N�~^�xE�m/�k��g�4�'��v&�	��@�����~1��_�J�z��YbJ(���A#۔e\8Ne+�T�[l�\E�]���Pt�2�f+�_�Q�Y$�/10_��=хھU�b�|en��h��k�Ӗ1Uq3��W���k(���+���2zT�Z^����Q�i�6ꔯ~��wֳ]��A�4n��A]�������/��:���կ�@�^�~�)S�V�����L/���|���뇋���j0���|��_�:�(�@�_`{�3�I�y(+�k*�ZP�>�>X��<�b�'���|+l�nz�ƶ�q� ,UdC1������	ߜ�w66�\�x�/9!�Y�)�׍��̛*ᛄ��9�>��v��9 70��%��#����	xr,�YP䙔_��U� �k�d]RU,C�γ?�=��$�hK������?y&�L!K� \fcU���x}b�!R�m~f:B���F���z�o�_��G�%�F@��Td�C\�[$s�`���עy���6n1A�'���}���^�蹅��)��=�Y�C�f�����P�i1S�w���,�$�F���� ��L%�����
&G�3��=��N���D��.�S���O6OR�yx�x��󘸒��$w���9^ƿ�q<�&�i��KR��.n]��yq#�m�O=�����]}h0�veW,H<{��\C�sr����7�יV}��b��HYy9,�0)���,'ehG�X���Yh���520`!�9u�@���]98��-������O?�6
�(CL5����M�֋Pa��J��}'l�;DwY����yߟ}�zNډ����ɖ�׳�[گ�5z|�9y��/1t���딚� `�_+y��)2�om1�RF$}���U�9��#lw��Y�DIc,��>������Ѣ��6H�[2b{;E��H��nA�'�{F�)o_fį�q�������$�T��!F=��N����ff���ώ��Џ�by .�A.��I5�cƃF��t���CX��]�'/�}c"�"{B���}�	i�������ɚ��؄�MXX[�����LH#ksu�oL���P�8ÁߧO1�6Ap�M�\9OP7��ce���v�/��nn��]�lO�=l������Ht�Y�u��Ɵ�\�<hмͭ )H����3�L����@����V7�Я��I~�����P�2z���l�������$X[����g�B$�ǟ��ZS�؏���L�X�7�n�y̫2U�L�>��\W�:�fSI`6?�i#�r��Sh�3KI��mH���ͤź��诧�f4�w:��ف�r����m�0������P����q�(O����y#Ȼ����y����?��8��:2؃�Jy�=ol�EV3#�SNThgA/3��?[\���T�TLKAp�B~��)�`�NtEd���Yߔ>��!�"��fWn�(����.���Ȋ�ѺԹ��GG�d���r-��~��k�㝔�C��u;�%1��K1���x��V"��^����G�'�v�828����iD��IB\��M/���޵G�.�,"��tn�X7�.�x�b�P��I�Ŏ�ed~�D�Vg�j��J�G��,�)8���kʲV7��4���m�},6��1��0%>R�!�����eꂕ��Z��#5�K������Ԧ
��j�n��'3��":��	�9����L� sZ��x2�]a�׃e��R�w�����[�i��=Vv����o�"����1u����7�L��KŒ1}�]��eO7gZ7�����]�W>C����-Ӯӭ��ھچ>�/��ˉ�)�mR�HFF!�Vb�~ա����g�9r,/F&���s���ĉ�m�W�W�D�ȡ���
s�R|7���U�����ӋȟT����'Cf�4~eM��=�ƞ��?����u�R��1ۜ��6��Qg-�5шC�Q�C���a��5����gc[s�O��`�R��Ӯ]	3ӬC8I�ф�\B��9��q�+ʜ17G z���QE�2D���_]yM��T�JXA�!�geXw긚�Ewj%��|��6eI����������̧���o�� B���|i�y��v��w��XӼJu�8��i|��8�k�bc�>���WC�O�qR�'sTg��l�Hc�Ձ;��q�ۯ]7�a�}'���S<����5�M����}s0����Jz3r���ԗ�\7���N��� ����l�R4���gfԔu��Jg�����IA V|�	�[W�;�$qĚTK+��Q�/Dy���nBZ{�����w��Z+Ԇ�z��exS��m�J5,�{�zYB��5��1��eå��H����\F�K����a�K��O�ニL�<�O���{���ܼ�W>�3��E�_)��en���zW�GT�����t$=��>}*���6�S{Z+?Kp#�bw����xͷVL|�
jM�3T[�,�[%���|�k`��URjyF���ɫ��������n��@����P榺	�9VV�ܴ���c��xFB��+#�=4G^�\�~g�-�gv�A�����Q�&������WS&��'�-��'�l4=�AK���uok��ǫkc�ܚ3(]�zN)�u�����R>��}V����s�����&�0b_Io�����U�,28��J���[��1e����Ϫ��?�a�U�8��UEn@b�W��~c90�`$R��%�5��Ss�v�1�`���z������6��)j��6@���05:U��ij��Px/��{C"��ԛ@V�ƄJ�r�J�~��[)�jA'�k�b��Y���i����Ȼ�Қ�yZ>�܊L��٘�5��J�Y3�zi]J��!eED���M����
��k��X
W�6�
a+:f���߼d]J� l���؇��[�z��ՙ�5�?��3���?���[�^��l�m_"}�a�9Ⲍ�h3f��Z޵V��]���.@O_�����o��E��Ka������P��*���Z-�6��`ˬ���m!הI1-���,Z��-x9��n:���`S{��Wa���=�wz�o�w�Z�	�D\�&�	9�%jǓxg����c��O����&s��K��m�`�#I�,�/��=J�M���%�
�!��n�mu�:%z���E�{SJ��]�m<k$���Lz�����ٔ!��9��\r��.5��%��d�HBL��^�r׋��a���<5<�D��n�pv��������%p�$� �G��~.�N��~.�@e�g�8W��k��ɚ\t��?�)I���d���6��Z��]��4Abϯ����C_^�xw���+z��Hg0_=c�̇���u��SC ��z�P�06n�I��� �\��鿸�,��)ÊZ~=��RCR@����+5*�[_M�8����$E:{�A���P)�R`�{�+4�� Π����+V�X=-�o�<k;Ģ4�^��Z�L#�
��2���1W*v;������-^�Gf_ono������Z��.��^�4,T-��T'���!����SKoS�L]��뒛�.!��������wJ���)�zT��B����/��{F���w�Z��Z{�dW�ͺ}#�A��0&a����b�2�Ѓ�q�gJ����q�	('>#�YX����Kq�8�~������g����V4g�w�t��=�Ԝs��g婵K�wѠ6?���>3p%���NC��W�9���j��Rɇ=z�
o9��P~����A���/=��kP'(f������p4��Z+�fP�N-�L苼��峒�0�8=��H�����ȦSR�56���7�g�3�9x�X���48a��e��$�%�{o��j!���%�6�I�G��_5�~� "\:�O�i��*/�̗�v�w�~b���	�!�򦌀�f��a�$
-*�&N�85��&�i��]��k�R��;��_P��s�g��3Q�ꦾ���Z*Ka��S�Pcq�;��g��wecv���⚅ˍ^�׸�q��6_IL��b���e�ҡ�?ե�Ⱦ�׉�LHw�ٌ������_���Mv���߭�3��y�>Uf�|S��s��J��������4{h$�T�r�_��Z��{�Mv�h�a{�	�'5Kj�Բ�-�6	)�����ׂ��}�2��`Q����k��(���7�aF�k���2�o��z��7>���I� ��gm^$5%O�7d5ߞ���XpF{��Tx F]ߔ���2���wޝ���.A���ŏ������A�Z����}�Ҩ������I�G9پύ*X�'����=Eʍ�2*s(+�1�F꒙[��T��	J�EIZ�%ww�{�b9�s�P"mJ.n>ߕ0�M�A�rU�mO�(�����/����n/��5$�l?���8�q�������'������ ip;��_u��#��2��lGX&�a�ww�9�m$��~s�x�w�k ��ƒ4ʯ	AY�kBd���P"�pULz�|ؓ��į�������Đ6s��#-~e���Vs��eB�t^�U�?W&9����|�9�n�L������k"�=�~әZ�P1f*b��t|-��fX;%����i�J��{7���[.(����@��,W�4�kb%��t�0[�#�CM�����^ݑy�V}VljYGR7������ҫ\��2�$�z��gLԴ�'nH�V*
I�ʅ]��-�U�9i����ы:�2��r6g,��H*��e��"�dф QZ�����oJ�ۓ��z�B�"�#��ӷ2�ʰ�t{BgeWbWf.�x�«��ɑ�:k����l�^�R��M/ƃ�bJ��\F	)?��� ,�M��E|�*��/'�Ԉxnnv0�mpgOVļ絗��-�����^��R9����:�lQ໔�}�`��*q�w|�qG��sj��fblt5U�@��Y�߈�%u`�"��CÔh�_�% +��u�#�#_}���N��~U�
�`g9��X����Wt��2��p�0����v��G����ڧ�X{3�Q���FK��F6�bx`��⢖�8>>ْ�W��4L�\hs��a���c�tw�{u½���^�,�c�ƭ��#�a���#�!m�==>UT"��MB���Ms8'[�p����}	ótC嶧�=o�|�yMi��ߎa:��oU}8�#fO��VLac�GQ��lե���-_l���J�S�X-.�"�^�Z��������N�Ў�R�9�Y%�q��*���H�=q�A��A��9�n��z��m�-�ۉ��k��(S��у"WA)P����:�@��������_W�2p��;�le�+�����C�6uv�O*[	�و���,�w5x�o��}(FY-T��Q����-H����rV�L�$���.�[�k���N��C��Ȥ�l�m�>��ΡP��p��à,7P_����V���������q� 2L,�� ,|½��@����\���aΐ�$��AČ�8|[ڕ�$h�?6hޗ�^,˜�v徤�BmKn�!��|�Y�>)������:�X��nj֗�{;jZ�wE��U���|g��9���S�i�����t���e�1Ce���D�֊���z��I��v�D�ɛR��䫊E�r������
od��Hc]��I�$�O�^���Lx�{�ea���y��B��C�oӚ�9���=t�������#Fw��t�\tK��� ���Q������P�h:χ�,����P�;��R�ڑ4�ݩ����4�	o�A&��r����e��o����F��X�� �T<ol�>��M ����EK�<�쓊QJ1%�1
��r�3�}��.s9�<#����D�Ø��� +W������$�%P��'��w�^���pCޘ� �w+ ����`�9�qг�Η=)�=���y\	n�`[D�}AÜwa�����a@����	�J�>��y5-��s�sfZ����2/u��.S<t�[��h����`�����d_��ծ��ڈ����BF�.%2�
eAdY`Đ��>�(}��3����b��R�5��;w7��k-��uL�mk��$?h��h5ebM�>��O�T|o�Ƙ��+S���\=���d��#�7\&*˼��;�2��޶��S�q���θ4Yґ>�]&�w��s�T��<��z�|hG��tX��u�<Ay���������Vl5��<G�l�F�:�C��^H�8��w�V�0��O�/A����pUϳ(P�0����痤��
��˰B�&D�W���W�w����Ӵ�I�ɳ�o4�W,�ۦ$K�ֹ,�F*�m�*�a
o�&߀�>�/��4��"m3��峰oТ����޼�4�8鉽P�Fa�T���U�,ь]��?u�m��M�L}��X!-�]_�ˬR�����G�%E��{t���ց�ۣɅ��n�``e��MSp�MM\B�x��'rsfX2q��E�,��8�
S�f�y8��Ɲ�q������sؔ�Q�eI<:'_��Cw*0��v�`�l�y8�p���UK��r���:G
|����')<�L��ei�Dy4�X�(��.��"�#���a39HK�	%KH�f���H&�{?�^
��U��1�#-ށ��]E���|sP�H�wd�q�����/����.��y�� 4������]$�B�h����gQj�z�������D�W�*%[�w���{'�t�G2L-I/x��*��I�R�J^�F������~'�݆Q����FN�EH�,�C�`y�D�����:?��2� ��r
`5z��8j�qL]��{�t����/� V`��y���[�>��{�V��)�,�v	׷�l�(�Z��Jm��4��˽��[�nke��9��tc�t9Of_�}8T�N]|6�<��Ĉ������g�$�2 
���9�\�ݮ3���\��-:21�OV���O_B92,H�#��]~��������'�T�k�a��5r��s	��dy��O�sª�U�h2Dؤ9?��
�I�M~/���
d����uOcܻ��7��>~�&K��$��sצTP+M�d�ӺCO@ +&�?CYڙ[9^u�Z
�_eܒ/X{;���^�y����AP@l��~=���̳�N^-��'�,j/g�  �����Q&�A��&0ŗ�0s��Ҍ��!�!UҺ�k!�]J(P4�� �W��$�k��D��^���q�@�G�W(�u֩��� X�y���Z�Tb���I��Fh!1m!|���v����LZe�z��� ͑RI��S?hm7���huml�@/�UaF�I�������3Y!�7kM��0 }Lw�3��3�
(Yr���Z��\�l��f!m���V� 3��^����L���kX��
Ӯ�Zt�V,|ߊ�P�,.jU��iU-���sò�΢u�����7�<<�ME����@�8��@� ]��f"���
�����ʰ�I~V�ՏL�Ab��ͭe��l̋����YXҊ�$�{�zpT|�|Bg��E�3���$L=�Q׼�I_ma�Ν�E��v-�+�L��/,G�-�8�rD(�1�t��>�9S���i����5�Mȋ��Z��S�\����>㗄\YC�Y;c���YI������'= �G}���o���k�<�2�D��x xl���v�}:�(��-_��X�bql���̄mTJ�LJx�}la#�Xh9�	y�]��$7^&	�s�2�դ��y\MVc�\X��lH��)v��`���j��(�..˩9�js�I�bA�5ҐS�����ʞ���z��D����0�oL���(~�z3H������@"��u:�z�� ���)��L&���Ǟ8I;��m� ��B@%'w��+ep�W�4���ׄʍ>~/̦t�����P����u�u��y.x��wh|e��m|ᱧ�#��bR%�Lmq_�_�.�MM	�v��-�h�m��{F3`lh[��G�з��TT�ǈg�b��F����)�[�C��{c<V}�~�APS��Z�e�9����E�Kӽe�Ո��<��11�*_g���B������D�7�ʏp ����sqM�&g�� wJ=�ܴP���uj=o���S�jGw�g�ϻ[�����g z:Ee�p)��M%�Os�6�#;�-���§=��>�Vc&�l�=?�ޮ�p���4�����Юák���R͎�s��[���n��m!t�d���(���(Щ{��At��恀q�A��� A_�c������?N�U3��ZIq[Gi������5rv9���m�H�"eũ�q��c���`F��K����.�h�п~Hy�ҫEbL�ܩGM��Č�Q7^�����_ (3/<�O�����<�A���UB��1���q��g�����C7mKPP�K�y^�AЪF߬�����j9��R,t<��?^'��נ���V��[%��0�1�5(r ^I������-��yd��E�ۭy�G@��4j�5
d��.Ä���<��iσ�n��Kc��YF�AO�$�Z�����Xs_t��MB)�l�oZ�{q��hu俼Uλ�4�f��W�͉��_e�J��V�l���y4bj6�����1�S;�. )_Ӝ�?�[-�c�()Q �������?����������juA�y��~������^b3�!*�@P�y�g5���_�zϴ��u�� }ﲿb�w�󠬣��*2k�c�[�f#���~�4x-6��A��{2p<�@�^��E�zG��Sv���!�:��Z�\�����C�a�l�.����Ѣ���Y�`#��uVl�L�}�?�V�����i�A^�hs�b@e(�6�`j�Re)ܶ{riݣ���	:�b�h�՟@^�rs>��}v�T��]]�▬}���h-ڣ�����b �  j�%ѩ�ԡ�� J?a���IT<d��ۓZg>�gW�}��4.���/�:8���i�2�������������sc�^2������g��v�vt�����
u�mǌJ�۴<%z�p��vP�|U�/�t�p�HLm��~�Y�f9�;���k\;#T`�R�s��彘Բ&����Z��Hd`�KZ�`<����~s �hbg�4����86K�$,��&pK⣟ �-��_%D�Ѳ�*t�hj֫\���I�}#��p��pN�ը���^u�V0ף��S��u�7峒,��7r���3�-�֦v#�v�?\	�^�v<I��~*B���)�/K_��L���s=�sB�;��k���y��".���_��l�`�F$J/r��M��2�����TU�u��o۴�ɲ�ImV���ފ.'�(K��a]��d�|����:��X:��,��T��T�"��[�kd�ȍ���O������|�xm��o���`�i��'���O�4�^c���C�~�2띨�����?9�U��z,�s�Z#�9�
n�-h*�������q��,�@�8���Ԟ� �$n�A�(N�����/�r|"8ySp	U&�?�:&8;@]@CW1�ml��
"�xhxCLv����W6�n^&�䱣�*�]�����r������+��"��8���${��Sǌ����4��R�E�� z��[G�p��J��5���Ǹ�������IM���u�ƍ�_��4�i�{�v���]5����{��ߎo�.d���J`��X�]�;T�n���Ӱ�Lg����`D1Xh��Fׇ������CV���X[#��a�c0�}�kz���0o�sP(n�G��,��;�v��l�kDې��gʌ�Z���/2��Xn��ב�;��F�k}
_� �j��{`��Lo���x-�|r�_�VvL�[l�2�5qˠ^�F�z>4T\Y:�+�1P�0�t�Ռ�}�s�����W���qG�_�s�o|��ԥdv�V�z��Ӧ6�L�����q�+Z/�6L�Tڟ~�l��Q��!��\>�f�,���fi������>�S�p!VF���Ct�+���&�pj�,��+N���4�?��X��*Vg�>���3�->�t��	��m����Ҳ[q�G��S7�
Z�f�VQ���N-�+A��Ls$��k���[��Я���T�~u�Mo�:�i��!��Ib�ӧ]�=HC~VF]"[�� 0B�z��KM��M^�]I��ey����FuֈvU߬W��i.��)��8�_<����itpgoYD0����|Àv�;����Fb�d��a&(��1l�Z�tSJ�䷛���B��O����1��}{܊bX:m�T�q��^*
��Z�<$T�� �=3*�;�UwO��f�U.G:gy��z=\��c��qB�p��|�]�0mwڅW���T$J����&A���WY~���	���V�/G�}�7(Q�^_Uap����)��TtKݼ��	߭A3���Y���IH!��+��}9�
=��;үH�y��b��/ɨ2��\{�gQ$/��]�-�����<����������&MG8��L�GO���e�[��Q2Q�L�
p[���*1L�0�(��?5nS�ןH�@�ڎ�L�6�3�҉�{l�wk��`P�_T����]�g�B^
�>�\�W)�4���wz��X�g1��'�#O�n�� m5���n�������t����^T-gӵ˞�'���=�9m;�����%w:e����3� լ��3����f������Oq�S��ơ�Zf��I��k7���%�������F���T����u���3���6���;�@�e�)I��Ž�����X!cImpz�#���_��}���ş�+}n"!L���Y��a"�F(G ���-A���~����1,�O%��%P0/���� �A�[��n��SS�2{U�H�;*��l�!:,1	)�c�y'U��>w3�7�+e#L?n6�S3���ۧ��)���z+m+�	�b��)ݢ��1+\�v�.��b%�j��3�׿H�L��G��F�&u�Jiz}�A�dR[sYYK&�0�?����O��:���^�ב�p^yk���`���t�n��h
� �8�_Y ^	_?|�<�h(�w>��/{�}RЁXܴ}��#���2�q�J���*�M�P:�D�g�����E�m���za �n��uo!v��b�MA=N����c%Nm�TM<q 6O��؃�8Z"`��������Xw_X�R�[�S��Y�s>%~�(_�"�u�����)f�D�Ѯ:`��oPFϟ�q�AJzu�~��StXK<%C���kl-V�̇5�i���Y���V=�F��׿7*���tc-����j;\�0+rQ�Vo����m�������Be��K��fΑ5z��(�u�?��Ԕ��e���UD������+�_1��Ge���Q�D���ΰ���|��u��&�5ح��Q�T�2��bԚ��n!��/&^�o[�pU�_/�5`n9|�\E���⩵�?u�*�̃���0~�L�t�;�k�u�L�YJ�q�+B|�݈��	lw�����k97Sc�G��S�B/5�ba��p
z6���-ʦ���}I�X����GD
��~�F=�����9ь����*a5�ʄ�;J^Mז		k�C�p󌿯����ZMG�m��{��U ���feq9+���Ƹ��|��Sq�mI�V��Ζ�N^��Iܛ�!�(u��԰z)�ǫ����5�n-0�A��*Ә��k4ƻ>
tʆ���6>���\)�1`��	�%.}�+��̽(��ϸV&Iݩ�g�����&�KJ�ڻ��4/ �5��	-�`����&�/�'�γ�W�p42�?��.1�оp/ֶ{ٸzP(��qBn}1&K[ן��滞Y�Z��*�&���!f�/�H���h���#�$X�&@�����=b�7��P����/q.&�0�AKGH�GT۟Kd2�r�d*��,��Tf�fk��:�Kq�Pzظ���]�M�05�`���f]I���Γ,�X����AS���8�L�%�{���uw�>7%�2`gy[��k���ᱺ1^|��B�=�@J�-Q�~�ѣ�>S�ƴ�����V���p�,a��o�.��#$��l����N�բF%�*XNnk�n���Z/�[�S�)	���GS*��"��_�N�N�X�U]������1�YjBON7KBL����
,�Pwm�V�(B\���WL�o*�����~v�ʡ�(s*�C29Za�'@� u}���Je�h�W�<AQ��VZC��= !����vy<�֜9k��m]��iO��d��:څK ����}��/КP�X��6MГ�f+��՗ä��Bʳ^�+���)k�0;�׼�p�i�.����S:���h?�j��	Wܽ��j�R�������	Z�yiv�`t�PΕ):PrC��f�jw��t����G������R�BR������r�s8�=�NN*<�j�{sA���~�	Dtl^�DB�z �j��#�\<ܨ��,/jj#�$.;�h��G$M~�EL�(7yBul������aݤ��!�f�R��
��˷�3	��T/�����1���|ׯ@�}��Q.crx�����Nǃq�!!��lh��p��$iEDq�T����\�~���_�q�v���W"R~����_!S
1��D�(�Sn�{H�ӟ�܆���)蚲x��*0�kg�B���j�%���5�`>;#(�� ��E�[GE��}ã�(�GPA��.��T�K�CTPRIi�f�n�k���f(��70�9��}�k�,\�g��������{�"�����	HI;8A��yfa=Щ�Y$ku�6ZN���f:�T�,��^=9׍�ekїM�qBٿj}&�LV��ք�oi�4��{�>t�^i3qo�������E�Z�ߖ�v�ݠe�~�A&~�K�Ӂ"�@�_���g�r.�êY��a������h!%<������J�@��2���ӷ���B��d���T�܁F�8�he/
F@�ad��e�����Ѳ���Y�RtC��B@R8w4RZ&��)�`�l���޲�=���?�[�a���9&����j���K�����5�
�._�K��/����G9:Nbǩd�W��㬯p� �����JC*�v�0�9Csq����-��~@�Q`�C`�"�ʲ��%�K��,�6�=�v*�V"��"�i%�{�"�ŁP
�fA}�S��QhlL��}pLv��xӴ�zݎÅV��,�oQ��k��~;\o�
����o��
�P��K�����l��
�Q:�<n5�&�B���������<|ĕ�4�C?n ˅�i�
���������l_L�"G}5�4�ԠJs�����Ƿ_�3����a��	Q8��J_*��Mp��er|OR�z2���OS�+�6��Y B����:���ҽ*���cX³��*K�qՓ +���>}��]�PI���]c|<����%i ��sCI�r양�rG˘F()+�L�U�f��a�����T�ڊ��k�� ��O(�A��[���e/��o3����s�X�*�^�~��Z���u�d��x����^�����9*K�+��l�k�������wO�5��OV��eZ��D(���8>���?����kۣ~�%c �g2zw{��U0�-��2띴�کP%�h)�.�2[����ݠ��rn��c{��n�5�2�mɤԧN�d�,�z����W !2`�w,�Z�z�],���s���]�T�hu�p{�h��LpI#�y��`�::�B2�5��<w�	��'dg��y���f�>&�:M��+��M�g�Jz����y�+U�X|��|�f7�{cY&�Co0嫥��2Ն���7m��r�L������@���+���`����*2=Y�R�s/��[�\����]y���2�$����%r�\�8�C��{]4�����_��.����Tl��E�?�t��kRT����M9��QT�٠��ց�9l`d}S���3�&)uF~;��f�s棓�8�~�j]ʝ�,r)L������ƞ6���5���ƮR�˫sG��W��P,]m� ��$W̿#B��"���H|�4�l|B��'��>��f7�G�+�S��d�z�+l+v�V��Zb`�i3Υ_����]���_��ת0[���:]��3�~�X�1K�7Ɩ�j���'�e�(��/3�Y��q��J�-Ixٝ�,*�Ƨ�`�$���c+��#�Z'@k�,!�az[,}`KT�E�nXQ����x�-&Ma�Y%���̓Zs�4v���,��̍(rV�5N%gؓY�5M��!ߜڛs��{�q�-ľ|���D%Ax�O�<׿�������w]5qK���q4�eTdW��gʆv�hޱ�����&��$y+m=B�yػ��h�qiFR}Z��xA����5�_� ��9��Y��g}{N���̢��ʊ��i��X�i��pt5rl�In�?x(/@u���:|����!�}�W�[y�Lbg�/Wxk%�w�����̚�,a����-S��.0��tR�]�;��S�\�D�"J�ܩ�Mv��؍�����I$.
���rdؖ�q��$�{�25�b��KG,���r��q+��3��<�fX��^1�L��|�O.�
�mq���J�6�2ލO�SA>E-,��F�-�~|�q����.)P)[ٳz����D!@f����m]���  ��i'`D:z���k�D}��a���prF�h��<����/��|��'�I�+N�DSؽ���Ʒ+�Li���!����۽)<���^'�
%��ɝ�yǎ3��O�P������P�'�Jn�Š���&YvjQ�c+}���T�sp	��:�������6����-yr���8/B����-�0PG){ �C�5fɛl!���+��vګ�j&"��|�����#��K���#Z�y���i�L�W��� ��t�5\�y�i�K����n �j7���� �ѧ�ӧ���ܘ���d�'�x�f��$�P�{S�"�X�#5A"h>@���z�����T��(���R�vv�L)�lٽ�d�$�.k�3.!���(��.`�c���X:{l)%������ӎz2���޲T4�#U#i#"��?:*=,��aj ���G*6��:��51G<S�
Ƴ�7�WI�^vJO���+ը\���9	8JwĿ)���p{������,p�	c��v��j*�,ٷs�M�=�y�5�M=�.��.n�6��ql��-�Oo4Y� \Ĺu�,7[~<z?J�&�� ��
Nh�AJ��\v�̦Z<�;�8���]Ł��@�[ۻ�
����ӓ�i�\���1�ffi䡻��`�(7�,�OD��l��썹� �v&k���L��g�h>�3z�����U�#K���;�B�W	�5�&��Q�1��S54��,�3<Ogx>��!�6�m�?�=�L$��鶔5>{�Ǝv��(/f;�b�Ł�+�xA�q�/Td}*�ZH|�<X�	?�a>�z��N�c��~q��%O����&C�0^Q�N8�	
td!������PH5N&���q&��ᏪFU	�&�XS�jZj�H�ko����.}&I*���!MjQح	y�:��&�a`�l�,�1��G���d���4S1,,TJ��	�*E!����&�J�"�E�NF����P�S��%	5��7�v�Ŋ"ڢg����6�ǡ�y��˒_Y�t-����6ˣ˨�(>�pE��G�7Cw�-�����[b�*ܧG���3����;>%�MA�(z�I��/�E��P��|qP�}=�I�9��ҥx�!�X�[U�On��ѭz�gK{j�P��U��Ðwg}�qɝ>:�Ď�8{}Nx��N
��� F8�8�ꚨ��(=�Q��u�$� ���+���~YG�����#���ߵ�w8`�4��5SҒ���c��׾���u�"MJ�0����!�.�nȇ� �Y�^1�/�G��y��^��8���w#��ӹ��T�;��ϙ���dE﯌���ȅs
XTНB�u�l���/dq�zi����فI@��͛O-)�Px�W�P�4��[�K-��i�?7��_�TUBp\��N ����$��(>)]��m�0]%�,;���SE�R�Y$�G����T8u�'��f��(�fĐ��mGL�5�01��}Z��f/jxw^zȼ�$@�|x!:>�č!�f�O�z*�L���3�q��N�!sy �*z�	{�Y#͡:�u����<�,k�+�>kmԭ��7��2/�#������.�s#ObA�6��o@�.,�E{��1[ �f�YXO��ɖ֨��Aw��Ŭ�#<p���W�R�s����A�9�قKL,��NE .!�l��w@x抭����Ԟ�(>r��s �爙�� ��8q����\9j#�{6͚���2�z XZ�斛���_�L��M x(���xo��@������W6�Tp�6K�Iܢ۟��Z�BJi0Ӆ�ղ��"tֺ:��<�ϓ81�?������"3�ݚ��uKCeMI��*����N������>YZ�2V�?����N�%� <����VO��)��N	�7��S���p3�����q�L<s���G��r����^���`Y����|��i��yX|��C���(P���O�|�\�Ê:6��ѭ$v���e��6H(�d2~�u�Bz[,��QU� �B
��*$�a���n?̷=�0�%; �f��74�E��d8@�Lm��}�N?��k.xRT�HsX:��1/^�XR.�mz�.C����;"G?�E�Nx�C��Y@b-�%�p��oŐ����a3T�J��� `�!^(�\����½��Ul�����mȱB��q6�n���P��X:�	���B�U;�/F� ;f�*�c��}޺��𱒜�5d���8���8����&;)�CY/���q ���
~oki#��8�X_����M��F5z�j��3y��g���{��]QU5���kM��d�Z���m��?B; �@���={�8|�"G3B	&�\�_�q9	�ڧ룸'�X�^J_�����U>��7+8E9�Zk�/��>b6H�m�]��=G�M���O�z��JӔ/��=��7��`�}13�ؖ�*<���0h._֜�"D4��H�O�병<�-+ ��[�s��Q�N ,L~j�2[�"��58�M4G�׈���Bl��>%���ӭc�^�_J'rd��ۭ����6jQ��H6���G��,J����`���fg��F<��ī��Z�R���&�+�\���&�9�
j����<,I��s�o��N������ڭ�(|����޽
�������~���Q�Y<_��պPb��h ���ص Gzh�Tqf�\�)��\��a!�n����G:�h��守iD��������Z(��(��*z/����:�?u"5�:���$'ݓM�p��k��UN�w��>e�H̀��r2,���0���P�vl�]C�}��vyB�iz����`/or&�7[�y:hwS�y�Ez!*�\N�dU�ܗ�o^&��,��~5G�ァ�ݽ���Bi��i�Ç���M�ʞ��|�Օ�����JS���}R,�Te,v*^�R�D�a��^V/������֥I����+s!:*ʳ�-\�3@I�6Ә��ЍzvwO��>]z"�y���{��z��h��:w�na�S橣��x��Jck��D�S�x���d�����+}U�Sq(��3����R�6�q)liE/����p�VZcܺU�OaǑX?�Z���k� j�2�08U&0���j�O �p�*��}p��̣Q����Fk���W-2O@�H<3}����Zޖ��{��O�),V^���wy�j���Îp f8MPVv%K(�E�2�tI�`��c��I�����p�Hdn�#�ي����4k@kN��z28'����Ie£��� ���Zah��I ������=�}�i�.�� δZq��T�E�i���iO�L�t.�h�H��eqz)C�l�.��t`n:L��X*�TE֙aH�8��M�*ѡmi��ӕŅ̷��jd��@����\��D�%S�4�ſ�z�����CR�����$�O�.<}�q�Q���8�K��<��}[��QC���d��\�80Z=�F]��G/#;�׾�ح�8�30.0������v�'��3�2n�t��V����+�p��.'P�Acf��DPrr�+2�D��'��z�!����S��.vKRBpyHn���:U���-D�A���wu�h�i�n]V�|���z���A1���WZs�������o6��ѐg�"|���.��jY����B�A�y�~��N���ϱ�CEs��~"�@y��?��L%��\��T��*��w,�f�D��)J
����� �<��
S.�M��85�:-�ХD�7�9��R��W�� �w����L��p��I�}�
+Vחɫ�g�b��נ!2ܒ~uw�bv[�bG���qN����s~i�W��jD���G���_��ò@�b�~F��}����r�ۧ=�#:�%"׍�g��L'�����c��b�u��x�7�_�
�47�PIZ~�]�`�*��R�co��P�*b�wO4����a���#�)Mv���;�k{�fzU�k˜�ᬭ���!�|�S��������f�v��c���h(C��������j���Җ�����퇿n� �C�-Ȼ�_�k�hsŷ�b��#�U)��-Aq0� ɽA�#J}�1r���=���@�u��)2F|����h}'�/{��)�_������Hb�a� ���X���� �]���d��r���I.S��1`>��r���*��^�Px�ƚT����| )3;�/��O�N��+����*홑C%L�h�|�z���ik��<�W����r�Z^�=氁|H���R��a���?���~G��C$�_ߥ�Q����\�9s�%ǅ�Z3�~S0eUG��۹//`�[�������E�ݯ��|��S�#|v���iKS '$Ee�A��h�K�#�-��!.�C��¯�t���E�,?���=�W4��>��R
����RI�b����R�epB���K��)�����Z�w ���
S�-��l��N�,�
ue�難��20~���a�e�`���$�^"L���T���������a @��

�ឩ�w�hd���M������!/���s�?^S��P08��\[��r���Z�}߼M��|
����q���RdnY"�[q@��q��T�������B�Ru9��x���J��y��v ��/v���ԖP�\�B��� �t���Tyj�b~Lw~ORm��2�z<ų��e$��� � iW��c��I�V6��A���Y�R�4��%,�A�Χ��6�Zs�~���K,y�}�]+�a��Y�& �̷Z?4�W����$h�x���N��!wG�c�Ɓ�H{C}eT%�}��R���n�I�[,α�9�<��K0�@Si@\||WC�i�s��d���j��Sa��E,	�ʼ��v�'���Y��}yq�>�M!d+y#P@7��s��T���%���X<V3"��z����4�A�P<��q-����o�6)����>�|��|�ф<������їp���b�	��-a4�SX)�}-晢�(t���m��Ed�P4�	9f���eK(|RL����bĔ���F�]W�ࢧ;�}#�-a���	ҊoŘOwNލsh�?4j:V̟Pb��`��P�y�+c�b���H[��'��}�\���NKi�4)��F~�$����z�̟'Š��c���l�{�����:=�p���N;q���,5��0��p�OL� �L�y��������!%v3����kSV�g�I{��ʰ	���u-N�3���j,��O�M�,����9�$�X2q��+���h���9�Z���l�ՠ�{W�Cb�\?Lw���nd��!_����ً�ڻ�d�.���G���X��Cf���aӝ���k����S=W�y2<��7�J����vcG=z�������Ԛ�Q1���%`����c+}{~7�6=��Ge��+��_��o�(�r�rS̰!�y�6�����b�,c�p���|��«�ˀ;xh�щ���Y�6Ou�E�-�ͽ��(�� �����:X�4��%���i_�|r$���7�Q����D�T��6jnK�*S�Z��;݊��= �y�֯�X�+w�ͻ �#��={p/cz5�oXiN��@����_��d�D~=*�=�%����ɩ	.9$HK��}��/֤�l\�5`lǪ��Q�9jڏ�f+CrP~3�o�]bsQ��y\�gQ�ف6�5��I#Ji��cY�VC�ʱ�Z��Z�lFӜ� \kuc�\�����wT�n]�׼�z�W2�T=���ϵ=e�؈�F�-�`�S�[�L�.w8g4:���<����O���ܴ�0,�Q��D'�fB)�e0_��*EEEB����9�YSmg��c@���xQ������y��*�D�����P��&$_����L���L!�J\<�B,/����]1W�Co����2���nT��C!'ޜE��b��-��b�U)�%�.ӌ���)1�h�FR�~M�y��(�b9-S^�v��O�A��_v�T	������{�2�l#5�����B���˓=�^�丌���Z@��S_˥�eg�o���_}�-p����|$�>����<I�K�7���k�he��&_��{�!А�Y�xa�iU��2 wC��;b>�r�s����Le��-��ݓ�y�(�_�e�� e�L-�TnH�����z�ד���
aE�,��k��n""�FA
̓p-���?1�_��(�9�r1w��i� W�Q�`Z�Į]s� ��E���\� *)�B5 ���C�h.�$����l�\�4O������E�EI�Eb���8͹'=�'HE����"Z&3�&�ёbS !@n/�@���t�
J,~���f- ����u�� �z��f@ڗ�nsqg�c�2��� s�������+��TtM]CE��������a�λkFS;j\R�+�HIW���>�%Y�b!�m������z�M,�c�^��N3��B(h���ʹQ�Y���~s/S�&�S�=Uh[�I;z� we�g�ف{>�ҲO(.��T�*u{����ϙ�yj�Y��2`�B�>�&�R�ck׶��sX�TliA E�P���S}Z(
8��4砄����<-�c_�|<Y��%����G��T]��؅uǡgpd��ݧU�E�wjc��'�ι����#a�<��X�'�$XN�&�4�8�[� �X���n#������rEm�_[I���3�t"KU@�6R��]������n�HI�8�0`�|�q6~.��[�8�O���VF�c�ae�RT2�jh�7���\�0��uf̀���e�u7�ϗ��A�t���ւ�+�pR$�ʥĐ^��A��9��t���\�{�2�h�G�Luv��2�/^ty=߲l�'!X:������׊���H�U%oW.�n�=Г<X��nUQ(��*^tٴ��J�༼��Fe��W�08ja�y��O�K.-�;����s�N�� ��Ԯm�?Z��}�2���A���<u_�su�0XxH/@P�nZn��ӥ<t��{>Hr|W�@�0��nH�nxOo���>����(�����TwiƗl\��O2���֕m�B���gX�:w��l��D�|��D�zd�I�4�V���&���H��O�$�yZ^<Bo(���g�����\��@ة�=����p�J��O�T��2ܪ��V����N���E�RY �/�ٿ ;;�fou�^�z���bkK��N25;;�	�X3�U���#�5�+`ܱ5��+�W���F
�7��Q�Zۘ���7ߕ�Yb��N>Nt;�\�r�u��HL�zU\��,�<f�@0��=Y�δ�r�I��|,���)��L �8�9� ��⤰�����1�Fw�"��I���5ϔ�P�-��K6�T�u��X79���&��U��U3�O�VcPn�ٟ�۟�@��w�VQ�;���sz�XX�R�-�F�5;ީ��t�_��C���nF��/��|ѕ�=ةe�^�w�D������?O Ǳ�/W���%��!�ð��~ �o8����:[c.=�}KG����h<̈���t^Fq�c�����"w�c�[KY��/����������s�'�iD=����Sy�Q^9�n2M��сJ���������m����>S�.QZsY	����,G��֊�|�;b�=]-���T�b[�0��0�RX�ʰ�A��ی��޾w����\%ɲ�')���7�
��@�&-/����6O���Kv H�xR��o�\S�1ބJk��}��B^�L��Y�Th�騰�'�'�dMi���Wʐ(u��&�$���JS�fJ�ҝG�����SYLe� �T[��s0t��C4a��vw_�m��!˂��W �`Gi%7�2dQl����ԉ$����@���Cko�z�șy�s����W�b��~��;n��3��� �ߥ����L��ô���X�!�I%�3�8{�1]M��.�|C��O�@~e�B��I0����ed`��Ȟ)�b���88����QӼ��~�QN��n5�ޝ�ThA�(RV�,��^�qP���W���R'?58LS V��"��@���Hgb�O'M��RȠ��+�yY����:k�Ļ�~js����Ȧ�su�;�v�ف�l�3<�}�yi���*�:�*b�i�d���p:�ȷ�'��$���U;�|����T64LC@�g�8{5�=_��h�E/�JB�u�������=����G>V�j"}Z�.xG`oD�-m+
t$#���������S�>��>y1����dLR��|>���<�#T���h�H �	�����~�ӧ蕈�2��%�j��/3Ŝ����0�yŪ٪�c��4'1۷�n�61*�,��i��c8�A"�v��p�����2���EW�
���G��bB��C�;�����	: ��Ju�����x���G��FA"��i�z��wN��zNN�g�fo��
���-|U����6�g��Xr�⃮qCc����~r]��i��<p���<� Ή��:��S��nټ�o�6 ArE�� ��I�M�?Dh>�T\f�S���)9!Y\D#ra��dy����|o�#�R�:�Rj�3q�E�	ъ(�gY�BIW��!!\y�	�PV�6���6���MZ���Y�R�J7$eb�Kx�4�q)b0tK�bc�d6]9�{n�g�ơRG���W�t��/���IL4����I�3�lf����W@��ϴ9�GWkx<�I�����:k`��0��О�{�2���m�W������P��� 5��>Ԙ�;��SMa�u���O���0��޴�}xݶ�� ˺u����[��L��q����$�|���71bc�Ů��x��x�#���n��O�8֛`�?y����^Z�����L�$u������q������7|_����\�Ƣ��(�I����+�~��R�6#k.�s���qC����>�F�ܬ�g�F�G{�;?�,�v"�	9hdÖ+@O@l�U!�R�\�>�7���c��J�}[Ǜ��{����;�Иj�P���[̲��I�.�!  hLԒM�r�)�Ch�O��PȋN\H�i���l�T�qF�8��+~����L+c�����/+|z�
D@�U�P"�`�=~X�4�(�)���r5�}� j�:��*=��U����QI�>���G�~��
��b�Ο�)`o�ħ�[�μ_����p�LC�36��N�h��58�(�x�ڕ5�peq�ݪ5v}�4 0��^=0)�F])5���絿��db��������+��u��Qx��Vf)~W��4#U0F��te�p�J:�6��f�K�Tf�H�;�\�����b-�b�6�K�#� ��nF,���٪�p�m{[�e ��q��s-�M�^#�Q����g��ϧj�n�U?>5��Rl��	�4FO�ᵵʪ��M���KŢ�L��^�2]�T'ya��9�,`}'��8���E�3w<���T���W�V8��rXG� ��/Іve�Sz*��5�N�x���q��(�N�*{��Ry��M�%	�{�E����P�78�����G.C�r�g��(�{�	TH��
`���]����{̕U���5D
��DRr"�+Dz����w"��?��5�G��Gk�Q���u}���^��}UX�����q���R;�iI��9�xhB�D�&4��'G�EG�*�'��N��L��'�+���;BdR�D**Gu8���EHN��]���?��}|3��x��Q���I$f8�V�	���	�}���x9��a�����q�Mh�E���"�f�钔*��Y����
݅=ۢ_S���):wL�֪���ejD�~�d{��~t��������l�)p���li��Z՛����-�T�3�_�	d'`��R�˞J3����I)|�-�c�I����������/R�q�s�����B����N�Y*�N��_O�b�������?�I�~�1RY��� ����m`��g,4g��}�0t�謙}R���n��]sYb��n�,���CD�H�r0_������ɛO��]��B��u3���k�s��s���3����Ƚ����P	����Z$�T�Nі���T-����C�L�#Ϭh�G:L2�$�b@=CJ�}�v���V��˜��Ψ��,G��?��pv	h�����߷s)l8�z̢��P��y|��~74�-�k�e|G;[���W�x��z��KGC?fQ�"r2�
�R�n�-�R�m���f �����= T�|=R��%黅Gԉ�b�֊H,�1���ق4�������sJ�",7�uDh���j;áZ<�B�@�3�W�#M�h{P�E+� �V�l�N$1���,ӰNq�m��A��x0��;WY5��{��ʨ"����Ș�L�DP���U�s���J�(+�PV�=�C�b���˯<yX-��-ĘuKz��te.�((�&>���{)��K{1Io{#�0,S޲h��� d�o'�� ���$�ƀm`�����!�'F��;I� +Ņ��~nS�bZ�5��(�ڟ�.j�Q����?g�	V�ϫ�[p����"�3��_����"���v�J0�]��Q�w�t���9	�W%v��#�(�/Ei&�q��)�i����0Dȧ������aO�3�8���۲M���[�r�;�������L��<�|�4ϧ�Y�}I�jօ���Z���Ή�� ɽ��+��UI=mͻ�o�^���������l�r�g������\�ԅ�ۜ�L�S�0Y�SIl;� ��O=�p�T�vǞT���rph��OAf^B��4l�Ot�t�?L�M�Wa�2�"�Z+`�a��}���4����v:8�cA3�����V_��gfg��2�:���"�m��qꙎ/U�� �6g�I�ڏ��锇ʿ���$�j�T�vntt�v�3��:D�5��-�XI��\I���C��E��N��B2���%�]!�J1�rN�슥mb�%�~I���0�Y?Q4mm�Z�]�^�fbz�d��F�ٷN*��.�N����]i�h:74\џ��}���g�6�Pa����;��1;/��LR30���x
�?�T�E k� h),z4L��Zǵ���=/?^k�I��>�;٢Ƞ(�f`h��
�A�u�2K̆�K�DEEÞP��P�3\'h]�� ?l��>�μK4��[�z<�o���V��X=�|q��z�h���������g��xR��q����n�_-���E��q}��4�2#�Z�#��eK{=�h��=@|Ɇ�Q�S|�P��|�\T�u�����i-�vp(�n�	�gRcȭzfw�{؟+�-^�E��kʹ�||���8ǉsv�e���|��{��9Q�f�� ��I}���%��Uʃ|�s-���l1�p���w_�d䶱��8���F`�K�AO�u�ΰ�?y#��ܜ�`���,ex��h���hkn�� 距�JdK~�2��t_����|Y�
l��|��v��!!���������?�3<l�?�!a6D4��&x'DF0���Y$�wp0=-�9S2C�������ɫWihlD��̭M�����x�.W�԰�<,Gon҇4�����cn>�JN�#�ȶ��O^�I��W����
"V�'r�'�"�,y?@e?	)����XU�D%YŸ�Qp�ؓܐ6�H��qJ�_��l��[1t�:�ͼ�+;�lt�v�v\! ��M����!�F	cǽ��2t���`���8�����Y��r#�/w�Ō���q��Ź,Gڇ���j��	�F�/��V����;�/�ˀ�|�Ds {O���-@��h㮖��k�xR��R3�r~��W�.I�4���{��i�'�=�iX�`Z���=��LUT�Hc.�:{A�.������ׄ�l���^�U�r����W�7�M��2�J��z/|YZ��F��h4h��
�\�2�GU��V�j�"RRRi,,,2<�Č���	lw���;� L�v�>鈑�H
����?�z4��h��֘�d ��b���L������&�m�3f>-)?�*��٠�W��ܜ����ν�Y`5G�K�z�xC2�-J�nE�OM�a��5adj�е�w��7�Ae����)���|�X-^/2�}�П}�QV�G�(B���q�b��6޿�f��{moC�����]���R�ߧ�!�V��R��_yfcl>��,S��}��g�x�D"-��8����l.����x�귆�B�\���.�<�}����/�&�T���t
pg����LLL����#�H�q[H���.z���gT�:�ҥ�1
��]kW �"~WRb��}�9_��3S�����.�Wy^�劖�����Y��y��ҥ���n$�U����J�6ЈQQQD�;+**��{�Z$�������
��#�����!g�)�ħo��%���$麂�Z:�hO�÷:^V��H"�Vu� Ӕ��5[�R�����@]��`5"`�!ӻ�X���n�8�4����?[����8��L5���V��n����������%f����t�#�AL(^7�C!pk�sQ��c�z������S'�"��^�FD��塎���W?�.��c�q�p��{�o�׮Sy���i�@x�*ig.��GOV�7�E^�Nƕ~�&�Q��)�p�q��������T��&777�"4|�J�'65X���j?ʻH{���Y�e�xWkM�n�����_�p� $����!�`0��,���}gº.0��kO�V	��̱�-tV��$�[/*�J4F��Y�ս-J0&��M�i�p\���+��Jy���! +�:����P�T:r9-�^�l0���ɖG������;���׶��*$W��H��qwX�E�1Ͽ��J��1��X�j��K�{�(-�ݹ��?���C��ф���gJ��� �UN��_���lsqh^
yJ#tC=5D.}��3BZiʽ9���������3�r��"��^Z"�F 
��.fH9�*A�-���މ�x,��g��Vjv <D��4�������*=�'��;蜼63u���EIFn�����W_����`oK椧AM��}���h�x��C��g��V-ti��.P�8[����B �'TUU�������X��>`ͧp��C��!��F[�$����?�R)Ӧ��6U*:��:�ӧ[9e�<Y������.�]����%�t�k���`bN����]B���O��E��/�Y�Z���L�S�\�~����r�lÐa|,8�Q���?��z�N�=�3F����Uɚ�yMS�&0��
0�(
��_�~��1��*:c��4�62&�4	eM�B�)��7��S�iqd
i�R�������:�yԹS�d}��sr���m�bP�'6zed�1]�I4_��vRTS#��q��%w`��|$/�_BQ�7����gHV�8��f`��Y�!���I �t�{*�'���iB���"�'M���g:K}q�l̷�ׁT : �G��e;˕��Y������!�вWR3^�_��|���=k�/-�z ��ے�����2g[|�{<���kk;�����&����&�z߼/X5�;ԩƆ�=����n���615�i-�/]�Ѝ�.M��jc�#��}w5��:�������'�T�_�&��v]4�:��L�;�`�̤�O��Zo�nL�� #��|�>95!�FN�Lԡ����6n�Wv2�u���1���C���y0���m�,�V&�P�����z����n\*L*.�\��>388�W���e��{{���T[� E�q�m!�R���ZqQ�a��,����j�~��e����7�s�7�w�@w&[|��r5$~��q Y�}�E���e���QaF�ncUNV٥4\A�Ɩ��u�0�-""bUO�����Jz�w�Η�6\���Б�N]���շ�u߿��erV�" �#%B�Lgw��0��r��W=����{%R\����^��O)$0.d�7�:��l�-RNA!�����I�ko{zz���4���f����#��(�J��� Tt�GƄ5F��}�	��Gcyi�?��Vio��Z���
��9Y�����4��yGi@�7&,�K=4�};=��ߵWm"M'����Qh9�D���c<���u�����1Wܑ�m2(<~��Qz���M5�$%$��i������oՂ�̵�K�i 	J�=j�����A�8�*4l$�����@�e�x�0~�1߉z��#"Ybb+׵�xP�����	�ZX��Ht�J*y�@$��z�t^
�mZ��xA  �!����J*Z)#c� �iX��^-��s��`�]D��������z�]�44��ñ��Cn��I�9��Վ���^ /����a�o��`�l�z��6)H�/?���f����z'-�o$�ɭ���R#��
1�rphz�����L����g��7�f~�% ��u����X��������I(�[��.�f\��wƶ�}}}n�;ȝ#�<-����Qy��РZl��J�ų=:�z�E��Lrb�Y�������Ttt(!��;g^x�ޟ����HyFV<C�K�b���%!Lw�D���s�Ѵ�r^P� �T�޽�!`�ehx�c�/���an��i��GNS�O���Ó=,o�dO	귄:�7!t�.��&D�֣j$���y���J��Ptp�l�yyw[Z[	#q���6��[���w��!X],��Ȏ/R<�,r�j:L�S2�V��m���<�������N�!�~��WPP �;444����Y�s�F�^���~������t��KJ��!jg���;GHS��V(��o\]���P��5���Wg��KKgdg�����̯C�	�%���*WF(�6���ޟU̒TS���q]t��Z�+,�/tFq2�H~|߂��q����5��񇌁��R8Q�cz�S����v5
���)��xy���:����1�0|͢�&�������fm1��a�!	ߥ�
@y�V;����^�ם��@���
��溍$��C8�4�K|]�BM\���o` |����Ռ�Q��EC?�yϛ�-;�F� SRR�@0EA����L�����2��p�Êi%?��n�!���!��}5%Bx��b�����ɷT�O��d��������z��F+8�І�Q�aaaY��؇��X�|�_1�c``�.��d�r��^��.P8�%��������Ei���|A
bLղOKs5�� �8Z�\�F�� �
��?d�Ks�7�,tl4���]�I��7�ފn�_� "`��w�̓�xGlO�Xh9�-D���6��uK�Է�k;쬤�4Z�l��k$' N��lqq�h�6��Ҭ����	M�!��65�����(�L[����㝩����֏D�xPa����:�\N;�05���GI�f��V�tyF��\�95�#�8���@�K��>�s��+�;�����)�I��d�rs�cKV����Z����a^.��m�r%�B+�a�j�sii�[�����W �6���.2���=���l��RaIq"��;�G�O��x~�58�d+"�%�U��? hM�M���볝A&������y���+r��o�O��f-˺��P���UD��Fo��k�=����p,3s��Wܨ���˳���W�lI��
��0-�U�p~�8i�Lg||�P}���恣��1pq���Z}s�$��[Z[g�wS���%��;+��s�w�-�;bڥ��R�N7�,}�Y�X�:v���8�����ӹs�׏�+�����,���箋h�1Z���Q��'im�y�t�uZ��C��qCI'��=<&������-��*i��4�gҰf�L#�����@B�����ўX$����R��ܷc�߾47�3{�I��u5{r��AߟS��ZiIC����TEho7����q����_��kw�i)��N�f�������k��W}��HQ��R��⥉tiB(�	=� �NP�R���AzQ ��[$�WCI��?'��_�b)�0sΞ]�g�=3.=�Qt�!dwx-����P��{r5��"��j�|�AX����Yj�������kV���k�e�),X_`�Z4Ғ��ѐ��t���ĝ�`�^�����ƾ	V�����_��2��j��>:
��Ž;1�6���V=�\�ճ�G+� �5a�e��Y]]]k�������c���1�7 E��0��*@�gK�e�"h���_�
G�4�4�
�����Wbz+����P���:ry�9�������7u_n�f�	�H�L"���v-������1(((�S3Lz�� ~�<�c��oXj�������r����yS�|�=f�*�����k���/�l��7�9�W��^(Wc�&�U��#�+�����`o7!��46�̵��w}�����pU���L������xP���*-���!��,�%���`U�C[�v�~�p�"��<��^s��3%���[PO8�^�{٩����/��<�ޟ^�k�Ř�z��S�f_�����]oy{\lz8�/:�:-]zQ�|}:55!T���ƖY�Gy�A�=�C��+�ڔ�i�Q��	�lO̮����M�m��>�lK�_�P�Y��+�J��5�܂���3N���GX�h�)o����<C#҅�X����b�go��˗!AɖC��ۛ5��嗩g��uI�}�x�����YO��a�L�7�4*�4�LA⿂�7�����,�`f_�PW�ќ�b�����2�OF�>��- Z_KI�d�>9�a�j���H}y��!$���+O�0���N��A�۲��0�p42A,WVnoM�+-��зρ¨-�q��9�d�����M9`��-�����
O��o/Pt�F^���m圣ߴLX�52�,��e�k���Z��:z.F�iatA�4�z �Sz*��?��r�]�)���@�Ԟ�~���ߣ�m��%�����ޮ����f�/; �#��e�������2�a���o�^{x,��΅<P�n��a{��~���&�\P7�������H������)8�*�LsJ�鱺S�~YsH���K�k�!1uw�i��n�ѵS��_𳷺NgU-9����AMAM e��U]ӥO�Ԓ���P[���V�����M��N3?ۉ���>}��*+ua���+y�ֶ���h����kc��nY�Fvn�f�-�Llf��+�7�����^� ��v�����_:�p���bO�!|"oG���t���{�M�C'�qg�-�p�m��kB.�}�u�����</�R�,s��0�o��T%�� /Z1���L��VJ�!�`u1W���U���`Y�b��]`�_.�a[��o����5# Ă��	�G�bw��.C�6��8L��MFM�y��&&� �TH-�h�ͽ*&��!��ÙL͢������Y�n��:�u}�ׄ��RZ�4�, "�u,T�55��ĆR������_Ň[�h����9Q�C�\�wP�w�c������:<����|�t������B�����[��� �N�_������c����K��=STYfi׭�X��jv:�z�r)M:���tz�!��lU�A�÷����.[�v���e��k���84�0lU�0��穝ƴ���?d�A��
�tH`�(�_����튒4�I��k�� :rb�ѷ�ǽY�H�L� ��e&����|d!��.
�p���J�ysWˮ��PY��Px���P/���Kq_n��~3@n��~N��pM6�#+g{�[ʝ�%kS�+^�t'�4F*�?4��1ʠ)�w�c����!:��� �yI�0LA� �x�K�Q\�.����Т��b%��������p�6y�`v_�R�ߦs����V�5;D�,'t��]! ��FV��D5���p�0�/4����fQ���+�@��M�A�
�[�x�iS��2ɾл�RQ��(zѱ}LD���D�Cs����� ϩ�mhg1����T���hy�׋�L`��_n�k�Y�0����S�k��e�����:K��?��4珔$�F5;0�/���2��PG2�L�ݓJ�����*?����dz����cA��ThX�R7�VD\\���锝��R�ؿ��N��7�Z4C��p��W���j����Y>`��;�{GEE�i�-��݋� ����6ճt��~�~��l�ĩ�[o���`57dr)X�5��2���� �!��J�܍����]�C�$�����iW�����q�^���zp��co�e�(������*q�R1g'M��+v�ۊ��3|����yNj�^���U�������M��\ܖ��i���޻��+!�?�b�ʰ�����
�e�T��0������P7U�PԀXT�����N�q�{�a��EipL������)��m�̎�����	��0��'��PN�}�e�nxBk���29���Ė������o�SH�++������N��E��aEĦW�Z-�sS_N4\,)��}��=J&��U�:f�RGE����q &��.�q��bZZ>�5�v���Y�!Q��V�t����M耢õ�� ;9�����E4�
�blY�~a����5Y��<VO��[�c۴!_���,��!�Mf]�-	<���7lM�T�O�67 �RU��)CrT�7{�1R�#r��B *�����d�:��Ӓx�rv��A��x�n�����ܱ)�	'�V�$��*p�2B﵋;w[(�
�� h�g�d��篘��#���
~�X�Qp:����i�%N\n������]yꂥ�+���f��<!g	?��_\�*�_��8�~4Q��4#9���Ju橇-����>h�PI�Z�Xi��M/��"Z�]�0a��Z)WU�n^�?��|�k?�"����Ȍ8=������_��C�F"	��ڪ����~pLx�zu^Ҁ�ia��o��s�Y�,e�u��5_��FDc����h�2d�����b����U����'$$��]��De�wi�A'��a	���,W�UGZ
]�� l�@q��[���H�6�j�]sEkUS��Y��*2,��a.W%�����}W�0=}��:*����P�EN����y]���r���an��K&��DG����zZ��uſ� 7V���+��k�q��a��&��l&��,rw�\�e�?��?e�-KDe�r	0v/�ey����ݩp&��+T��K
��	��>��<
��� Z/�����:t`^�!�c'v���+��a��Z�����a"���g�T�
A+���5�U��� 3�;���ȗ�]yz�+D`Հ�|��{�l�1J 7�����U-�hgH;60�\s=�ͫ�o�Ǝ7X�39�},M+��P������E������ڛ�6����K�a��J��+����]��a#�/�ve�@�X�R�%�v�����K�L���^�I�����f"f�?��Z�1�M��sHc�>X��w~7� �������Y^�,]�:���0$�ɋk�K���<셦U��U���r������k�ʉU�O�ʕ��y�tT���F��O��}s�ln���駖�}����Y�n����\a���L��7��\��(��������xC"�ߜ����	��2ߚ.f����S_֍�s\<����\|�� ��s��(	l���8u=�No��wb����T����D�Vk�[P�sMm���9��v&�� r�}��N���H��%_Q^��x�H��$�r�|� |�j���4 7���'��P�ng�e�<0�m��;�$л _+J��t�=z{G�r%�W}�h�5=�~�v�:�Q0�t���چ�2>��|	y��'�ז� �xd<1��^Gf��㺟zT��ps΋���4�]�[�F�$/�t��Yk�Yn2zp�������ad��/�n�~���S�NKƬ�zz#7��d���
�O��1��b��,ru�H�	�����Lb@��-�8fZwK��Z����7����䥝�F/�cW�%i�ZP9�O���'��dV<2�v`ș�e�a�@hC�qX�U*+�Ž�� T�U�����=����fM[m�G����r�:w,{r�yM8�N&>5E �$�ڡ�Tף������0��mVQ��:�@J�af��碑��<]��c��S�I�zCe�W�^��^bl��E�*-n��66���0�w>�iS�����n�O�2�l�ܬ�����jQ�f��3�T�i�A�cD|�,��AWx#���t#��r`�I�b�w[`4�;��J��������KG�(&6Z���f�c８i�K�#Lؕ
~$ ��i�wa��ûK? ˑ.h��5r�T�# �h�nF�s�2\EUG]_�ү��������^a::�U֛G�v��;�#b-�ӑl�n1q.�ހ�]°1�۝=�Ym|�J���B��!���A�$ک�~������ݾ6��K{4Ӥv���4\nE��9��1���-}JV�!�H���0�b>=v3u"�[�DU9��G����߭�k:�^�G���e�
�U~��0�b~Zn�?}-����:.�32�,i�	�F����������+�-��� 3�m�e�R�>+A~�'IL�X 4OL��!Y������/%��]���3+b����TS����&S4G�]ec��E�$�6Ǭ`�<��6l�+����Y�ܺ���u�D=>��3��G@�����\�� ntc���9����K!D+lp{�M.�Bd�ڕT��]��CƼ��e�x�������4�n��PZ��*�JZ(�T�X��U��LF���[Qn��noo����a��Ҍ�әO\~7������\:w���~$�9-�)n���b.2A�U��i�6����~\x�dJX|��h�����O��r�xC�p�m�`4�g����;W0�G�֮2����}}��㉭�� ݅#7�  ����$�;YR�y��ҫ���Q5��oH�C����R�z�J� ��"A��5�o
�9�� �kk�@'ehఠMh��������=�@�����eU�~}�۪�h��z�y�X��G��U5뷭O@����~�����,�c��s��k��/����
��/�c�i(��
pPWR����zMO�:] iOw,�ۣ!�ܱ�.K���k�A�ځg9�J4ɋ�*�?C�	��c�g��:��6��(XE&���8l~@�!gF� c.S�o�_>|BU3w�w��k�9�(ɡ��*X\�)5�� 6��ѩ�#JJJ05����>}�"��.���0KW;��-�Gm,� S�-{�Hi��~��ӑ� �h��*J��|��,+��+�B��z��q�?�g7n\·0L�?5����-��=�p�}v�m%��7����~u:Z��J,��)�w���eAN�-�x���[�+DFGGZ���埍�һ8����n�{�}����t��S����|�=@�i����K�v�4������-�k�h�.���%�ɽ�}G]��J3��4 �-�g��5!f����v/�i�@> 7�E����e�vs��!6�?���s?x�,�W�}(D]�d|��@���nȭ�ʹ��\I�($LR�z�3��
�q��D欿��23�J�`���ڡ?%<��H�d��6�i� �r�*a��o�*.U@j�� R S�(���%�FC��a��Csꦰ�G���4fOXp��xl�~�K���3�K\��<� �Y�ʖ,�:�ƶ%����u%?�z�Ԏ�]'�@�P�!}]3)��ߩH�s�kcAY���<��	L$f:qqu
��F��3��_K��-$;�3�"w�����~oP����^� y6��ϲ|>)5�}����nʚ@�(���+��pF�D-#�]Ẋa��,r"�"Y,��I�0G�����%���ՃmHy�n)�i�G�l;@6�-�(��(�n����X���#n<O<&%U�=�RX0��ǄΠ��2 gU��&畠h�u{ �˖����2���Jl�Y��̘L=tK�	���C���w�6�&w������U!�z�_�??x?v�Q�>*L±�6�X�	�yuE�;%1����G��&6h.m�����#���P��uF��lm���h-�=Wr��dZ�l��(��HN�)��9	-WçW�P+��Z�n'+�8�)�:u�Ss-�S�G�J\�w�7�K��nў��s%�Œ�����Ɍ��~�7n21�^_��3�N|��炃��e�Lԝ��hz'd1?�gØ����G��'�>;�([�&6���]_ǔl���$���םb)#���$�~iYvy'�����0mĲ^��K�(u��������Hi���)�T ӇP�X3�X�^��'w5��G�y��r��e|��qg�0j�(w9Y�+�0���c���z�U9�{�E!V!Й�Y,�`w��j����O:4��1\e�� ���9�&[��4�vxt��)#X��;N���0a��
�� ��]s	)|����c�
�#ŀ����9j7���R\\tH�@���"Wҹf�|w�0 ��l���+��v]v��V�Q.al�W�<]g��G�ɇ��7�� hRqw(�$��� ���$'7䩲n��s360��H�?�u���k�30�aW�x$�~C-�8bwʽ�(�a�ފ�1���7�h@V�,�0Z���PpGs��,��Z)22(B]fg|ް2�`���V���ќ��C��t��h���Xb��d�p�� A~���_]�줫��b���`�@g���4l7�of���rD�h;�#���������Hӏ��zu�aY���P���~0;]d����&�~�):��{tA�8��^��oa}Nwd6��,{�s̮
�Ж96>k`{D����S�w�'W�|2�+���Pa]t0�)��ˢh�+3�[@�-���J�@�-(�i\܇�R��5��[P5{b�vLb�dx�����3������6/��֧Y~Ű���o��<�ϸ�s���?�6�����d;�Z�V>l��;��2 �h�Q_�mbF�@y�;�o/	�n/��"��|w���1��N�+� �GN`���9�?�G��uc�N�2��S��W(���`َ���`�q���{٥Y$�I��< ����۳,�6�|q��Z9.�B�y���/ѻ�}��r����,���ᝉ�<� ���aN�oO�E�=N=- 5�)'�ey���<K�(��r⇛=LX�{����^�l���j�V�Wy��Z ���N��^|¼t��Z�tD#ٽ���������En��f!%�O]��$c��H�@�D��I�_t�f��ᆽ�$\Bá��ʀ�It]s��ܼ�z����A�s���	,�sP[z�H�Q�m�g��}u���$�@9a�OxZBv�މ�p�����bBa��J%iE�(i���F�8al���a
1����%�zxw,�7ғ�N�!�F��5u����O,����h�^5��r,'��1�\>/��+S�3�mS揞��"B�#��2�-��י*�,};/��M�h&,ՕW
T�W�f��+,i��X|��Ny�PAy����\Ш�MY���|���X~khl����o.4H�mF'���=�u��Z1���πK�V!LeiX؈yE��!F���p�8�mX���[�W%��Gq:��m�)R�m%tB��>��W�ͻ�,����n�z��%��U�e��SɌ�а�쇥M�h�x�v"ʶ���ڤp��Ao�9??lb���,�|&;�#ް�J|�i=�}�i��	�7?G?Բ)9����X�3WU���1��q5g�d��� &���?t�G��?�֫W
vG�r�DM���<)���|3�, �%�46d*�_-
�p��J��2=�b�} #�� ��2�YGC���y�/N�0Gh^�@��<�4+�<�7�]O����Ϗ��mJ=�WWXCM��1W����fF/$T�"�����S��7x��bZ0��m��%jjN������+K�r��X��Ht�&�,d ��9����g���q<1ȇ�X��pȋ�����J���_>�(Y1���?>C�:M�7����jqiIM��y�������ӧM`�Y*Mt� ��a[ꡚ���]���u��G�>�"���ϐ�RRRX����t�40��5���15eX��KSSS|=�N��i"������n�;3S��8y`ķ���أ�� ���5�4��n5ӹ���_�����ٳg��l�:2������S6=����Z�za��vz|DD|*�:����S�:����K.�@�� ���[�>�������J��ƍPu�:������:������?I�.ZR�`�UG��.�R���~�q/�g�Mx�`N�L ����y�u@ ��@RV?���l�׬��g�bb�	f�v��E�K\э������3VL�:��~����b�VC������!�İ�Ț�z`�4�����z�,��4�!|~�:�����K�����6�x9c�����bN���~:FM�+��kk�D`����[�/2K����M����©{䔎ԅ'�G�q��jWhd��Em��`]C֧i���f�����!XX%�*T]P��ǿ�t�����w��8�^.�Y0r��/|�;<b�o1ٍ��j{����B����sB���j�g�ɮ��n��p
/���t��yPHy��=�ɯ�Ŝ�:}����o�pW�g���l����X��eo �&�����K&I-�ŕ۞[8Z3Ʈ�P��)ϧd$E�!�2!d�0|����M�����1�1?N�h�:u�c��!Ë4�={��'��}j����w�+����ZX<S�k����Hj4�����9�_��O��������8���{<]�H��p1gVhu���M�gB��F��=�-��M	�N���>�4b8�������/�.���7�f��_�`aN�U��i�Z�c5z=�t��!�u�bX�g)�\/�b]���l�\/�#��
�u�2��.?�=@d��u�<�J�����~(o	�]����!jM+�B\wLmR���#���Ko�_b���vcR2��^��P��?����-����]�8�(��%��F�b��'�&�a��ȔY_��Q�QT����qXѷ2���#[j��+�m�U�aK��Iݤ�@XG+�2D�?����"�ǔ6y�P�;>�>�e�q�ћs�#������z��Ϊ
�˘�-��+K����76�0�������5p���Oh)�~����S�AE9""RN|4Y�#����!�Va�LPm#ɍ&���ݱ��!�,�r�x��Ҫ�6�������~v��};6��d`R"�}b�\6��*�a\��O�������\;�����9u=�؃[n;�k�n��_�;849��V�����7�/��]o��γ h��G�cG�c��R�����5�2VK
T���;xMh�ph/q�����xF�,�ak������d�#FЫ5�����Ԟ͘c���qbw�DzZ5�v��k<�������.���\��9&�&@���ϾS�,j��g(�/��q��L`0/QO�&񣍻��S�(Et0(+����ȣ�q&z����~�`;h��̖*+�F����|�掤F�: }��i�x�Ğf��gi�Z9Br�u^S�{~K^�d���":״�-�ՖM�=/z��=����Sox�f�;ƙ��KD�|�&�
���s%f�f�a��h�҉�&_���nrm��?Oh����kg��8E��a���JgS����$���7�5��|�n�ۃF����tN��ċ����Y�p�~�\����1m̔(3��L6*�����_m�E(q�y�6�OT��lc5}\ kM�Sw�J�o��I4�o�#E�� w���w�E֎��w��d� �Eҏ�9�s�c��$F[�G�'�z��ŠE�g��3��9����X��ar\W(�I9���)�/��329���<�5E(FoL��'����Rp����b�nSw��a���Ԛ*q��w���/(,Q  �'��ߵ.�jK�(#.gj���:Sv��N�!{]q0J��w�����u��c���q{�`�e���N��byJ�\(;u��c(W����qE����9:��ތib�J��\�|՟9$tt����|驒��ѥK���ۨ`]�8�S�8�;[�;�g�є��:�(�,����B��T�nl���ұ�}�ٮ�{��J=f������/#��/C�����~c����(G�׽QCw�/�Q�in�Xɨ��h�i��!3��1�G����H��SR�#ם��z��&���&Oc3-?��)����q\�͗�h,��N׀2�4���B�L�����/�Ϫj��C�0���/cK��������\Y*�x��K��HG?>��zzh����ūV�P�b�y���[V��bg�4T	���: "���a��.�J�Z�a9$Rz���.#��<��>=�s�Z�n�i(��/,t��G�����w��r6���OX���f�ע;r$�9B۳x��`3YqԸ�Ui �)���?(;�/���62�.�G�������	Fꚛ��4�L�L�H���yN^�+V���og�d�k =$�h��z���M]U���T,(�&��O�?s!�<�>g��tȚ"2�o��'.�U�aaCL~��[߻�����0�6�q%jʔc}��≧���L
���G �QҜf)��ŷ�Jo�lԌ��i���.:DS�8�җ��\8,,���@'�:܉i��.��$��ѧ�����!*F�Ŗy�j��k�̈��TV�޳���c��+���ruԲ�s�<@1K��J&��>omz��R/����O^]gp[�>�<���e�����ܡ�8^j�ZN�y�xn��c���Ԡg��H�����X��~�qK�I��:U�w,�$,��'m͹����n~�'���\��7��Ὼ x��ɾmk%�S�y?�J�wN�[�z�MZo�;B����K��zA��狠�r���H�ִL����:c�B�7��Ew���*��S�^�wiI-}��HE������[.��x�_�?��j� x�_vM���Ϗ2�c���W�ڛ� p��Rc��������:!yU��Ax���K�Q�����yhP�jj������K`a*�{���
�t)ʺ�����\&��/��u�gqG9�S~� ��1	#�>�;�^����#.�L�F޷�L6�Չ����i`����.��@��6?�!�X1��P��5�{%t#3+3�N�gd��)����墜"�R
CB�W���3l����P�Ӳ��xmyQ~J�-�BǮO�<��s�y9���MK���k��������l���f~��ɇ|/�����˾��\k�1���'�w9�Ȥi)�u�h��%����r[:�G�c��aRt%�6��w��$�ܓ���q4E��5D.��*�8h[޼�� 4 h����ђLʋ������.�+�����[$��&og�PN)ޗ9lq��3��f�a���m���j�k���.!R<�`��g�M��ɼ��L*ng�-_LCX�שc�npL���{/���rc�km���zU����.����M��Dr��IO���:c�,�z8��}�c%[��m}ֵ䏶?��{p����+e<􃳂m�e���V�S'�-�PZ�3�%p���N��y��ژD�"s�ƹ ah���%�z3�~���X��t<J��gU�a������g��O)�ѫ��]�W��QuM8�l�����6���+n���zp3[��25�D�u�V���� <�i.q�m����Tf
h�d�z&�q�������Z�	��M�7��n��ϋF>��'8��[�����~�x�Xau ��/<34���J\nߊ��;����J�7w��ᴿ�à�u�GP���^�2�u�Q9Yّ����7 ���R�gMUy6���lL��Iq� ���Of~d#Sq,��=B��z��aw޼�'4����ڡ09�#�e�2w��u.d�v:�F��Ε.����Vy��0�Á۸{㍯��3d��5�%1��gv*ѳd�B�OA�mN��ǡy�:�Nɽ�%��.�Ƃ��O�˼P����Չ'�_[b&Q�6g�w���m2|yt��d;Y�1���ҁ+��ʠ ��g_��y�}��Qx�p�������9���qV[fɢP����(ܞSRw�W"�9�eE�Po���9'9����V��k`Z�����h��x����A˱}�����D���a�|��I\�����Q���6�>�>]]1|�uN
�k	����ѿ����  *t�!�L�ֽA)��Z�X���uPl�ס����!WV_HI`C���_�$N���������U���݉�4��Gh	ҷj	߇KЀ�p[eX��ߎc�׍�K�Nm�%,��TjBN���� Uee'x_��#?���'�X�Nf����n��>���+6�S�ί� �Ѓ�SlxJ ����-�����?��X��u��B�Dq�R����ӚQ�,��[$���,�,տ'�m (l�v�A�Ӣg���kJm�\�D��d��3�C��f�[�?���a���Z��W��H+�j��7�����f�����$�+�+���s��8��z�)���������9�';l�Q ^���%��4Yi�PY՛�� ǹ,x�;�<].*��1�𳔝��Ű���T�=��F�����̹��W~��u1L��L��J{�8�%9��p	Զ� �T�Ib�,��i�K���.�,���}f#� ��j�f5���ؘ������	�4�Yei2�=���N�_��[V�(Z���b諙Ug7��J��lE2dh�[̈Ғ:uF���	Alt#ot���9�Pq���M�3c��b�G&4~W~�3?D��P7�1?����M���ǯ����9Z�t�J�S�9ӌ�]��' ����� NFZ�!�Â_K�P��:MϨ�2����0Q�XRX�,*,Ļ�ϫv�CK2a�����.����Ȩ:���	��[�~Z�~���Ӵ)uНB��ܼw'W;V�l���N���2�S������T�{y]Y(]���2�r��7{�}�(�3�TK&������ �$ZZFfl�2�O�0[>ۯ�w����FZ��ӋL���4:�����Wz ���U���hr��B�ׅ��N�'+k���0;5�¨��!�e�_�0�&�c�@Э]�_-4�F)~��@��bJū�U��|�L1|��%o��rA��ae�H��k}��gs�9��K�E����{k+��oNC���L�tD �%����8]�:�?���mr��V=hes���%H�N�ܜP�x�`�J-�O :��44}C�7��
Z�f�Ų�H3��fծֽ���HyI[/�ٲ��t޸���>0O{|�6AKYd(���K�@5��j�ң%{�O���](�6.LC�,��z`��R�U�Bsfa[�Q��EeMk�iO���!�$����7����|�A�z��z��ͫ�\��-\�����:Lf�8l�����H.�}ć4480�B�e5�f�ori�z�TA7��ɾ/�f�Z"���j���U�5q�C�P̡o#�u	(e'��ߣM|��m/ޯ$���S�ݠNܞ��Po�r�����TDc���ω\���V2��i����[K��v60�|�M���e<��g�6��գ3n�	]9ȋ�B�譧B���4>Ḋڀ�;Hç>��V�Z<�p{2�xptxГ�`k㫢J��~O��Zd�X�l���GpH�~��6T��
F=_HP�q�ؘ=;#|�Ժ�� X��
�KͶ���H�"��d/S̅L6��¯���Um˚��BS�n9�`���Y��RtPl����yM(�x_"����� ��ǤQ޾���RJ�	�8�zLo������'��&�Ͽ�Okj�p1.���������!���$m�P��kQk�!p�rhY�/���做�Y�E�lV364�3�%�$RM��]9��>���Wl�ayh[L�D|���b@����/#�z^F��.5�D�E�@�^LwC<����~	Ջo�STu����O_�Z�y\��ҭ ����r�d�TPAiOtQa�d,�u����ox8��҅J<;�7���	��BmG7rB�>q�3x'�#?��VW��uS�}S�7�q}�"^�o�����h�j*K͋�7��N>����`��jB:r*�Iގ�t�Xޒ�ox=���W�dT��/E4Y��JK�g����cCIiE�V0V��'`��z٣t� �;Y=��E�{���%326�j��w�&����:A��s�c��B�v.�`/�~.������>3ut��(آ^-�����"{5���O�k�߈ S�SGcq�P�����Õ��-�m{⃱� O,r��}f0/0��a� ۈ�^edn��+/JA���)�q��c=�8v�N��DXSS�DE	�������_)v��z�mo�����4��('�iQ��kz��� ��C���s�LE���r���br0�JuC��\{@���~;S�<����#kkkP��I+Q��vg�&�,���8�U���^Z9ʀ��]<"%��sGz�y�)�p���L�37�㔇j�#��j�"� `f�s��~Nr�}�(�����9υ��ܞA��ɩ� ;�e�P
m��,LQ.�����L���e�k�`=��\��cL�`�>��/O�G�_�:,4�߲��U�A�w�{�J�Nqhct8|϶��e�����긕�W������$.�fI����T77ٌ�=[^���&2d���w7� �,�	T�C@5�w1�:��G73�p����6�<i�w��׵%�6{Sw�T��8RN��Y�Zd��w�i��$������_x�z��t�LZ��B�8�cSSM����4�TJ����R�΂Y�/�� ˮt�5������lU VJI� 3�?�Ҹ`�z�L�v�U1�X�Y.[*���:���Ϊ]=$;z��A(�Qd���>j��V�M\+B�!�q��3��'�����ka̺�<��.�`K��Xg��q���������in��kd6ʹ����"����v���o_��Ӭ�"6e�3w�+綒��$W�0e�bN�;tNh�n
j\�1����oؐ��PR��h���e:5��Ú+�БԞ������ϸ�����A����
4�� ��D~5�>����!`�w�ʕPVڷ�,���L�\��m�m�RK���ճ��fz}][f�\@�JqI!�.(~�$A���)�� �fS��SQ�f-�Ƽ B��bk74���}m���Fn���7۩�4�u�@�V��Ե׬��6�~�*���_�犏Ss�?�,_e
4i�Y��+�2��@-3%~�-l$T},��l8�r��I�^�=BU�:C�u��Smm.�w�瑱�/e��7yҿ�I\�t_�/LZ��p W�,�l�Q{�)�EP�N���x�%�c�����oF�n�[�%/��y+�'�,��p���(3N�l�_?:!{4vښ���i����kB�7�� ��̰�*#�n����@ܺ�0����o�O��bߊ���WĈ-�]�5M�#�6�Z��ݦ��#��'-�Պ�Vz�󣏫��L�\@��Jn�ϡ�Tt�F�wW���W�6 �_y} �[����B�x��� /�wpN}��f�(O@��5��s[ӯ�B��&���}xX�$���T�4#c����Ẽ'(���&0�,F�����1�@l��Q�Ԇ��`9)�Q�Y���57߯珤�Ov�>��Vj��K^��Zl��oV�&�)\�`���"l��ky�ܜ�$C�Ceޙ�^O�Ϯ �.\�).�t�=n' �F��	���s#
P�\s���M�#,6�� �O)·��ty�[���-%E��Iӗ=�����Z��g>��Â�^��8���r=ӆ�>B���,D�����3e�����.��8�V2��d�#s�S�1���u��ΰ�C͋����;�aCc�T� �!��
�M�=$��S��������R�ƋC��W�f���ke]��}��S��yn��5㉌��?%�&�(+���R^"z E������6��3�2�7�
�"����I���|ҕ��8��7�Ys�:s����:1�/���7-<gvO�v�� YD,�t�����W젉�/" �����a[e 5R�]�� ?��
��D���
k-�WG哃)�!_?ݣM.`~�=�e�<L+�Z�9��({�Uy�T/sOÌ�N�T��4���eA�(��x�FX����I�<��qr���/��y�`�j����xpa�A��۫�qX�"JK9:Q�+bذ���.3� ��4�E=��V���v��F�z�K�>��#�0�R�bt|���,!Ҭ+��7�1���.	�S�������C�]��g������FN�-_�1RpU��1��o�k��zg�y6ۇ�ֵ+�c��[���Y��0��rD�xT�Z~�67��A�D(�'�>?�t^}��l�����<����E&�XJ����I{�/#�֣jDr�,ذ׫>\���p:����H�J��-���7�� ����3IM��(����`�̬�J���r���{,��z��xp�����ΞQ9�)�WW�yi��Ƈgp����0��\�G�gb�ڵ�;���W��cۈx5c�~�v�}�lP�������qR�y�w��u������R'�:!�g���QVy�/�~ݬ8|��L]
~ɡ"�,��]����S�K�[�t��\��=�nm��3�F*�i�
\�{��j�A~�F�4D}�����:`�y���1�JA���=��7n��#2|�>��sk�?��N���DX��A>|u����;�F牡e�	wY2_ `���A1Yӟ3�G�/���'N	
�����k��x�MCꔕ��> �>}?q3
��~���h���zy]�d�~������G"�Jg�`b0������--,��;뤾�e8�C~*N<���addds�e�h�_F�g���z��?1�Dm:�  _ 8��ܡ��{��J�R�G&��a��*�=�i�!�^�M�%���3�8�,T���Ւ"�s�<�}qcC[ꬕfc
��J�&��R�G�Ŀn �:CX0�y���l��c߯�K��X�X.�&��"O#2��G�%?��Ӗ�����57O��~�|T���F��7�G�Ё��%�~{^܀����ڨ<���-0kXJ�O5�M��u\m�۬���|%��b���:9d/P��X�p�� k�2� 8?X�M��3��L����&�ik��R�����Wןؓ��<N�3�B7�ϯ��x���<d�Թ \uY
t*��<�"�-�-a/StY��n|Xn�G�d�����+�{}}�7A�y5�x�Y]�|�,m	��>Z���/x�%�䤻O�s	�ܳ��ǍٱXR��V�y���U�����P�A鼦���5�����Q,oN��W����_�<���<�������@���i����g���Wn]��_:OU{�o����ЫH����
�*�.\�iiQR��n��6 � �ݡHw�t�t�Hwljҹ�t����Ͻ��9�Q���ff�����Y3�1<,?�L���b��Y����8_		���y����|�i��V	c�n=������2�$��ݹ���{�;�0�J���u�� G��[�������o�!@ۯX�gm�H%�(>�_=�!�?M ��-a�k��⇴��Q��������,�p��N��������f>ϓ�4E"Z�4Xy��¯�ޞ(������N�{���W�O��7��3��<z��G�ׁ�M%������\�$���[@*��惺�L~&h��V���~��dɀ���ٙ���������z�iN�e |c�q~<���6]gg���ݹ��0k��d�W�v���ᰝu?P���,/��:dI�~��_�`���6��i�����ʊ�u��E����"�ճ1"�y��G%M�'����ɘ�2oY���7�ܞ�9
1��������PP��h����4I-h?��w��ɜ�W��QiW7D�/8������~�T��H��㜳r��ؓi��F��`���k}0�Z5���r.	���, �B5@Ā���1��m<���	F�L��3�j'�������68O��
�"��{�o�W��i�J�TT:���2�ʘ���223�s��D�� �������G��̬��JDXXUUug��墽4;l#eEH��{${
i*��4�Qc�j��2(�}���jf�'�?jns6�`�.o�Eۗ�3ȫ������V�����{�Ez��1�����cBl&�CF4a�� =�,	ͮ(\��e���YG��͡�.�0G��ݭ���r�� �:��]5����o���gb+�;��L���7A�&ݹ��ʿW!}�j�x	2�;:aҐ"��7��'���Wu���T;�-�ȽO�_	�lL%�a,��FW*4#O5�v���le��f3�#`���~W��.�����s���?t�V	��]�`LŻ�+��R� m���O�l�%"X��؛��¦�; ՟�4�p�.�tv�F�p����)�K��W�Ky�c�k���I�������x�bzh�5�g� ~��m����`�?�E~�а�^�\��ՑV|go�l�>A5�<��#�c��i6<��n$��� ���0�mI�f'�=RO> j�;0.#�褙�G�ytAr�-L�]7��,��[C��0}�A�21,��׋̃�R[uͼ,�O�D��9�6�@��o��+}�H��x�({ܜ��U�f1|�W� s��$A����o�Bery�~��(c�*�a&�ru�0H�8��/�;�|Z�G m��<���Gz�,<%�����/*�'���
l.���L���^���̼+w���w��o���?]�Z'��^�9�=��[��ͷ����h?��~��C����H���xϳ���쌘�g���� �H����B��~�ׄ���7�f�7�$��͝�������5#��^zw��D�7����J2���A��b
�]g�����n�ܯB�bJNV��[��{]֤o9�F�{��Z!�"MMb�d�*�KR�˴=5��OB;k��8z�����[�]����t:�o;�%>��σJͅ���-f�����ۑ���̃MT��|�:�D�#P)�����,�3p����������`��	��2��^������v�9/�:�O�6�v�c�mS�|��w'Ap�ٻ[���f��1������7�RbC4D��5u�Y��~Dϙ�����A�����yʲb�q}
�? Odf���Zq3�>]���݅���{-T�
/=��x���xWo��>�	|�f�Ҩ�9���J�����0:psi_y?����e]�5U����%��]򖋇��ޅ^��e;U�k����:�� ni1Th?������I	
�Z�0�B��d�X�Qx�W�<�:u"��zJ<0�f^�k)nu	"�r���Ei,���_�&A��B�l&p��)���'��/�^����:���.��e�j:���ϳ���vTm���,�:w�Dޕ���qy%�.�����m���D�:�2Y��ƅK���<oy���4�ʮ_�ԛ��HIU=r���ʌ'���Ϳ�����L��x�#�x�i7	�S���&�˖�?�I��C%���{��gG��B�DTlb>VE����?�ə�t��Y�<�����,��==�}��wwT�BF��h�?�S~~��8F���O?}Ԟ�3h�[�5���/3�o�O�Hۈuv�Uon�s�������B�(���Ud�'��Sl�#�E����J��C���P��?���{7rjZ���\o�Ѥ����lh`k�,6a��"�c�k��h���&�o�����]U�W!6Dō��\}\s]�.E� �p�g��x���bn`��S�;��_������!?�Z+y����pv��t�<���٫B�\�+��Qׅ����D�;IU�MV�WOX�m�;��?w>���Ru�0�����,*�;2��~��ŦB�8Ϡ^���I�>γ{{ԣ��9��a=`8U^�d����������6[?p�X�f�dQ��%PeG>E���{2�z亢v�y徲�����j?[��4�y�A��h[Θ,+͈c����ԏ�Wl�.�������X�)d��K���a?��Ro5�"��A\��?j���\\HLn���l~ߧ�Y]����w���射شVV�%e��_W��_���Y�okwTR���=O��־ۼ���������>����Ɣ��ۦ�O�P�$��Z��j�\~NxH�6c�v��B?�W��@�!����yxe�����i��?��b�di&������p��4�q.�)��^��ﬠsAye���-�o������Ud޵�Zہ���	��)��*&4��H����`�eF$þr5{p~wY~�-��+�M�.����r�?	��������\�s[BR������؟.�P^�|�3W���� �E�}��r�����~+�����*'���ҒO��m_�?��N�nԦ�sA�c֦��W@BJ���c�7�t]cs�VI�w���C�Gū�24��U�H%��>~^&���u��,���}�(���\�������Ib��# �-�7��c�z���+�|�Pez��J��H��������� ^�F������?���
�s+���}ί>㏁7�G���J��d���D�g�&*�J�9Ѣ8��c�t=��xK���3:`�&0̴�������L:�_��r�*�.���nT�<�!���n�s��1`Se�����J�SK�R4�?z�"�ǅI����b�<y�9g�`Ҭ���&� x�E,fc��\���ޤ'���f��B&�h$�ҵP����4�#�bY�#�9���&w#FYJF<�cLLL�vI��m��K�=���#\�s�[;��ô[M12��\�����E�.�f�Sֿ@���m'f|Gܜ�c�Ȭ�lD�ᄛ�Iz�>w�C��SK��6��r2z�ޡl��VVRd!�\@���D!�����b�.�	�h6 qLG2D�9xzk�]�Mz���_�C f�ɕ�&�/�'���LMMov�Rds�R� vqs�RZ]��M�Zdx�d�>����`�|}����Q¿l �yJ.�0������ؑ�˃^m��=�^�ӥ&L�z�æ�f��u�d��bI�j�YcD�h�u|�X�{�|G�B�tt�<�3\7g����î�ꮭ��5�PPX(����o�GB�Nj����H�߰�Q�g
��;@�,Z�hB�fL��b�Re"��g��x�%\�;��!�H��{{t]g?�����+�~Um�T2go[�d6V�@o� ��d���9B,�y��i��t67�����'"N~��������>��+�ćJ}W�M�u�D庛<�����h;�|�A?~)��ߘ��Q��:���2���<�ӷ$��GTt��c�\7�)��$�R1(�@�P��ED|�:ْr��D�M�*|32(��`M��̃�&$*{�A����O���_���#n�����`d:�v�7_K\e� �����=�'��\Ć�Hg�Ҙ�?����qq���5�ۂ�L0�C�K�e�kͼ7C�v��q11��0v�c���?8O��0X�ЉY��f����O��c����i�B�I˳3A��4�ɵ��9?�+�Ǿ�\�͓&)l�<	qA�C��Z�l����j�z���{c ²���\}�WOǗ�k,�+�n��vg?�X�
 |Bge���_(�ԛs�{�er���Vh1XH[v	h����,@��\�$گث��QTV�F%wX�P��)&X����P�)1��Ff���iH߱s���R���O�U�&�YD�f>�)fc��l���b�����r��{H\�0!��ͨF���\Gui��r�����еD�@��B��U�R�lR���q��"v���Ւҟ!d�O�T�����C��^�r��{�6\E����M�.u 	��� ��zY9&��X��ǧB�g�����=�IIU֋�H���9�14k�-kxJ&I������q�͍b��x���a�>�����Pm�]����ށ��7�n����P��S��=/O,ۻ��Uڅ���U��ed�\�RVP���+���Vm�|n8mޙ&��ԑ�Q~R����M��B3��_f�<e�^{׮�a���_(d�DK"cM���Kz��}'��l�\�M���p)��j����tYf-9"_��L�z]��B��j�CǪ&�_u�9�q���y^By�,ߕ���VZ���$��g?��џrW�O��{zF��_�2�8��7��[�����5d��=չ��'��PJ�͞���.i�w����EMD��	���/��EE�;�g�i���'�*���}<]�j���� �͘&1������x���=}��i�+{�F�\��1��L:5p|��k�}JZ�>��}w��������k՘�r�9!K�w�4���C\�Z�l�/��3��m�!��+*¬hmm�K1�������\�?�X�/��Q��~	G���r!�'	$���`���?�v���WD1��g�o2����U�|F��@��Vo��S����TS��Dn� w>��T�!��ra��?J�V�,F��X�iS�;�6c`-��H4�H܂��q�`b-E��_��J�Ia?������K:df��L~_J�.v0��>�H�� 2��%9��Jv�Im~>1�z�z̻����N%9�l����b��T�������u��9�!@�7��Pe�c����-�{u�p��=z�z	�^�L�]�ۍQ�x}h�Q�~m�]yN��-&v<<<�J�'�'6�/_J�,x6 �	�"��������.��G�?�`�!�L�����#
V%P��:���N��]&`�74��7!Uh�ȄVue��ȣgc�'��̎��E�l��T�������.�K�d�<H��4�k�Ӊ���C����D�4mֆ��b�;�{�z$q�E���`FQG�W�P14���vܚ�?�ǟ��"�Am0_�.1�v�@���^J��e .2C侥~?���l����)��6Zi�����5Y�`(�6������Z��i{h����w�j���`y�����y���a: R+�ٗp먙o��;W�k��褆K�[F��5����������L����O����3�������rr�d��:1C�����9��b �I�6�oT#в���~����.�\����w�5T�-K�ģlR���P�ЩƂ�6ά_��$��[	3qfy��d?K?	�����-ֻ������gQ�1y�&˦c�i�e'Z����f��>%��i+#赢U�V��_�T��Ts�S^�0e
v����Rf� �6�o�/��L�������'azk��ܖ�<�"�	���O��1�[ؙ�p�6�K ՗��I�#� ����i��Ԩڭ�O��z�~�~D&�L���Xj]�m��5�VY,�W'c��P�;;LEk�8�G,.g*l�6����4hYA�gh��)�M��EԑkȜ�4�!6"i0���^��}�6����R�[U�1����,L �x��c|�J,�
�������edl,�|{y�A���M���X��~���:M'z�V���6�=�mwf)�,~)�]溧mUUr����=b����H@�CN�ό;j��	�gP��*Z?vu�� � S��5Cc�"���@R�U�����[10���X|�	�R �'
x5�`���D{p�~��������Jܻ� ���������XO[��C(Z�ﾁ�H��a�)Wy���Ӌ�!Zh���{ۛ7����wn����xnJ�Qұ����=��8��9��f6�x<y�W6W��k��D �6��6s�,%������2��_>_J|��:�@�	�(��I�V��}�K�"�z8��K�%[� ��Y+��:��;a��ԙ�<�
�3��9��:�[��kL����uvU��e����v��(��)���,�X6�8�maR��ׯ%��Z���>_��q=��4c)"�I�ߍ{J�Bh�ˏ*�&���աI��#�;���/�l)�4�f�q���a�`>�T���s�f�G���q:<2�X�x�V��#�f�X{:�v�/p�Vy���� �Pb���wJ��Z�� ���&X��������;�_t|҄�q�g��:���'[X��$i'�
N��~��:�N��i�'����bmO���)�ܬ+,j%U3;���Y��g7�6��ҭ�z�uבR�?�^}ͬ��خ��Tc��q��.��ָ�Z]_߾��Ml��S���� J�=����B�n���*������|&�N}$�-�=���ż5j3v�pzJd�++Y!�<�r/�ED8gyO�E8s���ԗ����]�eU�O��6�>w0.���ƭI{ �'�����w�[����~��M--�-<L`M��n�� ��<�C����a�(.;�9�jk�u�U����c�`�z�K|�iD茀�Ӎ��k��wu��I��S����0ԥd��i)�����q�$dt�o�0�b�;}��+'R�M���%@�.�YY��3ɹ;��DZ���j�$�4��n�H�y�<>H��ZN)�s��&���4@8;)m{�bp�YG_�X�#U#2T:��*'jfn`_�9TRaH�9O.=��S�虒jb,�ͤ�'�`�,��'~Y;�m a���o�<)�6���TΚ�[��5:��Җ�a7S�K"""�<�<���ɹ�_i<B���Om�.T�.(,Q��Z�@߷��>$��^Li�s%I-ʅ[eHs5���Fۨ:�y`�&�*q�jWp=�T>ބ(�۠��6A�)�i�a^�F,g���Y�������}좊��m|����\u'NQ��Z̖W#�nRn3��Z%�AQBBBq�е�~�ǣ*Sp販'j�lR:�3��j^-�'cl���ۥ-�t�)'��[�U�F9']�^E���oo�'����w�����
����(3���U�aw����<�X�&�N���z�r��=�0U�1I�u�2Y�r��$�;��aqf�W[(��L��s���U�ˮ�ު�X�Z�?є�/l�;��kV\b"��Xb�J�Q-T-��u���$���Sb5��U��V�Uz^��ݜ-�i�������ŏ�31RRR��%��Q�Ԋ8����g��jGEyE�����;Tŀ�Ȗ���t�ȿ������Ww����Xu�'�(�y<y�0������p˺�G��=�Ec �M�'�W%��+��s�Q&+'�Q���%r�j��m!��3,m�Y�j�;~��=�AI�(���"4�쏸[ �c0X�J���l	�0[7��kO-��ץ �����7�#�@t�w����ڴT�YN^�:�J�t\Ϥ��՟-L>��-����X�4U{c:gJ�_?���тMq�y1�����Ɖ��e����������O��6�blIy�v8	i~D�y�դ�|��ж�a��WCJg�׿
qU� ](�/:��}��o�¥oP��f�����bp�HP${����<����N3�1x��j�˛Ǌk��ܗ�g���fK���2>�� �Z(�M���3��n-����Č�j����`ʁ��|K�|[�j��P�n�Hu	��$ƺ&1�#�z<�xf(��#!���'y�S�w��5�#q}+��_p'8pG-��2�l̎UJ�?7��r�[�^���Ț�3��l�#
5)� ��jC%Ϛ�l:�}ijj:겞b�{���ǉA�[�s���RUEŌ��z)�� !n�+ϖ�MG�Sߟ#9F��J;D(����.��.LU
����q���6y�f(��UJ�7�܈QV����~�b�)�+��捰�Z���#�ْ�g��?Ύۺ|�W[�	uy:�=�~[��l�Y��\���ư�&)q�p����g�M� 8�������)��X{�ms��o�e0�8c�r�E�a�H�����(,mV�?�>�HH��3�Vh�͇֗@Zk����E��S/"q���T�����kW�қr��cAQ@�ޞ㧰�}nv ��J����!m������Db�[��|�<�|:4�L��������h��wn[�%*Ė���Փ:�uS �$�q|�?h9��]zh�N��S�G%�+C�%3�)����>?���	�+"=�J�.m�q��y�F�a�k��;�����^?�{��<d��4�x'���}5[�{++|��X�8���}n�#>I�k3�"�4��  "G�nwA����9Q��{�+O��pJ�u��(�2��6�L���o�u�N����y889m�,�g"deh�?�����z|=������Q�qY�0�6J��J$@�aY��߆� �f��)��:��X<)읨2R�R��`�#���§����̓�����vֹ7����<�s;�d�\�p�!�O���pR���tOC��� F*�\�)���fc\ϯ=�cL�*�eA=!�/E˫��v�T����B%*M����Õ��IpiG̿�p�jٸ/:}s~*D�8p��q6�f��/J��e�3K\G�R\�VH��C�^�=�^�pm(vt~p�ۮ�E�gK�X�\ߤ�ء2s��W/Z�,���s�4'K�I(>TC�6�0�������9�6�Q�&��-���{t��F��7�|�_�?����[�z�n������̃��);��n{��������xM���VC���/�����a���=�����Out���AH��u	0(x�H�PM�pN����us��[������"`׃��|��q'���k����q���^��P(��Lk75���ݫx~O����~��ϳ[��U%1�3�9n��2�T��W�+k��wq/}$Q��]�H���h�DN������fv��	D��vhppb�c��^zOOǂ�Ҥ�WS�h͔p'B�e�ޗ���N)��aX�>G��e����k'><�Kj�����|?�U������e�-E��_��5�,�
+h���zs�_�T���a����Y��R�X�|�W	��W�o%���Y��xH~�K��n6oS�r;qx�c��ٰ11}�1t��P��XHH�5s4��uL�\�,�T��O�t�i��]��\��5�e�^m��6��ko�G�A|��.��tx�{{�N��p�>¹����\�NxX9u8��C�m�=��O-�v�"�<�<Ŷ<E���*,�B
���)����sDJa @�9�,��~1���l��|��+Vmr3͖�� 9qr�4q��tg�Þ�^h���X�����d����M9��A.1H�E�eU�����������*�׈A�u�B�Q3�H$�-�p0e��s� _�{�zo�]�}������uXU�k���V���ƭ{�H��Fr��MEbF�Y�����[d:w$���)��PB�!ő�����+o��WUʬ B�Y����8PUYO��ky5Ng�?i��8�����~��f�����������2�L�6�fffX�v5110�ݙ�Twp�kgY񀛭�)eZ���#%*���h��h	)Y��=wݦ�򦩳8-M���a���-�\�s��-��Ln+�BU��m9yz�(�]B��m��ֱ[͛�\��Ȍ}~�N�z����d.��K?B��K��&E��͐ok�a�
�6#�[Kr3�@�{��/?����6A�ynu��<�0�f䃒��v��r�9�ŧ���UM�������z1���,mT�O��#s�J�4�����V˶�j6�ѕ@����q��7<�����f�K�2%C_��밪ss��1���)֒�At�\�>7��@�e0��C7	�U�Y&��Y*H�/9B���B�v�	�-f�4,�:v%V��{����0��8;p~��C�*�T�]�i��@���g�+[~f+������`&ʅN��j�F�*���*���M��[&�����͋IBǔ�p�-Ug"S������w������d�̰K<P�6���E���,}Z�)� ���H�=9�[�ti�(�S��iy�U!�W3s���^L�:Lou��u	�H�T�vT�R�n�9-
h��ʇ�����pFH��~CܢPx�b����)+ҙ�H�ѡ�Q��H���*u�zSXi'7� I2��������3Q�\�,
i��X$�Y�Y�� ��1�Y$˹��B���Hդv�ӂ��-�:"wSs�L<8WTS���&�b/�0'P��/���%i�p$��| o�صXC���@Nq�#�%��J���R|p���3m/��4���e���<F�ߺ~>��U�"m^��+�E9BWg�?�N
���Y�֠���ܕf��}D��G�-g��|iX��8�bL E6A��FN_�m�J�� �{��4?�+��.��s����`!djB91+[h�*|NthߚE��3�P��fK`�h�X����]@�ި�z�O
L��yT��[B�K��&����WU��y��s��������2[��(JNT�N�;�g�ș�A'�rgV�.���ͼN�L�vؔ�G�ݬ���j�k ����)��-X�f-E=a�8����R���]���������\S�@ߢ�#�����<A:���Z[�>�ZI�/�+�u�T���>�OZ���<�r�$����v����3�h��:�+{W�S���	�bS	���r ��I���Ղ��.��첕�k?�w�:�>;��������Iܑ<��S�s���4r8��������|���x1��F��}�Di��L�W���#L���R���4ΰrX%��@*�<Nq,Lv�`�"�7`��Y�_[ѫօ��]نϗ�TRGi��;��o6��H���Y�!r�fMq��k�
�{�U�`�fA�!F��)l.�kaS�":�y�v��m.�||�2���0���-s�� �/�Fߐ�o�-T)Y"�[6ww�y�i6��\&rX�R>I�}֌	��M�>�h�ۀq���d��%���N�˞��ރ����֪�q`R��+E�.	D��q�@F� $�A{�D���q������i��-t�ZU����PPF��E���!o+2)0�-r�R(j6-�ۗ�>n��|���D3��À3:@S�Bq�2\rU�!m�] :55��������EW���ЬL0�E|��v���?6e�*�{������
�9g����=z+�S2%�\t9P�!�:���ou8K&QG��&[*E��:k@*�m�R-�d�f���4�hyt�]����D�TP��z���"y3�b���8�&smmn2󠏾GT_y��A�o��*��@؜�:��x���*�U���:/\sϗR�Oh=�P���mSs��$�tD1��G&����ZY�����_%H�*�B��h)����rC�^[��Ig��ӓx/f�=�XC��$�$(�*r<�pU�����e�QF��KF��W��e���@�����> S�]$tJc��d?2�u��u���|�\$�z�~RP�}/�Vs���
DC�J'�^׋kT����8AN��40�h6�ظ�Q��Zߓ��.�O���<�e���]�	��(�s��@�n\��kaGg<l����f'�u���r�D���b-I���Rf�C�7p"y��n'�~������Q��0�C����a�e��{?�k�4�g��ە��hn:�
�����{��.JA�dp��
�==8O��!ycc�U�/�Ү��q ���2Q|��U��7#�z���R�bql*	w����)�ө�߭���w�������^��?OTY�Rw��;mr��@����}�/5('�V�m�XF� ��l_��{J(6�H�;���Aj ��rRx���>gAM3�0&@Q�!?�D}>& �����s8z�r\f�xc
i�������?� ���<����&���!z��~ޗ�(�!�����~ǂ(K��{	|�����z8#����?0��1���8�]) �;>��(����a�I�@p�w��ưK�<�7C��f�� ���B�L���R8��UؕMܼ�y��!=�W6ujh��[��O��O0܀DUP�
}
!�,�Vm�Q2H�6���-�h�J+H����i6�?"�v���I�_k�J;�ڮ;t�jf�1>2!�c2|��J�y��K��Ιf��Y��)2�ҶA�!��F�*/��s��+A˂��'M���l���~�@�w��<H���qg��v�����F���T�w�#��Nn�x62���gO�׵����BU��Ft�v�m�����H�N�7��'qh�9�Ĭ��������r8��ZQl�u��E���8���0b���|kf��:/5�lđ?�X�(hЙ+y������`���:��|�1�:���א�`0t
D�տd�ʨr�!�D@J�^x�+,h�1�\Dev�W�'2:r��A��ߖ���N��94:88��[��b�Aߣ��x��x�X��ƣE28lE��
����\�]�AF��?��9��.U%�q/��@B�_݉���1�2/`|6�Ȃ�����]az����|	�N���	�W���{zy�N~#�=Y
oO��6��F��Nғg�M[O?���k@Y���ЬC������������|��qV/��4�P��#��(HY']>,^�.�GwkW��yq�#_�Z�GZo�_�\1��%�>_^�Ϧbh�R`^����ܚü&"��?��x*<��c�����vi��#�/����0�LVb�Y1ɚ ]eNNu��K�l
 R����
�Ո�����G�b�/Qa[�z�z�k�]C
g�*k��t�qga��X|��v�]H��" +g�u�����ɱ^2B�s"s��/n�P��m�!��3M�'	�d1��{�q�}�%����P���ԭ{��9�y�d�\Xyꛢ����`0=5'(ٌ�� +0�o��^(�b�Ht-B�o�<R�"K\�L��h�ɀ�|�HM�/�tߪK&��!������i^7.s.�)9ŏ�Q}c��4߬w���F<y�VV�k��O�$��˥���f�D�� �	�
��vX�F����[ϰ�qCDʂ-�J�;/c�Y�c�fJh���Iqw����m$��
*���
F�Y�����b�$�h���&QÇ�N��N�界'�;lIj��0�ӗ$X/_�t9��C��0T� D0f����)���C�f�F�*�{?ࠟ�S[ac����ԯ��2^����Z<÷�-��7��(�~͏�fz��!�A�s�+������p�Q�H#ݟ��Ujk*�Bkm�ry~��U��a���IV	���ң`�ܽ����2a#��V�}� ��~s1���W<5�[��,�@�C%��J���n��#vm�g��8t[�&��n�m�H��H r=�OuG�!1E��Ub�+���1+�l�m�	dp.]�9�-◒�{�M3�i�	�ǻv@�_�w��?�K�5>s�~�<��"�F*Ho;S���<���G���Ur��=�V�N��dK9���O�OC?�0������:�>��<�R���2|5I�����l�����#ۤ��ފ&�˕��x�M�����[���X+"Ф`����Ԁ����}g���0�#�����
<�>��k�k�ʍa�zH�9��I�����OQ��2)��
&��i���3�	,��?�a�� k�Y�C��B��$���d�-pRʓ���.�E��3� ���O��� ��a2:�M�z7e��Ca,�Oo	���d�l�B0�����-��j�.���nT�>i8��VEt=���<���P�I}z�I�_��/.��N�.��u��x�ÔaLR��D=��-��W��pRӱ��e��(;��+��	�`[��� \XB�;����Q��+q�ۿ�q|՟y�W��͆d�&T{5�P"�[)W�;.����&��ʅ�RXFL_�ig�?��@H���[1o�#�������?8���`��GD5�[��ζ��v��6����X-Og^61* E���4)�7��:�]"��_���<�ev]gUJ����U�r@���p��+&H�IB�e����"�O�#��?v�P	���h�O�W#)t*�n���<x��B˕6�؁�>NiW���'w������v	�|�7���"R�~nxd����9���~���)Hh�"?Z�n*��*3�N�j(vb���ټ��t����{�.��F���i�`��HF��|-�b�.��J_6�Az�q�E���ZMڞ.#�Y�vD@��E�_2h�M���?dl��A�Lg{���C����B��-�h����>R8����r]���2/�+H_d{F�n$���@z���a5���0�������X}��̉�5�cp��m���ÿ�[��@��)ֶ�Y�)�G4�{mk
�ޛm�Dh,��Ij�

�JG}�/Q!>��o�����|����!�D4�2����v��|�8s�K�'�C@�O�E�i��@<� dQ1'v!x�$�RknZ�0NS�)�:=T	|͍�`b������}Ľ���ZzI���)Z�F��w�IrXd�]�Z�C��q���A,�cG<��!��{ܣ�*T.����%W	bͦԨ �et �B���r��-�j}�:��c]	높�@·F�o��Q"�d�����{�?��;(���1Tك<N's%G�g�1�#��l���ޣ��^��r���TY�h�/<���KI��2����L5ͷ�����@4,H;Ș�)��z�-Qh���zU�8Z�M�_=u�E��T~�faY1���V��uj�J�[qg��1�@�P�E��9�]Ƞ_|~G��*�v:�X-��Ǚ�P�R�����N�`�˗��,a�'	�\�6q1��|ɸ���C�R������"@�[���K�W������W�GL�f�Kq��O/�~ ��|��U���j��R�?�F�5?��0D&K>}��{g#��������#��@�� ~���LY����(�n�X�N��Ց��c>8�pHJ����dQ8[���e�b�~��0��qe��0f��y#}$��:r�}b�4H`28=<z�_?"�y�����t� s���ӓxq�p�+����&HiR��p�������c��ܛ����s/�l}�����f�Ar��ɼk=�Z��h�V�Ն
֦���0������.Yx�IN7������?�!�c�� ��A�)�-Wgs�\#@ �������������ݸ�@��NC��e ?���w�:�����"����"�sֻ�s�!ƙ����Z�x��<�{5%#�5Df�6�-6��ɾnW)m�޽/Ho=]x�
�҃
ec@$�f�xy<��, �g���p���8�W����<\C�p��L��#�qz�zJ�[�0�U�u�)c���뿃�u���7g���I�6�O Ja�?g*�A�& ܦ�����g�T�z/؄3KА�_F#~w�S�ҥ�����=;�_}��N~o�t1iyx4Q�&;b�|��i."H1V4������pʹ��P@��lQ��ޜ�gM�t޻z荧l���\��ԡ�I"݄U:����1���Ä�GHt�R�7�ܜ�9�n�`��˼�^FQ�kd!b��=K#KxR����?��<Щq��,��d��fPi?�7`�x?�%�NM%�b<:F�-���]F�8��T�yO9$���z��&���n�&�D��v���e}KO���F*��=�2��k4�(4M:��5��Dz��������Hi��.��`��<2b�������6	;����M��YI��r�z�p\���v���/:��nJ+�H�������HV�w"F���[cj�)p[��#*M>y�X�4�����%s�d�	]8b,��{��-��}}Nh�\��������Mƙp�����-���ň>�����·�Q�.��-��E�]cn�'8�"�#�ߧb߳��_Igcb�2��b�E�P/ffE�11ύ����������晩V�\*eæ8W@@0���q"����<ٰ2b�(�!U8� KƩN�Fy����bA�)��n|��ǰf�t�8�g���3�5���
����0�����m{-5T�Glrv�>�&��_��aVT�XH�h�b�Q��N�����Yܹ��b��c�A��@������3O��(T�
+������C�M.�(�2o�T�֎%\����#�k�݋cg�6��;�]�m��:�7�/b,A^��v�˘o��#�{~�lJ�hsN����!T�5[稳�wd^^X?�r�.��E s �rw&�cL�6��	�y��K�		y�����E;1�k��L�cL��gO������^��zQRZRQ�Tr�P�_�Qrtӗ�v�@��6n[�=1ꇒ���n�'�(4�� g�me�n�BMBއ��Ԏ�NB[_��_٤�_�jt��a9���{w��E^������k���-&��N}*�B�l�R��C���pG�_pc#	*���(ǐ�=d <�T+#�s��5Ӯ ���#2�!�������.$�}:N}﮶���~R&�ؗ�x��)�SQ����A\�,�W��z|&���l�4��5�� 2b�F�ܞ,����pOY���֖8c^ӧ�ɓѹdB��ʻ��1�7J��C[I�q|�֘�gc-\cI7��e�|�eY��R�`�����u�ch{|�*?��V�؍�<���E�骃��9�>�mys���F^�S`�=R�t�p.>@B���,�<ڃ�����9?$x�#��0{ٕ�?���ςB�4����LF֦��ѭ�TG�d��ۓ>����w���F�q3��kJ.�e$&v�N+͞���������١�f��Q23��l������D� �A�*(�Nif�o�o��eʣcl�HO&�o�zbI���H"''���j~�vp!���J���*_���W�x��ɓ�,Ջr�������Q��M$�;�Z��ʼ�"&vw�ƈdl�68������A����~ɬ_^�zZ�@�{�CO:(H�coe���.��ª(
(*�te���(�5t�(H7HRҡ(�� 1 ��H�P�yfpw����w}\�׺��<'���9�9Z>����ط'P�hO�{aV��"�ы8�},B��ٓ�B>{*]㊔C"YЪX &�-7"��T�y���Em��1p�N�㞜+~(F�*w##4yڕ� 鵲K&�����S�+ccoq��z_3�/w��<c�-�U���=HUQa��2t��� �א�S��/���o|�8j&G������2��>	{9�,??�P)1��N^&�?�8C��
=�l(iQ��������斍����VV�c%�{No��N��iky�<���� qs7k-*'�ɫf�A>�Q�[���'۠��-�»x8��&ڔ$S$a�\/���Ttx��ۃοǵL���-���*�lܙ���nuZ7�=�uzX��⣚��S���T��|�2j����fo�������-p4uߘw k�/�������E|��j0�s���'ߓ��y,V�6���\o��7���֛^�!7o�{�*_���kr�w쏫�A�G7w�����o~��vn޼��cF�Հ[C����W#�'�?�¶i/�@ޞ@��1P�2��ҧ��./���sY���[������J��?����9*�Nr�Tk	�f�)Jct�������'J �~D�,��g�/�c�f�L����.���s���BM1KΓ�:/p���x�)^� ^b{�ɠ��lT>$�pP�M{�y��Oѽ������ـ��o���$�� ��ވ�Å� lP�z8���&�Q3����H��*$�r�3�&6��5/9lO���Q���{�%tU�h�Y"C ���U�6�\M�����i�t���@V���߽�N�W��S{Mpy1
N��/�钒�v�גb�F���Y�_��_0��/��V��.��ʨ/��y����D���v���k�p;�X^Lm��X8R�����A[��-���TrJ;l����Fי��
��Ӓ	�+F�5��s�]��0Y߿��}�I>ȷ#�O��u�힄�¿X����	��~��M/C����M�ʇ5�ɍ��|�*�r��]�4%?_�E_��[2�p��3��v��89hk���Oá� ��ʶ��$^�E�*;G�8I����2 5{��y"V���a�Q�fn{fw��y%�������G��B�`�2LG/��������ך���e�Z�v����X�J�xO&]���FNשP�fJ��3�������%���qÌz�:,����[]M_�r�6��X��B��ĳ!�н(#��"�yV�d@2Y �񩎳ʥ΂g����&�&$ǭ�z���B�����M
�1�"�� _�e�k6������ߎ���z�^�7
�T�ۓ�o;p�x/a20y�v?3�_�l����͜���6^���{���@��f½>��"�?��ގ�(?��|�/����l�u��f�L$��b�ŵ���$����q���06e%�ld� �����������}�4[��N���S��ЫMg}�ɾW��n�]��/)�M!9�oL�f{�AE��l�z02�݁#���8�����O�H c+� ᑺ`m:B�\�e�F?� Mu�$�]�ɣ���T�9j�y�'3�2ǥZY"��i�k`S�
���� ��6Mx^{~N O�(cp�%r9�Y� �Uź�*:%[������ſ&���ń>������Իwn�^ݰF��CǱY�t;'�!s5�5���
�*��]�ܓl�/�#+���r|]'q<tJX�� ~��J�2��Ւ���|[�F�a�q@E�Β�wc�9���|�����@}Xν�s>Z��3�=)��k ���ƶ^�n0rr:}&��)�� �h��/�*0��?F�ɼ��z'Ɠ�F��nll�׽���E�6n��d;?G&�h��a�Ò��"��2�ۍ��(IsVJ�~�S���_e�*w�|Ww|�v����ER4=��҂��rE�~���ّ��]v�a�|��I�4^;��F����.�V�Xu_�̯�z��^��i�Ͱ�u�ō���J4 vjּ��]7�f�>\33H�ϊ�p�D�t��vh�43�Ȱ�@g>*��`u��L����뗁�Uq�	I��j��܁W���lͳe�,�(�2�0&��g�u�+g�� �~�|����&����A��0R�5��&_��\��JX.�*u)e�Y㦶k12�b�Ŕ����Hl�\֘8f�q�^7TY��@J9I[�k�hfd<[S�5��!]��`I���mTT����Iy��?���S�8*���9-3��!���X��^�f�1=
xr��oI��/{Uˤy�W��C�+�/������w����G�Ye6�2C�a�r�]yCQϷA��l'�$ϼT�Ҿ�\_T�닕X�S��հE��J$������ih�_��	��;��۷���o�{���d�UUq����6��wLw$���srN�O9]�h�>�6��c%�-��ځ�"��H&��&�9_0�crWt��Y)u���� ��2�ÏVL��,�hPX��Sl�W��̄���p���=C�7��_��1�nZVq���Ӱ�ͯ/��/����`0Y�V�.�`�j�d����Nb| �D��]0����@�\�;�I�����W��iғ�i&����u�/��G��:)�� \��Z���o<��d}WG��ܝ����Jy4N�����1A�/u%�7|��>��"���Ɵ�)p��prn���+�i\���X��w���rT�<x1�|��-���jW������9�;�gg����?��E�_�t�g!��D�f��|N������SM��&>�Q<����TmS��9��Y��ۣ=�1��R�,R�Jf(�A��C��bh@-���v'��{��n���:�M�H�0�s��'?��g4�mu�hi|�����F��{����v���n�l�	}����ۆ�2`҃���&�
C�Lb���6Dqs|=�_g�Ϫ,�wn�I+ʐ:��v��OM�o�UO��k2�&��s�?�{����d�J&�&�k��ܛh�禨N4��̎�Dr2p����mp�V�������B�t��&�wM���=1�I�E�8��כ�t[����� �<D�)c�Ppڙ>���0�� ,+8�]���/Ee�ѕ�(��H)�g!�9�e� �q� Ɏ��B�r}�ǅ��%����t��!Tj�z��BT����R	���O5b:~ֻ!��C�����;��^���:m~�K�\�3���-��Ϗ*����j.��I�X+(����8u�� ��r����dg:s�|ɛU=ޭik[��zQ��3 ����\��|cϪ�����Y��u�	aO�����BzgYIq�B�q�ݘ�T�~=��]xUM�\A��&�3�!���A��*��.6J�fS~�OU���&p?��?��`���6��J!��ԸV��k��+���ʻ庬�oT��٧�P��{C�+�c<���W[�����gP�-���/� ��FG�����2g%M�A���rKĞ�84;��0��~v��er��� �,����rMb 7��ȭ3�L�9�MZ��1-�`��
[B>ǃt�JH�.��b,*�˸X���%�2���/��������Ny�8�|v����y��əaY�l "sN��(�� � 9�������	�8�-<���,oB���Թ����l&ϖ�^:���ё����(ȎMw��w1y )�]�ۤ0���vO�v�B���q�*`��sS�b�mmѝ_(�~N��x}4�+	��?�]P}����2 4��T�ТU�����.s�K���C�ځ��񪂣ʴ��a��pQJ݋r��ni�gk�Fgg��L�ͣ�Z�Dy#�������Z���s�ˎ���(�����ݓ-<�a6 �A�c�w�FwO��Y�*�����v��E}+�V8�����e�2Gii4 e�����F�ltG�A�ri����H���8oC���-2N���#��ґ�Υ#Q��X"M�kjp��nvE9�k��o�F-������8�U�����!��T�"-����)�c�R���v�uȧ<��
�s��{�
�9u%%�sWzt�9Y˸�M<�(k�6�i�l�(���Ȑ�����L�SZ�o��X~��D�"�a���8X�ʺ�7�~���������/n�H{�"�ſ�N���9/ؚO
۪�Y�\*c�;�OO��� �Mh��y\���߽i8�pz�l'�>��'�H0mҕ�_s�:��t�0IOb������;ɉ�eRoj�㣏-�ǆ���K+$�n?����+�d���^��%_a��*���h-#��E���ץvG���O�@�a�H�=t���8�]Ü�L�g�AQ"`��RJ��Ʊ���d����&��B�/����O�����qո7,���D���S�A���w��Tsv����s�r�����]���N��*p8;3�����x�ˣ��I�uR�\ҘN���3�^�6q�o�k�ſT=Q��_��?aP\����[
����F@�Qu��8G̎!!Ɋ�׬�bd�+U���j~4с	Wc�|i;��Y��S�~<d�K�� QZ����"���0�̔Cw��4�����SY��*��2��s-B�=��o���BM�zj\���lUA�_7�R�W�NQ��An���m��c����+�������;$Fגb@�	 ��
���s���"o�7/S��ͨ�.>~A�-J �2��?���2ZQk��,����=�a���<�ߥ�N����-c�{��`=m�i�	�[���w/�� �OE�	 \MG/{��r7�/o��f���}���m������wc.ہ�(Y��{�Q�FF?^.��ܶrTp��ebb��P�W�s_⅑y�}�'�Hdd�!j����W� ~#g��ݩG*�?�=�h��˩�r����ş>�}�_�=V)_2�Ҋ\OOc)�p�����oo��ۘ����A���<��5G//;,���!Θh��Ң<�va�����WE��̣$oNjiiAۆ�ڸ�R���{���$k&�=\:r�	7����8<\�ҷ"XEmÜ6@�j�V�0�мx���3R4�I� �z�����f�w�7 �9�Y$�d>_�~
�������RhD7*�#��o�s��Q�)��� ����r{��R����S��:�}镙����mqW�`�l�6;���vA8HF�
뮤�!9.���H`�+]��G3;x�ڳS�Q��(���pn/�[q�e��ޤd>���Jqi*�I]L����L�(q����]lW�������'��A��_LbB|���.ALU� (ћ���j�!�1@'�K��5�BTT�X��������b	�T�*,�i_2}N�nV#�8��N0ɅY���`4���k|n�J>�=����w�\�S��.U[�dK1%9R�jeڡT��|sb�JbӾ/���=Z�����R�f;��eҁ�(�Bd�Ez0��o�,�r��t�Y_8ߊ���wn�
���"Y{��/����
"R�-�Av�6=G���,[7����K�=],������ ���0�5e8.oSy�ק?g4��F)\	�:����6	��;�>�S���W�V���V/���'�HInS ��~�|9JO_���W�)d�?���̓8��X�1A�z��P�8Z_6gQE�N9E3D.3@і���Gٓp�9ts\��$���Y�O���"Ɩa՚l�Fn%%*X~��|�1���{�;�;��n?�,Z�|�W�_��I�j�B�	�v�����+�*-�d*S� F�	��ε�`��w+�m��g���N���c0���em�^ةf�L,����E�.�IT�U&#��f������ў��ש�4b�
��(M�?K��Ą�g�N����͛7�o�q8�J�'f�yN�m�NN_t$Ԅ����M��f����(�<ds��j6���P�2[̔��"D�=oĥe� ��=C����_�����%���A��2����7Eoz}�>HKK����y�MOO#�I~�%�k���[uhM�!u[l0\��_;R��K����&��#Fs��;�!|�߇��v�<:V"�-�"����ڬK9ݭ�E襤���7r_)���d'�_�t��$���*��R<�y�a���������!d��fSㄺ�.DV�+Mm�Ob��<��F��@,�I��xl3{tt��P�4ta��Ȁ[]�++���2C��9v�UL�1#����y�7���K��r�z�����/�K�`m�<]@�@'?���Gf@
�Xm��$���h��(���ț
f�Y���o�ӯ��Yqqq*i��ڥ�Jw�u<��m�DfK%�}���NX�Z>+��y���z���ȃH��+Z����%R	��77'kkk#[[��q`}���$e~]]R��	����"����[�="Ĺp�?;�D�uu� ���뜔Eo����Ï�4�L�s�v������u�ذ [!����9E�C9���@q���\�vz��j
E*�w��GD"eq�W]�gL��o'˒li���"���f?�Ɨ�^~����5׼+V�.�ao�x��"�FP������b�طU�f�s%���(V��i$S4k�����?N���[�^�<׫��˯Xc�l�������oN��q"E�uڷt�|�^3'�@�W�!F/;�I��o��� ��!���.��f����iC-����&��6��:����G�����'�~t��o�E��]e�2wRoD���<Ue�鵘�x��+��V�]�X�g��J�{9��c���$�>G�P	��q.��7�?��u++�,����]��jy�0n�5�VKC�N�l�q�߀;���%�+���c����\g,Ȝ���Ny�y�g��b��(m0��*��2_SBv�?���a=�2�
������+Hi��!��,��-�3��oT�ް�}�iYW��]Wx#������|�H�e��Q%����_��K,�����h������>��9�Z��S��1a�(bbRK���=������L�aO��Fe³���Z���l���ݛ�)n���b=~+�9( �|G��6# �x��w��+e��]����$Χ8v��<�y�������H�TLL2���3����� ���~Kǲj]����������ݞ���>�(��F֣�6���W��Hi#����%�;��rP6��(��1=k�'ȉ�fޝ�Uf;{�@u��^�qM����a���	�I����@k�H����X[�'
؂�|���P�}�9�^�c~��*���Z�`��=��|����ƫ?�}�������u����܆�t�W�Ff������I���&��f9
��-K����0e#�9x���=�{�3�cb�����г��xO=��"�(Cjq�hL�R��+�P��a}6v��S�N*�yg���&uC�	~e)  N���I���#ᶳ�sN�t�e�!�n-��� *7�̈zu�6@�����s�"ʀ�z��P���,`ڀ���z���i�˺�&�xK+�Q͎0�o���'��A�}�@�$�o�0���G�*/dbFzP܀
�5��EE���2�|�z�x�'�%k�Kc�/a-�i{~o�x4�������J�;dpp�pJE��S*�~�r�	�a/����8k�/6l6Ҁ�Af�:E8���ޅ_��_�s�;z2ˍ���5� ��au�B��{@[`&.�y7��"�S����)T��Ǯ���j	'Z&x��L�]0t�A\g��SS�:�.���T:A�	� �%SRO:�<�_⳷�� �{T߈ч7x�#�z��+��������3�&��{u��,������c9�*
L����Au[k��h���G��Ŕ���s��zWW\�t�~�z�ƾ�&l��=Q�+:rr����8���/8�"��ڦՈW[� ೛�7���3J΅|��ώVd��vS����K�t&�u�? ����V~8<uu�u����Xs,W`���9���m`sظ$'�_o�Q"޾�Z<�N�/--ߨ�,g������R��C�x�p�X���f�[q
BD���x�4�ݴ,X�[�ݞ���0;s#�:�X߱A�}��v�^G�U���75����l�����A7Ј?I<&W��
���:����z��(� �c��x�S#Ϧ�Fl�j:�b�<ځ]��u0to�b>�f��!���zns5M|��v�*[���(ɝZ::�?�%׻����xxx�b��C�e�s@)	an�<���\�~��2�~8)���Na!Ҟ\��������h���}��^AE:���R3���4��8_A��萴vr�M�n4(�*��7�ȶkZ�p�$���)�|$r�m$m��%~AFR�Ï\8E�9�]7Y�U���:�џ{��v��
fY������wXXY��`�,U-ՊL���������]��m�\.��#-my���6)1	�Sگ8�l>_bI+ޟjܲ)�����|
�.u3n�ދ����5X=��~��qXFb-b�aʄ	B���mq���6�L��כ���*L�(tc���W�]"w/���?~�$󈧜vƁ�@{�[��6O=��ӻ�|2hSE%E�1�'��"��Ԝ��(��xS�~;����e���Q���x�l{�����Mxv���~D4��\�����_�k��-�S�@�h�i��D��� K�U|������s��Me�s;1���C�i_<yeI��r��>�q���)Jێț^ƻ�~=�N�/��6�}����3q=���[�=�`�!�.��*Ĳē�@'����P=u�s�EV9G��+((���pq�Hz���^�l����)�Y���$o<�]��5f��o�k�;�e�D�;j�S�Km1�m0���[rc��Q���2
�k;�C��^���~Lpg�0�dnn�,��8��H���44Zi��u��U��J����Q{`���Z�p�a�3�]I���`o�n*V�_�"ط�� и�����6Йz�oO �[���=��<�qOy��q�����S_Xh�Y£�H;����H_��j|��_��Ĝ���]YY	�s��A��omP<�!����#0�nQ�v��o���4������!-U�%�������:��}�b�_(7�U�C**h�Â�=���X݌�$����Nd9T%�گ�B"�h��rR�	X�O�ABUC��@'#���� �Kl�`]�v�h����PL�Bm���D����n���OT+�P�C({�����?�A9��upW9�H�2=�䈾G)���{��T�B�� �ł��>Y5n����濟����s��q��|�la�^��A f.���t��t:� ��2���������i�{]q�П(�?�;���ba*����90 �����a����hl���e����3��4�a5`3Ŷ�w�A�QJ��������'a����
`ʱ�+^����W�W=[�����g�

�b聹I��Bgh�C��y6����} ���qɋ'@���WXE������O3�h�F66�a��U�J��5��ܢ����ɒ���QD������L�L�߮;J�:dE�ue�v�5i���;���o�ޖ�b/��߮W�YJ(�=ϯY��tia�>dc�]^���׿w�ji�1�};Y;��VQ�+�^EB��x��D�I_U o��n0���;� {é�OP*R�`�l)Ը�Rc��T���-W:B�pk�ƀ���_@Zk��'�X���vVv��%�WW�Q�[Q��r���`v4ʨ�0ޭ�˔�t�B_�"n{�z��ث�.N�'f�kUc�����
N��֯K��aC���	������4%&&n���)Z�&��N��Ռ��ñ�X�����6��#�\�?���JI1�5�F'��������͍�ܒ����2�.D!�K����E�  �k�f;"�~H���'�kuO�jV�T��ҩ��1�q8?�֘^�ȁq�r����[����a����)�X��+�0�p���<�h �m��{�4�L x�'M^�	[���|��l.|�:�5J�ihb���`-�ӌ9MU��Ý��J ezU) ���|�={���]"��[�|�s7��Z�D��)ݼ�|:܃C;��y�^��^�̋
b�}�X�DY�mE{�sK+���.���=��y��hh�yуҏ�hc��H��ϧ���%���A�u�B��c�.N�m�&͊�	v$��h0דd�DQy�Yy�9��*?��V���?~h::����x�9Xwg۴��Y��Z֣�x,���me%�҉:��E���Warc���Z��9Tr	aOE������w&Ϻ[u���Uc�[�M�rP�r�	�>;�m�2��&�v�7?���$�#��`�_�$�-��V�k4v�X!&�Q�CI�kT����1�%V6���-�(`������ۆFG�Pj�f�	���]�b���âu��>m �{8t�/�3�?'��CŤ p��yг����s_(y�٨R��l��	!]�#�]|}j�����\�{��Xm', G�=�6|��н:��LEђ��EH�`Y<�B���R"Wr�\R���v�K��	@p6 i��3��(�ͽ�>v��0^�3g�,��ѣ �U��ʣ���kk��n�_�F��=~A?V�A�C����uG��p�AS8��;��<Q�f�<�<�P��Z�$~:�<N:-���O{b���zP�K������X���������y����	Rń�
�)�aQ���
�����޽{ ��i�x4��u#�|���g��@R��\���?��o?�^	�&��4�Z�-��ݕ&��q�p�<��Þ�_}��{��7uri�S�>n{����� ���6���D�1V֫�yZ��_� I��Y_� ��ge�Jd��Y�U���X��Į�����Z�X�_���l���?�"9�� �M�w�����O�PN`��'�������T���H��J8iW�P��ԉ�^��4��E������4x{No�	�)~�^�^���� %W7H9l�SbV�J�{?�|�I�Cj/E��{Ɓ"ST����h��D���zR~Iɰ��ڥ��%H��N� ��e|P����%�<��5J�á�&�*mb.q<0�KO��&X��׸�+�$y{{���ߓ�$I.�c��|����@]9���P�Z�Jc��%��K�}�c����>uD_9c���
�J�S~ު1���4�<8�E�v�嵦β ��S�2d�j�� e�d�d�yG�
ٱ�bX���W�g.�F'/j���g>�ty��-�E�~
�o7#����
 �AT�(�@x\��	�S~zz�{�_fS�pCE��Tzf�=h;$��OfųM1f_uѷ�v�7E����� @���xE:��Vx`ǚ����� u23/il�ߙ�
��X��#���Z~�4�4tt��i �GFX��4~2<����Y���Z���߅�^W;�6�.���v~�Gκ�-\SasM��Q�8W(�ĝq�KxC·'�Z��,��~-�gs��,.�\ۻ{hk��q�O�)H��%x�[9�(P�Lm��e����mݑ�T��j��ʄ<Kr��V�u�f*
]޸rV<g����M擛�98�ʣ���YO�٩�u� 1I�#��­TW̣cc�B?��\�*,޶��^nַs<��J�a��3��)d叽�����R՞I��S��㩥�{�2������ԣ�����!H�n����Qe v�OII�n{�`�ܨ`V�iG	�@)ł�M4�͓�������-s���tU����L�0>�ݱ�Εm��x))�����ڙH袠dwyq�k�r�й�[���L�@{u1���mu'I�229�lu���i��D��JY��}��#n�#�N�� 뢾�M;�HG5����E_����~�����Ai,|YJ+B}>�c{����[,|>/bf�O����$=�VP|"�zl��`cﻵu���3��}?�����_�ġ�b2�x���sth�E�\����8~v��$��GB��8T�!�5�e���E6��h����&cɃ��J�M�.�X#o�M��c��5�.V�q~��5��n���|0h��T�n��Lm\Ȝ��2z��F�gt	#����Y��1��8t�����o���k�/�`WV�&W�?>?m^5��� ��z�d���C`>Y3�9��*�W�id���9:�ߋ�����į�����6V�V�+e�M!9�5jt���X����9�?�Ф�����#�ư��7�(	�|��C��xmF�]�ӝ�.�JO71���lMF	2�����T<0nq��U��v�1c�ފ.W߃�����Om��o�Cᡫ֒\��5��VCe� zoYsss�|�+����-��䁻8��4�י�#I�t������z����|�����7���s�e ��Γ'㩱>^�y����C�^E�R���|��C��;�]�i��n�=&e#��HUGǊ�$�x/���㼹�9���e��PW�ω9�9>�ӚG����^����Ο���WĔ�?l����سtgɊ�F_��5�"��L�2��C�ۄ��;�d���Ӄj��Oҿ�bMP\̑�σ�����������v ���Lj�El���4�g� ]d
$d�F������2�K�1L��K�-_��� ����0�3�Nߵ�.�mZ��4�d�\�D>���u����$��xhZ�9�Yİ�+�>����{�NVtT�#I`�������#5���;�ѵ/��ĤY��W9�wV���j�-B1��CQ_��� o�=�s�_C�[�Lt)�Z�4��~����[(5����l� |�Pc:�q���V�apHǸ(�`#'v�9"NF	��u���`�R�N� �:g�E��ho%�����ŷ��z��b��So4�q��IJzM�K��ߦx'W�溱z�����w~��>�����'����d����y�(�~Iy�'��O�]�#5���D�%�{���%A���m~�İ�W{�\����l���A'�tC�0�Io�����0���Ϳ �#6�t
23[T��[Kcn(%����>D���r�p�"��+�2RZ���������!]����7ϟ��@E�q: /���)�?MN^a�q~i�b�R�eveR�kZ��p��8��n5�$O^$�u\V�F�:��d�J
������������뼵[��-���Zͬs�_����|��"G�D}rS����ޱQ�9u��G�����ӠZL���*��|�F��4T뉖��ؖF�����(�
������r�#v�с����LPm7?'�A�ؼ��K��l�>b.��b\���Z�,��� �Ed�v�E@��k�j�LK�fư|��+��E�B,m^��8,��»��j1
JU�;�zj�7�0?��lJ44�)�Y�p��>\V����s�?����u�9T�1�΅*�PlaY4�(T&t$�$��
�^��i�&T���S&RAס^t�^|lo	Uu�^��S�ӊz �!e=7g�R#y����p����7!-EI,��Xq$���Di�'�Y�L���6,7[4cטF w�bXf�å��ӏ�+d�u��;��䰸���'��U�<>����h�):+޵G ����E88�q�� �,��{�Ms�;)�����N��[�C�U9`�{{�Q<�dO�>�^���X�h�OG�VE�H�L�n(�"�,QEq\�z5⩊��~�uu}�V;��1ӹ��A@u���~�����V��}mʠ�zê�ZUk�ݍUjs���]
n�k�75�mU���vě����ĉi���9dco/ #c��AK`�́X�+(���7�q���lv\b�S������܊�A�kV(�@$9�O8m,�5��ݏ�$�����+�+�l/�'J͌���^?]���v�sc��Y�i]� $�)�ݸ	!s�P4�nx)[j�Do��.ه�>\����&P�v�I��K��*�Ҍ�e��e�B0hog��\����L�ih $T��\���y��VJ�q���\�Z,�@��G�x��㣳@��o�F��=06��W�Dr=u�n���6{�bbرf�,ZIac[j�2�������ht��3iQ����� #��W�6��5�u7{8�E����V�7t&�9�mʷ5ǿ�<Q�����]��iLܣ{u��ٳP]T[A!�o4H��� ��Ĳ�ƀ�;������j�t ��3~A[M-�P^f��S �5�>�w�}I�LN�=���P����fck�;�a��q^Hl���>�]���F�`f��|��F8��l���/J���]ۇ�֦�z(���۾�|G4}��BWn��S� ��J51U$f�^��ɇ�����5�|����Y���A
��e$��C�w.Ć\(�&p��L5�ڛ;y��}������,U�/�b93�Qt�8�<H��M.,�� 7����$��S�ZD�NY�O֮���lTgo���D8�$�&�p�ʦ��]?��<�D�#=��UI��`:������F �7��
��<
��x���[UME�Е��2�z���ϟ�⃙ 3��%D�U:
�O��!I��/fgg�k��Jj���������PI��ڏx�i�ڑc=�ު����d��v�B����,$����O����0+�۬,����7��v������{�I�Ц�P�|RX� c��V~���Y�*�3@v�;��2։�"���а�E�XS�	��NBe�Z\���G�E���S���e@�&n8	d�m����������xXa0]_��֖�p��^�K6�%��k��t�"y�N[wߏi���W�{����:j[�L�x�QH���<z#�?E�*�I4��`��q�ߠ�e���}������15��E�g���U�I��nwI�nC�Zӊ#v����{�ɡqzM�OV�;\G�@���*,��QjW���z������(��v)[`��ٵ���t�w �דz���;�M*rkR	ijB�c�Fc}�O�P��0��S��&D(�bf�߼gn��g��W7n��m!����j����D~c����%Q���@�R�|y�t��=ty��{�z4��0$� ����y��(㬹ߜ&���OC3�8��ǝ! WP�����T&q���"��_�� �.��ģ���]#�nH1��v���g����!�@�d	�Bz����$!G�ׯ����':��!qxR��:���)U??q�ۤ��Y~VJ^��bN�����ySq=Q��>�Q�e�2ν)����vpȜUWA�"��u����"�j��]8�;1�Yekn��{W��Z8h�i���! S��kvD�^P�+:�t��F�g$���H2 �:�Dݡ�%t��Ǹs�:�����n�m�GAqq/�Իh[Ԙ���P�C�	d?�K��H$J��PH�"�o�79��]�K�:N?hO�`�S�pPS�N?\�h�]}�^�Xz�����F�v�pO�5��+�l��Y�+��Ȟ��6d4߁]�G�hj�%�9D���][g�z�T����ד�,�̝���ͽ5,��,�ږ-c� _n��Elj>V���P����tu��/��s�HE���=��---
]���HZ��75���.0B�FFŀ�A����������}�~��2���|�}�*�q�)\���}�-��[	 ]K3h�{�����p���ܓ�/Y�+EzVTw����ј�h�T��z� f?M��C���o�.�ņu� !c
��c�GF�0�{w��
��L�L�
-��a~����
���3 ��!W��Ư&aU̙���!l�������M#1a�LF$+v��S�LnE7!!r��J|�V8�e93B/nG~:���P?6N+��U��%0�?�ajCF9��^���y���\�����[
7�O�D$��ȭt������@�҅��C����ᢪ	��F4�_	�9&;++YNNN�i���F	 ����e�� �n�8a1_!af�Rq>�S�R�<���Lx�f��0�5�b���e���B��7�2xɭ��Bwe*�_fMϮ#�U���ʟ�&(��e0��9>9kJՠ.�YE�x.''��ߥ׏�C�uE��SP��Y2jt�~�S(6U7�J��������THv�R��S|��4P/^�nN�Ra.���%��Y�������ʟϋ������֟���88����7�{/ 9�h�m����k�m�o��+�r`����re��5�S����c&?�������Z-����%�=����ȼ>�����/��^���zhh�Âo?b���}��I9u�˃�~��;. �?�'����A}%�b�xJ��+��#ԡ9�I��ݴ)go��d����'��<��P�㥦Y� ~�Dv�{A�G#����Vڵ��y��ݷ]}%_~����l�GpzbK����x�1`�.݅�K� ������֏�L�1h�<�Z���#�x�r�;���l7�WN�.Yz{_9��m�%�2��Pű�[6{}�#*/S��2A�r��X��w�^�-������ȉĿ�:Y	�e	����i��^K�~�۷�l��U���$����:oa�f�
m���R��qR�Ƞf �ݥ���0��|�ug'���'�Β]w�^��.���0����Ǎ� � %C�b�<�{�8m��w)�@�`Re�L������Tg�l�E��&��#�Щ/U�&<`�X#̾5لڅ>�z�j�4Yd�2�N�|6���crXhߺˣ`%��d&'t����.A��5$޷mq��"�/t�!sv��]���i�JWI/5{A��-�⫛�� �۴������������5��0	h��20;�cş�%���k����P�+��h��v7]o~ɍl�c�a��	ǀ4?���5����4��� /�b�6�7���lP����nM`��p;X
o�x�7ܕ����f�����K�n;,l�m<(7؝}7�)YuDZ���ɽ4��e���RdZr��(b[G�8�̈��OE�O�����t%�5��#���c�H@PP�����\;�v�T���ں]��}FX�
��������z>��.A�q^(�y��.�&���7#Y+2���}���Y_�c��r�Jtg��_�\��ߠlo�Mv�����Q�G����/���?mFI�Q�8��=�FH8𝛇GR�����B�|�S���q���á����}l�c����Vb��B�^�\������̭x<�`��g��͑�Ӛ7�A��Hp�!BI3~,E�ѻ*������� ��@�m��=}\�����H�- �'S`���� k��S�^X�.1,����;]����MT��=:�*�=���5�E��.7Ut���.r�XS'�ݍWS��i�E��d����u�T��-��0����{��h�݄-��&�tgi�O�T�ƣOa�P�/{�N<�M��A]���-*�A��	LM�����j0B��
x,�Αdu�zQ��*z��γ�׻q��o��
o,�{k~0�ڸ"�~�w�+�jdz�j40��/:��*}�V?�֞���D���Ȥڽ=r�GrK+�m��91v�G10��������I 7�/?��l{y S
���:hqU'����'є,#^���c�̩g�_�����*^�.*�4��7K�NDA����l�$�k�lq��E@�=�H�(_� g����t����c����h <��4 sZO1z@�	a��EEE��W�**+���Q=��80,�������)�R����n�����,k��T���>-�	%[��G2���Y8����r��<7H��b���5�U��)�k���i���OyHmF��+@Dˮyݜ�Y�����uh��R#��Znnlć=�[�04��wV�����t:Di�[���������<K�?�w>�9��9����5>�A��c�̳����G�Np���p&o�c��_��]�p���	h�wT��\�ؿ&>�ŅQ�_�#@=��KwPEf��r���X�!Y�UQF8�%��=���9����ٶ����N6�=���W_��*�?�	%$�YRD��Ai�X�DB�S�A�C���i��]����"~��^?�����Μ9�yΜy�Wgp���s�Z�}G=��NMv��)��K�J��8J\gt����w/)�o@��g�q��cD�7�&����}e�2�`��W�VHF����Y���k_�?/ѫ�c"V��6������Oę�PR�����,'x��t8e�Q׻��G0�ȫ=d�s�bmOً`JO=0��y�V��oB��=,)�E)Hq�z�IҫH.��d�m�,��hfkcm�}�5��~5!+�����9R���WT� ^��φ���P�����&���	55d�R��tX� E<�|M�����
�w��Ԟ�|z�Ĭ���'"����$�}��뎞�#W�yπ?2��k��������'�ɷ����l]�'Ǆ>S��.�;U$��帉"Sv��VG�|��2�vh�w��ߦ�8��L��w��~�Gt���TW��)����u��++G\Ü��	�@�Q�*�U���;�,=���ja+X�Q�(�(��H�ȹ'�b<����1��'�������D���?�-�T�x9�k'��҄���}i�~Af/C��׶��n�6���Ю�F�y�d��㦔Wb���QW-G�Hs�g�i����<:�Dz���Hs�b���M�Ν��;F���
%2WM��Kݦ T\s�4�$��JZ�~O�Ù��k��5T�ʁ�©�DL�`Cd:W�cc�z�4�2m�t�i˄`/ ��tu��q@g�����<�H�U~����l�x����\5 ��M=#�Nv��,�*`ד���/3)��:zId�z/��i��~}�w,������6%�'����w�1���is��$�uz��.�/P<�ƱLw~��(;;�	�:�v����<�0J�*y|k�\5q��҂l���ד�21�`�K33�mJ�Q��i,%��O�k�-�&��Qrp��ay1$�;���u�/
�gy�M?͇DҦMq����{�!]���[r�3�<��$-\r�*�����pnJ[�`D�Щǥ~����x���{��̓�������h����GR��kv-8�@n�2)�4��uϰO���T��Ȉk�|�S ��'2��O��XܾE!Y;^Kn$����I��f������PWq��M�(萬�� ��ëÊL�����]o��׵rx�l�kc���Hx��m/M^~��M"��w��"����h�Mk���g��N�3�^�Kx�*fR�q�YX�Y�gΝ$틝+{v�~6����� �sC��cWAbx �	tQ��V�p'N�W���ٛ��P4��+l?�(6���n�z�6'5 ��^�]��i-�6�g6�უ��j.8^���\*#>��Ǟ��2�Nֺ�g�m#V����\���ù'���=~��^bXR���a��3_/,(�q�E���'dfV(�ߣH����b7���0�rƈTy{H��B�C�Q.ͼ.P��Sذ�����i��<kn��� VOU�5kt}�U�"J��z�`�\C��а6���eۇ��#���Z��y��,`�-�ef��w1��y����7D�r��o�mt6� Lr���<�s}{�?�3��A���]�i'�fӲ-J"ojWW���҂Z��;��� �`���NJ{k����d�?���Q�XIOBJ��ɞ�K�6(���b��n����[�#,���:�--6�5q�2@�f�jD(��tMhyu���M���� �d�}���*o<�
Xcf�E�L�B��,��������}���#��O>�C
�v:|�g۷�E�� J"\꿧Ֆq��ui�kx�J���5?e��p�;���Qr���-�	���k���+���^Ű��g�F�V�ԧ���)��(9���$`���؆J�L��s�ز'�H568iz�5�{)��̺{������8�����á	���)O�QY�9��6ؕ�`�4[y8�ΒDy3�o%�.��.ץo�b]�^V8��3�:���X�x��V��=�_�|T��xg�WflSě�=�xRte�,��c�o^~�Ggr���X�UJ��}i�;�R��� �N��E"���&h�T�%˩�-�8t���d~�/�`P�r�'%�M,���S��-����B�d��=���az�7������K��]Ǝ�8�f�vP�%.�;$��֜��?W���k���u&˩;扟m�b�&��Z�|^���aeeb��M���4���5�k�`v7R�7<�0._�de����2Q��8
��e�ŭ�6�V	] ��n���B�3*ؾ@{��n(8vcT�B}=�ۯ�x�����˂C��v�5nypK��#l����R�\^yGB��mʻ��^�o�#�؜W�}��掆:Лݕ��Z���[����(4�O��F8�Ngtj�8B�bn��2��Z�xM@���� ��3�t�,H%'^{���駗������mm�S���4�ͪ��F_�?wl�j����ޑ5c�0��O�7g�_��u�<�]7Z��;��bз�b������VC�O�����.�������0Ei�5}���t��w7���|�qά*����ő���+�<�~A<e=l5Z��^����K���^��g�r��b�9�M��g�
����}pbPߟ�?%j�Os<�
�(��L�di��E���3��؏�Bஓ��l�T�,F}2a���!�_���/�ȫ�R]ΒC���N6%a��G�����I
���w�XHC��� *;"�:;�i>����+6�ʻq�:`�9]Դ�=4އM���j������'sU-!]ָ�f���K��5���Qؽ���@������!0�C5f�m��ڦ�Z�C��SS��o�ѝ�(�����+�Hkf����	��)���x��^�6���nd&}/�������I��I���pv��V`r?�aJT�0�����W{;�-�;�c��
���q��'��<�rO�e�rUMH�'kr�T���^�%����Ǐ��Q��A�.�?�Q���Յ���gs��ܕ6
��H�KP�c�:n͜X�͉����x�����Z�f���Lja����9�����o����sF����=خ��Jy�e׹<?,������ő�A�1F��џ�����~[ݦ0��C�D ��6Lc��#��X����j1r� !1�Wo@邏����ݚ�y]��/Vŕ[9v���dӥͨK�ww	�����U~�I1�P����j��7�Q�x�S:�̐�7�r!����'ۤ����n�ov��	��*&7�T�d��2#����{�Ħ���nX2��0CI�R}0ť�k�O+�Z��,L����V�%�;�R��-���SL3эv&���R�V��J���(��:�w<��E킻m,�y��-���Z��C�7'��s��p㏵���>Ϣ�9X��d	�0�)��&�
M񮷱�ǒ�I@ۑX�KXԌ`BeJ�����.^�Ձ.rO���L��,�}%k3vύ��+��Ϧ7�w��OT��P4�I�.5������>4�2��Sڤ��[l�:<K����uK�kc�Y;n�u{R\���md݅Gs1sb�d,�6l	��:��U�{��
5�תTT!�'���,�m���B����5��-�C!u�/��=���4�����mK�_�<.�*M���f��.`�iƱ��K-#*����y��3LN����~���9&n�X�9J������O5���E��4>��By6\��N �r���SѢLq_��]cl`w��Vz##{�����	'�=�a��;���]{���#V�TA�,�W���1���L^	E�K'���0��`:��.�:P�ۧ�P�~,s���\�b�~�w:o����-���q��w0�^H���s�^~��:jb�^�?
�h���V��0c�lBccF���g����柜S�w���&l��z�(��g]���8�T��i=5�O���V��zs�?�t6/��Ll��<�'3����A8�<j�k<�d�ږV��u�l�.�4tV�(Z'̎I�_��>�8������,��K��vv.8!nu-970��eom��e� \L�$nP*r��(�`9i��i�q|y���N�����Z��u���'/	r �;jT4�R���i�K��G Ŧ��o�R,�Y���
�G��"�nb����N��o�̓�i�,+����>�Y2�Y�6	�)�u'X��@	w�� trp(^
aX��c������u�Z~�L��ҭ�t@������;�n�yiDl��l��6
���}� Bu��(ؾfS�c2�~E@������:�#��kyq�`qK-l�_P���������3��<r���Y::�~�o�p�kQ?
�<�S��<����W��wF���|�B�7[�:���1���!��#[�0|-�\�kv$EL˥99�&
���CT�j4�)B��+���7��^u���#C�3���6Y���R�e.ڟ�l���d��>�ĺ� 
����Y�(`����J��ݞH������:�Ɇ>�D�2w"�VEf��R��ѫWG�'�8&?�B�.=>v:���ȑ�i��ƻ�Z�S����v��m�c4����N��{�<S����N��y*?�9�G86�`ѻ �B ^Ƿ�@5Ns�5~h��V���=	�*|�O�Ǔ�w�(�z|@�Ǜ�rP��[{e�88�B	��s�0
�{���Z8Q�Q��$V7U�N,0.(��}�v'_���d�ϲ-g������kj�-��g��������}�.�V�\����bN.s%�Ae��)�F:���%�m5fkKo�'Hu�{�~1zZOU;vL�A��Y��p�|�P��fs%����Ǽ�|x�נ�Noo���Wh�������S�8�j�|��00�	xy
�'*�g��Iw����	���@�����ox��uQ�1�ۇRL���cP�����zܳē�5ν*@���� �.v+'2�/����.�)*�vh����Ǿ�j��d������_�ƫ	$��p�e�V���.�a��rP>�T4�ш*����!"���|��F}ҝ�Zş�������^��RXq}��R�zE"<�Ok�/��f=��⮗�������#��X�M㧺zn̜�h�U��c3kȠ�*R��x��Pt�$N�����/ⶌ��]�ё�[�I69T�nc_�p͉y��	Ji�ȋ��_�0�>W4�ւ�u.@G�`��4�3�E�r�3Q�T-v��'�%�g`��ݮaN���6����+�#�c]Z�Z!9�&��@X�bHhi��$K��}{E��U�B����6)���.��>����n^�s����k�����R�D�c�7��&j���D
N�����^VC�:�
�F��O��^�8�X��]%�0�I��n����w�ݓ�p�Q����
*�b�4�[���Ӝ��YSD�'��+Z��kQ��*��R�y�" �����
"Ï�{&�W��湄��V�.�@����	R"TK�zb���QP����7�� �^��j�G���Z�LG��Qou~����߉h�">�I���C��/�w��*������� $tO�]�P��^��<%��� egHć�É���}c��<�(:��#�R�}D(���HA���ø�_�~���3P귦�XR��g�{��Y����������-�*C�w��"	K���T�ˉ�� �>!��N\���f��3��s~.�-~�(a}�"��ܚ��^B���<��		���)��r�����~��Þ�~ s�� 8j�	Q���;v�6��"���y�zOzWl�-���&��]��>��1D�[$6�܌JR�<`+s��<[)�W�G�\C4����;ܫxe*{��fl���%H��;|���A4~&���,li�qC��ظ�n���tje2vf樾8�a������ɡ?F��|W�kȓ���h��6�ũ;&�	�H���~���Vj��k}=z�y��/ʷ�2}�J�'t��	Ҟ{ T�0����>0��M��|�G�~�~�mP�-k���g+C��BƫR�ǧmyy]�o�{��m�Qeh�z��Oa���V��jxP����r�Z;������ܕ���OEo�uqWS@�3�A{�H����8sFs)Om$�/��aT�;/o�������c�#����JL��c����P	��ZsqeI����Ζ�Aa����b�w���(��=�D1!أd
ʇ&�-��/r�k+�[<��G��TM�n��zG�Z#p��+A�6n-ѫ%������Ye����<C��T)���w��E{�� ɓ��� �Iu���É�XV����J��l�٬���Kq���/��E���]	t�('c��7�kbYY5@Լ|劢�`���܎���î����Ù��iaiJiB��Qv><���wG�Lc@�0s�t�%Aۃ� ���/���Er]"u˘��]��}�S��U��V:y��g�w
-'�ߗ�R`l�om�ޡ��8���F���Rt����)L}�+HLCU5
��ad4��J
���?d3tLș���#�f(���k�N���أ���>W�12\١���3��O�g���qU��<�]7t�\�H_�J���U���z���t����G߇=x w#��H�6O���+L���m=<���o߳rU�>R^~����nM�u3n)h4ZA��5�9�*���&�m��]�腕'���h�Ј��C^aᒑ5������li��;	�6�;�9Ɖd`����)�s5oY��q׮�}PN�M�z*�!�E�Of9����N�:
+�����L�-����=� 8Ȅjk.K- ����r�󊒲������h�-G���6KY��O�~�U~iV�C�?�B�Gg�[K��W����S��,J|��ɑ��i��\�o�B��{'=nyyy�LSUُNp��3!L��/fc���a��n�Xm��ɋ0V)�8.�XX�s�)�^W�tI�q��ɸ]}43K���G��aBhhF�n������b��R�wC���c?��񂢢e�-"�]X���|�Qt3��8��F�n��{�<s���f�s>�l'H��>f���ي���Qܽ�M�vV�rg<�I$�֝HZ��p������b��a,qrޤ�x{�o\7��ɍ�8�ʠ�zX��V����@���g��_ۻkB+LC�}��|��� s�Y�5[����lvCL��R�wY�����o��������$v %I��ξ��.G?:\h=rFID#Z��	����5���h�"ǎ�f�:(|��w�����Lpf���-}ym����\��`I	ｵGT�z���[ʗEm����pd��[��[�X�c���ǿ�w��������5��&�^�NY�SR�n\:���>%W����^t�w�(+5}��13#�(tFݪe�;��u��p���sؔH��KqCXņլPW�"��.EÏ�����?�%Ɩ}�l�����*�R�Oxdf��'��"��>K,���|<�.�|Lom=�
�
q�>���{(��7>���Ւ�m�(@9�v�Ѷ�.\�O2�u�/}���p*��垞�V�N���Y����/�O��ygy�z\3^�f\�_�G�O4e\�t�n�3�j8h��C#M���;�̥D�NR�A�6���YJ<^���|�	gTE|vS,�E��.��$���m3���~e��W��/m%���c~�VlCH'�� ���6�t����Bŗ�$aVy�阯9|�%P8�������B��1Y^����rD�T��FN�
�����.�ܷ���1�mz��I'>&��<�5�t�\��`�ݗܬWՓm+�f��+Ԛ!4�7�W��s�챠5��o� 4��]�`���-~�n\�ck��dm��Jt�j0��HEl��a���0gݶA��_Wf�0������u�������X��b�2:^�~~��h#�^�x1D��L�&�����C�PX���b3j���A�ռ��Pw�aig�z!L�06�Z��r�5i���)2sJT�����ntF�����C��ABy��bܖI�<_���<�zM߳C�c��E8b��i�:$�!y�Dv��[���+�6ϖ��t��ᦄ���Y��'XE�aS��o�M���f��� Cfk�w�K���jb���WQ����X���܉pqM�_���y�@Xm��
���H��{�$��x�N`lF,S�z�=���/lmG�S�>_H�TU�_>n��z���I~Dp%�.a6GKm��5��m��HɆ_���K�o��P��>11"r�e�s%"9I��t�i������&�ΰ%�a&-͖�%k�m�ǎ������Y��/ x=��႘�='a���Ld���\���EȺ7"P����"���?�=��=��-:�Kg�^��6���9^���m2F�o��P8��\�+';XtI�Û��^��:�Yg��%���M�j�m�g���8�I	6���9X���s�2N��o�B�Q�����ņ���m*���覾�HHI��et��ɍHs��>�suB����vRc3�n�;f_�#��͔\«�jkD�ˊ�������V<E�06�.�$B:)��F}~�3�4E����P�b�;#cc�K8�h�tS�@Y�(����-�,7���jg�t����N"�9I�׷�7���z��b�S5\�ss�a��ϼim�q��bB�K��\n���.�fU��O�U��s4q�bk�,}�� .֞P���L�˯[�:�e�8�m���Vz�ڣ=�F���qA�?h���7~���iC��W��O�B5����R�*���S����`��NNN��ЛU���x�f��l�� ߤ%�	zH��z�ߧy��p���M�j!֢?1sm�L��'*q�{EO��f)n��x��S9?��C�S��3�z��Fw0oZz��.�(�W��i	x��s��=k��i��basG��q "M9��Tۄ�%'S��U,�ޅmz@����k���cd+++!������r��pg��U�T8�_��B"�p�'�q�O���iٛ���`kr���$�I�0�	>{5���yG����nN\��/�3O�k��}@��D[��\=��V��S�G)Vr�Y�����C��'�[� �O�J�Btnmo�<�]�V��N$jiO�>�w�S1�3�q�Z��Ҵ��quY�:�K�zl�����{sAK��˼#7��9s23O�9h�F��ϵ��ׂѢ�P���7ta�7q�o3�N�3������{��ш�΋����FX੣k��)����M�ou��E�S/�F)��A"K�
-Ặ|)��IC�`|j��,���Bֵ�A�W��d�b-�W� AĖ_�M��>s.��RF�`9�Z��,L���ԯ�h��z�r�=Tkn7�:�fz+�6X��������4�'z��8�A�y����R�������ZҟN''�� �*<$��#rn��*����Z���(�<�H�l�iC�9�J����Ӹ���u������3�13�4>=�y�q��5)�^��Ɋ?X�!��0HV�>����/��gff�R|��K�M&�ʃ��\]G�L)ޣ�i�=,	�=�2=��J���0!��p\�W^؞�V��Gv"0[8q��`^@��L-�#���.�@�_��'�����\e�2]H�a�O����h���4���]��څdK�:�T^��ƍ�vḷCB�/2�E�-��i���y�ڛ;-*��p1{����455��J���>j���`��~�*$����Q��P����K8cw�JY#[0B�K���o�fjj��y�<��P-^�1���f��$'��^&ك�!��V�G���8�GGW����o���� %��-9��oO�a�"�8��|��+��~�
?��@2ZV����b����]��Ǜ�K+]_�XX�>����L�އ��^�*]��Hf�����GvrQ2���T1�$dd}�u~����/�s�=��Z@Vp�%.#��l��T��=8����FIB�p�{��f*T;�Y�r{�F���ж֔c7i�2��[�̈́R.&�i)Vƚ^�~~0.�\P��|��?o����"�ǧOuс�z�2	|[>tpS����:���0/O��y+$k8�*�˷o���-�$t�s{���A�7�B�[�=ys ���r;��p�����]t�l���D���AK�ї�M�hƪ�܀6JEZ:(9%z[�?����n�Zؚb���D>��塳y �ڮŦ8!��p���\���I+P��h[���>�8�`3�q�W�aդ$��͖�	}ʜ����=����o�)4����_��g����\ޝv�^ꍃ����F�i��+���I�^��C}��
�l�xxV�+^���|Ms$Nf��;t�0�Y��=ٞZ���;/8/�q�4��s��B��Ѕ�<��&��G���џmMCC�񵍍��b��,���Sر"������nk�3}�t�.zh��4(N;������]\�=�$���ƥ��M���6ڊ��\�j��{Ez��nk��KC�������<���x:�q�}G 0:�v�Q�$�j�B���� )��=7D���Y���rr̦˚,��h�:<^pP؄��v`6V�#�y)�r}�w�h�M��M�I $EI~���X�,��<t UP"װ4f1VRu��pJA�u�wy�V2�a�����}x�@�
�C�x�Q4�#�lS>�_�y�M���Y^�m2ҧg��$���=e���Ҁ�i������>�H$�-1�G�g�x�"��d2�\yۓX7�FgA�S�hFS[;?�۲��^��Tyv������������������Ʉmmlz����f_����[���+��a'k��w�@�E��=}�i��s5P��6L�8:2µL���B�cR]+`Rj��5�����D|�m��|ĹYF,%�`/�n���.N����j����#~�Ït����j����Q��P���2  @�.�����5����bv
	郍�;4�������¦t"}���|�0xX�8;'���Tk�>*�?�9^�˚���Wv!�,^���r�O^\)�·�pB����R���xyye�5TT>|������`x�T,�A[|��"~���+�:88 �&R��HPP��q��w+ ��PȯN�\�r�x�W�{������˭**-龫/8�wl��0�T���Nc������{��> �斖�YY�G(Mwwʘù�֬�����+<|��m^��	0?5� z 4(((F��0��2� ZW(!��AZݲI/_��  С�p����T�|�j4ONm-X��Җg�>�	~���Rmk�4�*k��b�W:E3<��1�l������<����o�Ù����˵��F:��@���������u0�ɤG�oO��N�'&&�E6�#D�R�������|"[��'�hьA�S�R�t�V�*�	.���謯ܤ^4���N[���؞iG���a�~(ƅ��s�n�����)Վ�낪��u��	������W���V���!�[>��L�������ܐ|��+!��ɩ)H�D��l�ܬ,�P2�1�wJ�_'��`1�j�	�x]n���N��&9�q���f.bv+�+���J{���5μ���S*��0�ȅ3��ӻƣ[5{o�9"9'8���WwY���B�%H�LSCC���<��3�+4>��Lօ �������1wr�A�:�Y��pk���?E��M��f�=����1HU�d9y�����n�S�߿�=�&f�U 8~YP�Ch#����H
}F�}�x�2֔��	D�6���|"�{)��o�����o�
���<���F0�еsx�5�3�w�xl���n!t��1�萸��CoŇ���څ���K|^5�
l��AQvvZ�N������'<gJ-iY=��;� ��yKO#���[�Y8���RfK����'þ���%]�w�mf��o�y����쑑�3'8�H��^���g7|�͙���4��(5�Q#�^���yy�G�:��d:��{�	�*E0�6��{�K0v�#sw�_�w��;/�d�z��`"��Ar�V�h$3m~�
SN��a�xG�-��uHIz�'s݂��2zO��^Hɇe6� ��3�c�{H8{~�Y�B��|D! �*gP�<F�5��{_j���8�@����"P2A6�bֹ�,��5�b�|iVś��[pB��Qr�'�27���7*��uT4{O
�D�x���ɕ��6�'�c��� ���g��qr��C+�(OH��mʎY���&4���%M>����d��j�WiE���K
�.S�7��PL���8��ۇ��[�gZ��n��1�����·wh��:��������L�P��o�3��� �ܫ����;�b�;�Mי���n����O3�������&��N�y�)���}��^l:Q�W��$Z+/D� ���ޤ 9�ΪO���}xi��ۺߢ�������h�x�}�RF�/��9>�[��?�4��C=�S�p���4�-��܆pX���n��/���DŦ�:Ăg���� zB�����TXJBHq�_@V�*Z��[Zyj�3E��vDw�Ŧ��G �z�r{j`�g��-��%�-���\W�w&���Ҁ�8���Cwg�#B�3�Y~�)�r��|f?�����O˴)�������{� ��P�T�Ҕ�m�ȡbO�X�z/R�b��c��{ͤ?�Z�h4����>���}}U`4�6W��j`�TU��;9>,=��� G/n��T���`�`�]Q�Ң�3�Z��4s����������������!����|�~�Ը�˂���{ISM-z�e����q{PH��ȌR�`����g����PN0�L(�~jo_1-��u�ζ��;~GC��#!Ε;7iJG2J��ˑN&�Saa�3�]�c�w������82��BK����Oթ����9���h��p���.�l[7�>���x�ծ��55Hq���+ �iH�5 yBK^�up���g���FZZ�P�"Y��E�'l5�j%a��c�����fݿ��Pڎ��"}'1$֢ݺE������72�����n�ś9�>�>�i8��B���
�e�"@	�hޮ�c�vT�k*���u��,߇�f��L�$�1�s�!�����=j�[�L^�7V�Q�J ����É|�Sk���g�����6:��(ࣷ�{�����g|�����\ /���K;��AK�zz�9#,�& ��.g��Чb^�$,թ�%e��I'�.��ׯq�0� )���s�K	dx]�U��폊)�D���R�;��h��^^��~��HG�F������V�X$ �ɏBUD7�A	F��R�	>@�x6}�����z���m�N\
|�ZWp"ɡ���I��E3)rH���W��g|����!� 9?�6������cc�%i��Hȳ���X��>�ՅG��]�����\Qy�z$W�Sr���#b�Y��V�L}��B����U�=$N�/K#�(I�n�mC����>$���k����Sy����ݫ
����--/�]2Ժ;� uK�������@|��zRq9MM5LJ�v�I�{oM��C�ZQY��VId��rv3�� �U�.G����qn����,n���C1���抉$���W�N�:hoA*��47OC7ůj֭�5�E�����'_�ЕRv��)�#X���-W��p�꺦l��[
��/%�`�ia#ԣQ{����Wu�e��J�p��MRR��!��'��V7m��CR3�G\����@X���[�>���O���SW`U��t�<�xX���tX�+,���MHD96�GŰ�[�� Ń'�L�����J�nd�D�ýX�H/\�
�~+�~[]�s�[���j�B~F�OD�逸��؊�ȓ?�lY�ᲃq成�=Qmy�/s�����55N:)w�B��yvW͌��z�vc�4Q�H��#iI'��5A�Z�W�6��{��L�.��U@�+'�ٛ���k�Fw��+�T�(@	b���9#T��f�/M�j{��*Z���������,=��ګI��P=���H�*���Z���f˓��^��_t�F��с�d��?�k~�h�<)ɋ�ia9,y�%S֮������n�m���u>��zӆ��R8Ru���1��3�)&d�~���Ց�[y���6�����{.3�je�V�}�|��@ ���k�B�5�r_��ӧ�HU���谸�S�7ɒ*����A��|M���k_:%"%�A~��6���ǈ��V��~[��N�&��Z��KIY.ˋ�k�'��Y�o���wp�@��ېB��x�8[_��q� �S���2���.�4����2w�p�f1��E�?KȪ��\ֲ�WS]��J��)WO�^oH��W����o'��V×��h�x ��lû�-{�{��}^��5�$�6�V����-|��q�(C�#gs"e����o�ΕΫ���s>���Eތ����%��d�G8<sg1����ߺs��b��e;C�����g�m~�j��ϬpR���4��<Djb�l�)6.n�~') ���]�-�G�����9�#XU�ü� �� %�����*��Z�\P�
���%�r�K����z@�v.h�`YYb�5�W�:sM���8[uL���"�#��B�V��}�!"�����?��������N���NM��a�Z�c�bM��]/��STbr�g-�2Q�:�{_m[��s+�s���+�4n"-uDq~�4�E�7��Tv�[[�ɼ�|)����1S�u�V�B�74��N�h���v���Y|`���q�u��[��"��᪓)��	S��0�{?��m��r��T#Z:�]��z�V%�����%^��}:�^��l�g�[ib\�D�֞Z���3���U!��.	6m�����Yݔ����ann^x��r�*����$��%���J�C�q,�E��FJ���BVn�S!�u��M(�FN8��o��[��9��؞H�#��O�w��Kr��٠�(���������R���((\	� ;5�R��3f!�JW^�ܸ�-�wj��-�g0+Gj�٪��ܠ<��`L�=�����A�D�%R3Ud��贺��)����@�3&�;��_��]>[�\?q�r�~�~�":Q��&J��A����t��=�q���jW){�zM�]���#:{��ʩ�!C�"��",�L%�w{{�f�k����l;@��F�����S9zH�h�uCBBx\�@\赨�����E[��\�9�[4�<x� ��{C�t!C����}��P;M�'֭�  3x���?;CtPf�ȟǓ^�(��7�w��W�|���w��t%�c��Q0��U��Ǵn���+�@�ͭ�/��;��}h�c&��v>��s!���4��M�s��	G)�e���iJ���ŵ�Z���1[C��F�K$g���.�1k�wx4��:h�`�=�m��ϳ���������U*c5��E8�4�w0�~�Q�L�a¸����� ?�b�t��a��j )��H��y3����
�-OʭƵ�,�EY�rɗ�
w�Z��5J�O�I�]�W4(m��ߺ=k��d8Fj�f����-*(Pn_�D'3=� K���4�I���u�\�����ESO���:@J�g�A�����:r�r��S��j�\�� 1�#�]Si�}���rߏӿe��K�y�t~����omu��^o���/��j��pPm�H��g����J�82�ͫ(̜�۫	[��)?5�l����%�Yk%g��j����ݴ|��{p";�O����f��8[gТ�0'G�]mE����qtf�t}�8����J��xxx��Uuu� �_��������ԧj��zL�|/2���}���>�&x5��sZ�W�B�g�}����O�EY=t�J6#���s�n���V�|�CF!�����Hq���.@*n�c�*��	ZliY7Y{�_H��|�x�ޔ�ib�eV��bI��N��M93#�4� �� _�1����mw�ɇ��._��#,|����m5!P�㘸�u�񜝝c�A�\Z\챐���K�11�tn�_�@��Q�!Y?o�����N�z����bS��6�[�ko��+��+���k�����Ma|�������R��O=�"��v��b��t�;�.,򮟚}�/1O��i�~zg$(���
Y�pG;XR�=����zT�}��Znn{SJ�=��q=PM9��!��'���	S�x�5c_�p�B|ݺ��
*���v=&������H�"yϨ��Fad!buX�{wb[��������@����?_0l��*����/Ūԉ9�?�ȋ�����H����o���Y*�*ٹ#���d��K��W�eo%t�{��$f�\���>��&+'l�<����ˬ�f`���q��/zc��G�cr��( �ⳟ.��Yg�-�&�ȩ��x5+Ñ����_i��)0���̾T'��%��'�[F���\�|��R�j�M���9��kcE����:����8�W/�����#�F��f�llj*=�Go.go��u#�q��qO=Pj��˻m~��r99��&�&�9=M���% "��vkE+N;o�|�=�ƴ��ѷ~s�uI���8�Ie��v. ���D�d��)�d��P������$�l��R���T��|�=��:���Z�^X�%���������{ID� W�����D���z����:����;Ϥ�v��zՊ�
�������n�Ր���������_pI��i����w(R0p+=]g����xJ��ԟ9�(�;g����Od#���{��d��W�H��t�=���"> �tʲ�_G=��r[myQ�]��[�����I��b>��N?q)~?������W�!��&���i}���7��p�w
cd�ǔ.U9���*X�B1�,�r�(�/{{PH�M���$m��*>d	�Pa�i���EU*�դԫI�S��:LW�,1����pÊY�0ӂ�o�o�D�6��>�S�@�GSsq�r��O� �͍'��H��W�͠^e��}&1�fP��ROdr�.�?��3�Ҁ:��Qq^�z��\q�S��r3o���25�c�wT�M$s����-�I�����M��v1��l��]�fKL.�֬K�e��O�A�d�����8�w` :������p�y4�������[��]�e�oO6�Y�҃fo�|�+��~�����/�2�r�(5TF[_|P��h��oб���� ��Qx�H1߃��N�>kk�DD�z/{7��Z[�K�+�m����� ��ׇ�6��"��p��
}ZyY��
)[�B�`�;���9�~���d���2��D8_�<Q=�bX��O�0��X�9��o?q} � z��!&�L��O�	U.@	�g��z�p	��,˙D���|7�n�'@��oD��x�x�ߝ�ŉ�ɯ�g�m��|�q�����g�����{;���U����8�jF	�"���1��U
�V���:Y'�pg�'�D�~U���=m~��}]�SȧUp��n�V�����¬��������۷H���]$�e�ꫝq���"L�=J��Jt�D��oD� �UL�{���h ܇�6��R�MW�5���o��y�*I;Y�Ք������N;���������mJp9>����`����<�
��3�v!�0n�n�1/��'��n�?̽wTT˶=�r�k��((�@R$K��Ar��AA���dԣ�( 9#H�"9�"Z�d����n~U��w����c����Uk�5�\k�]���x�A��F0?���B?��p�>%!���l�TE׈�l�^��w��*�!v��/�6��@q�x��}]xw-��Z��wD�X��^�#�$��CO]ͮx�H|⹚�_�_�N��G\�9K=�2�Cɦ�;s/�6��ͅ/�T��:�,ѷ�@K8&:w��yI�K�G��Sƣe	LS33e�F@(e����Xo�D��aUS�/����y�Ƈ��>ݍ�vA��?ٳ83??�� �Bl��+m�'��(v>�cYI'�>넫��:���������o` n���m�[/�T��v�\��:����Ļ}�W��d?��J!+����,Z�ru���͒��tW��N0D<̱,���M����������u2?�jxs��*������/��l3��O�b�e��(P��� J�jLM`��S%f�����:�P�^����ss+��iQ�� )�]���}2>z��9
6#y6�d����+��rkuOx���.6�\,ML����%#|�������
�����率cF�l�f���5��?��?�@���L�@.�X�@�y�ϕ�E��X�R����N�����Em��H�2ӹ�Wh�����E�N�P�����q������.{Q��1����̹'@��DK�����+��P�%���;]9���m��h����8�m��ҋ���n�i)-u�Y ��#t�G�<��e�)_֋�ݹψ��_����U���o��>��i^�ւ�m\��[���y�"�r�bq9�gMS���6�e_���kfq�,�ZMEW7��������)P6�e�����,�)SC��%�Ǔ�M��V*��P�;e7�[���!wsn:������ Ǘs�"g�/F�pk�GN����Ѱ��܎�:w���k����K'�*����pD��<��s2a�;�\�4�ǌ^�{W%'�΢]ԸjC��e5����6�4M���:4����^߄������O�|ic�RK��
�ԩ��\v^6���JkJ9�|yp%�X�3!;�p����M"���2P��I�	���j���7a��}EEG�����{�d}�#-2��0F�P-��סɮ����o�Ē�i���ܻ f8* ����l�TW�v�-g=����d�h7�Ժd�uG�����)Ij�/�1�^�>���j0,9o�ol�b�������%$��� {���T߀�.�=� G���A8�Q�%>�C��z�0����vVU����s�t��IU?�^��cf@a�I�bw�Yh<�l���,���#mˢ?v��7M&��w�R�.ix��J
nR��(������Y��*v!bJ����� �Žk�Ϋ(����ɮ���3Wڽ?�)��P��В�t��/\5���m� �M_��8E��u�1�
HZ�'{k�r��1Z6���:	Ӓ���9���H��$�p ����`��ͅ~�P�kxO�2�7p[�y�9m���FZMx�w? ��� ��fX�$M����则�%n=$�ifu��<@���Y�It������S'��' �̞,��u���"~���Q����M��@�uC��d��%Jȭ(F���@K��/ϰ��" �R��h2Y����=bt��i|>Q�?Rb_)\��q�HX�e}��V�9��=�<|W8jK�WJFO��=���wY���󻒽ڈՊԸۼ�_�� .��G��%�:
��BPb�1��=O�Qb>I��^_�$a�����B�*�%��5�P���� ;�\��-��m��l���L�g�m�yl�������|�`���j��w�J^NAa
����]Y�?.����\Jg�v_,�4R�Tz���eY4��p_��$�E+�~0ӕS͠9����лsYEL�91�`|n`��6h���a��w�a�+��Z�!c�a�5���ko-�.+�8�C%P9�Y-l��[]F��O�I^{���oE��=���=��#.����M�
6`�>~�����#J�N�_R�yY7n���;��2~���'K3��qN��*u������)G�4�^���_7��z���I��iX2�L��败�6󰓛z���P|�?��=��Ih�s�k�-�3I$�rt��ٹ3�!fbWt��+�@QX������W�
klL������4�����k$�.���T@����5�%�󿠷%��:��9y��O������Y��T������YRT�w�Ц&� A�������nf��Ѵ9*W���>|a`+ۙ���^�p�w������3�?�� �dV'�|Da�В�yN�4ũ��^���7�	�#h�33i�߾�
����o���_�˺/!��ٙ8�0?�,Mw���MN��{���7�B��f��p|���s�(��C���v�$]S��폯���J���+�h�}=�%c=7 �j�;r%�A�N-!+���p���uⱚuC�]s�!i�T���d��ﴪ�HR�×o?iK=Q:�DԖ&/o�D@����l��\�2]�X �'7(�ϱw�_?DOFi�&(>U�ϟ%�5ʗ�l��ګ�,@X<�Պ����j#�hy�w�O>�}8��C��V%���<�p!&fT��fc��-)��d|�� '"������tUDk�7k��G����E!�MP��N2HX]]]xC����P�~}:44�Ɋ��_9�2|�f��M���B.4��l�_�$,�72����Б����Z�Ί����8>{Y�u�
�������8K+����7\� � ,,V�;�y:���^gC���$����a�׾m����O /������Ve���_o��7���}����.���ٳ&������j��/nݺoUT�[DF�^�SQ]=�_@ �+E�[5��0 ��ֲ�3�]-B�Y�fX��@(l2��×�̯$�����_�̨07*��y�g���G�V�\����C����k�'){�>3�-@%-�f��W���7v���$���{��{�y#�51��a����� qS����|ޏ<��D�b@���%�g@Ut篻Tj��� ��KYk����Q55M?}�̤���4n��5���˵�/#h4�$�d3���v#���9e����̛�Y�~��v����j�+�� �͇��y,\�����Z��q�Vgg�6J�(֍�~���J��OJ��=�]��O���]�_�y�V�߶IXX�9Nvw��,�u5��?�d����)G ��[�����YwJ*��89���a������gώONL01���O���^�Z=���鱍����j}�ؾL^|��ӗ�i>�T�V�	&]	��_���%�̌8-#��P�0�{��&yy�����.{�ؗ���%W��b����v��Qa���gy�$tt��'jS����N�f:����.���?(������/����3δ� �g�u'p���� ��D|�y��_�����
h����R�W:l������E^3̋���#�s/�[�>��#���0�;��AeZc��R�֞��ӎ;��yP#lV����%UgX��Ek�t�H��y��iǙ!>C~��n���B�6${m�LF�,��R���]��j2w��,*3�6�S�GmZ�LI�yN�+���#�a��Q�@�r�x8��L�@���E����ٷ���a�pྖI%�p۔+�]`�cY�?7��ͯ��;�ę7"�iߘ"W��xO,�|t}�X�!��=��ä�@��k{D�mS�=�ϯVj��?���􃅦�i=K%�=�y_��	m���xVN��S�D=��k��oz`�Z{|T�l@@�٨�{��֩õ��Y�.UѝS����S*.�Ʊ
-������H;����O�j��_��U�.nx
3h�0�$�ŗ:�?��sw#������v�����5��6��EI7�� �1>K�����N��=>N�mf�JBs����6P���CC>����g�Z�s:���5��{�d����ș�S7����k�Hw�E��)L�������������
��㧆KSt���\���F���{��9=�"���}P� �V��~ġ��:�I+5�a�t���p�~�
Bܾ�)��5��a�Jfq�H�y����6.�&tͶ��Z�!L��~cᑪ��yw�d��A�o�(����z@��rI�CkI�J��& %'0nX�=	�;dx�*��wdj�/礇�VrS2j�?I�F�[�T�Q5�Q��}w�>�1��U�͹G�0�����JUQ�y��ǮX.��9;[֒��:�?�X᜿bk�E7���f��.�y�Z-��b�{/�<��S9]~�2����U����?{YԻg_�p�X]�֘���z�?�m�ֺ_`�^��s��SY 6�±��]�]v���qR��o< y�H�".����C`7�2xL=�0}G�Y����lN!�x��믤e�$�����!�^����������~7%����"�9���fJ�'e�bw����9]�ޣ�O,��]��Umc;����$u��L՟�+���ā�68޴��`�H��)>!ԡK�v�◦@0JSu{Q	�{���J�;�}�;�P�����ÙQᵊ�z�iXt��՝�ϝ��)o���0�>�!񘆆�������Z�z�h�<G/�uu�Bf�cL��>�,i�\K�ұ���'��6��ǖ�-�4�?���lZ�"^�\"��W�1p�A�y��T�,������W&`� �\Y�l��$	FjA Wa�U�p�3��L�|�}я��^�R�?+ş��i��7l��B�������d��4��mw<��{ש��s�ب����J�(�����f������v<�R֖�p����F�bt�v[�ZӴ�uWBG�f���@'.�n��y���N�|���?`���wс��ן����D[a�co�֑��|�������!w3*�O��Aչ�D;����[�3����#G�%fu���^��"�rA����ש�;ү�^��}���D^/MYvo�O�l�й�n��9if9��^�ſ�t��YP7�Qy|ڎ�VZ׎E6��㠻Jj�\j�`��J6Ze2���F
�x�N��-�	�·�>�\����Oa�eY|��B���N�]��J�Y��4�{C��h� ��d�A�e��v��O}՘�����A#O�D���w.s�o癚b�f^�/���9襀]�#�5g�@�H�h��d7��E}�/�DF�#}&Ks��񭭥+mE�w�Mؕ��`�O��rS����1�Ԥ{?���w˔Fl�%���#�i�e� ���Zl�����j�^'{��P2B <o
���@N�������É*��ᨈ�����J��Ph���[��"�Y�� �.ሥf��3¹��.����-rF)x.v���5���`e�?P���n�mdP�==�E��w �6�i��ʧl/���"#8LO�5��6�`E�7�0ۙ!d:�.��^�G#G���=Gq�~��e�
�X귳��R���ՊS�sf�4�,�iӍТ�΋Y�?������Urv:o�彍�l_xR�_l��}[Ͷ@h}[Co�8�̴<Re-ycd�����@�o��ܘ�m�l�M乁����R��)�6���ђ4����h�˶OTa��F9���8YD�H�����D�I����_��n�kn�ٴ�pu�W��xLV	}�Hƽr`����nRNH�ވݶ4�
��ָ���oF�'��L��:��{y��×�9��G�G�+X�'��FM ��x�8m�#T=C�6z�a�2^3�M��B�lXi:U_�#g�
���/�
��df���x�9N�LȂ��<yk�2-�˦b����e��G����M#L�ם�5�Ʀ^jl^�KF���F��ˬ�W�G�S���su7s�%^H��ձ�D�8�|��	��kؓK�XEl��]˚�G��+��	K����K������Zݴ��"Z�d��Ɛ���Ψ8���oF�X4z芭��ܐ��(9{Û�B�}��qw4l��&���4�5o���Η��V���9:��m�|*]$$~)�����s�N"��g��'����<q(���Л�BC�&��{�M����-���[Xې�G
"���)�^,�前 ����7k=�u]��oR^*ɋ쌽�,ΌQ��dc]��\,x���d�@�}W��|��;���Tr�=$�.�v����u�EW�c���AH�9�(,D��?ux��.`�>'��Ǭ����#��2���Q9�[0Z��R��I�?<��8"�cOhPO�6���~�'�s�ɉ��m����'|��Cb1h���'>7����:����?h��p�(���vhH&Y{C]ϟI���]���΀���lL8 �-h�&P�7�DG��5/yvh��Ж���r!@�f���2�mQî~l���M�8��ߌ!�	2�	*z�������|��l���/u�[�ts0vM�r ��"�&���@��ܼ4��d6_q�P��d�@��B.�F� N�D���ק���Q�ݍ�����; q>���V��k�(���1C�~aE�QQz��q�ۗq���۩Ω^49��sS�c��� 椠�j-�b��[o��ʴ�m��g�\���l�q�K,d�ta.ɷv��B�@z��i�B��>�]LD�W��cM a˻�h �"JW��z|q4�g�?uN��Q���T��*)c!M��s��X��>]�6�!���+��Q�5Bv$t��C�pn2�&.=���záMƃ9�W�k���M���_[�_ۼИc�?%e_CdYȀ���'g�>��y�<*��n�7S++����S9��T�%T�����dܕ�[Gp�&��C%��t��]�:�G�&!@��Cܪ �"�>t�d!W�dk�%_�ۃv=���0.2�a!ӠF���|#M0�<�Ĝt��$�K�n��2��|c�G[(�6�';�9�q�y5�,J�_�9�4y�`��!�&��A�3l��Vuz��:d�T���.c���͗�������+���'9�|Ӫ�����M{eeU�j>|8�4	��['�0���_����oƅ�V�&U����M��8��WcH��o�@��G����\ �7�n.��V
��|�NEF?FL^6��K��k�%	�H�(�
�;P��ܞ[0���e^D�)h����w����A�R�8����a��m�*���j��g}b�qϸi)A?گ����ţ_M0�������p�c髙�U:�����$lg���.MC��^D8���1�2Ѻ�I�f�]�UR�1[]YqG�I��u�%8��Y��Ռ��o͏�vƐ�1����tw0��
ht �_�����Ls<JV��u����ZM\�;B�a4�Rҁ!X7���T�<���I�����~� 7'U&T1�8��1�73��Sl��u�N�^�w%���kuUM��=v�K�yh�h�p��Ά��?��Mۄ����X:��n�6�[�156�ɕY�"|��Q88�U��$&il�rӷۢ�5��H*ሂ�F�Hnˑ��\�l����2��Tg�?3��K��ܚr*��LR��2G�*ߞntX(j�7�~�w��}\���X���-;Y������`��"c<tR�3�Wf��֢s�	V8��u��_��e��4��i@O`��&�]]:n�i���4W/z��\��</߸����R��(�߱�lx�T��j�aƢ	�~e�LȍO%���{u?u�I���]Ɩ�c������ߔ������ݜ��(C	'��uw��{��VÝ�q�ӞP��!=��oq�cP�zS�1�,9ǲ�\����f&���~ݞ	t�k9�FJ�0��b}�%�4#��:|�V���E1 UZ��>�k��MT�V��j�AR��g���i��|��P��5ť�z

,�WL���> 5�̗?�߬R�p�=��K:3}fxq ����Ú�.
&s���?�iS��6.�t�*J�=�p�������b�J0�ve���H N^�P�7�;
�K3��c
?��ȩ�2H������-���a�X��g��?w�͇���w��������(ݺ�;�l��53��r�����y����t�2�h�P�0_C���P8���L��*A6�/�f�F�T�Wo΀)u+1fp8NL\�V�G�9i) ����v\�v4�- ��W���0���(��d�*]"w����]Z�5���9��czR��-v�rwuj�C5S޼����1Y]v�rsz�d�����8(:�q���|��WJ1�7�:�T啿�[�{�o��44�,�� �#p�IFO�Q�E�dճ�r����<[��B��d�	�30$����d�X��zL�9n�;��N,��_wT�����=��ob��o>�Y��2_6�6�ڼm��BV܋ ��f��m�s�����'�pB��Z����3�@V'!�M�-ڝ@B�b�^����0��/@a/e-�:��X��M"���S�92U��*~dlQpd�{�:�0���ej���u�|�c	���A&B��FSUG�P9zl��a�`G^���@Y�
8�؃�!(�}r��3�&��I͍���zs5c6�ɦ3�������Z���g��Jq��P���y���2?�i���/C�k�+�K''�1G|U�FoLR@�s=MFE��9����Ӝ�q�)^6�@��.���C��-��3���-lq3���E"��<;���+F>��@���V\��Y��0����p��7�V�lj�qwz8��/��n�_��m�za���6 ��D�,17@���7��}|�k$�5��g'�o'(���YQV.�5y$,�l��bu�k�].�x�|Os�A�Q�K8����A��Ns�{�Kq ֦@P�t��4�d�����^�����r�Z��'�3�'ӏ�
<Q<��E1�i
W��E� ����3�����5�4����� ��� �
�g_�t(��3��f�m�����a�^��u����c�:�l�=��߽�k�x��w�pƓh�f����@��v撕:^2��q�!Ɛ��2��a!µ��yO"����W!)����'��s�Ut�����ț��g��0���;�|EA��Eoy��if��hq��3��tk�0�����1��u8�(wi�C -��<��c���A��Y z�0�#�cӍ3��>���t�L�F���?�:��U�Ze�,%\�Ԏ�͑.�H�~����f�??k>%���_��	��,���K��i�w���@��!e�Ќ{��J�_�������mRٰ��#���.
$��X����i�x����E�>�Ӿ��x�H�+����0����BR������
S�@�����'� O���+TQ��Ø8��T7�<&� YAmB���y�*�����������Ic�\ppc��r�'`�D=��Ӟ���y2���Ց��g48�����K�*�9ybA �+��b���/��!��<k�|�պ����&��%p�|϶�Y��w�j[6=O�\r^��]��#i
�+���O�ۡ���?Ì6b��d(S�i�..l���)���}4(��P`!31�H�c1��y�)\`DL�L�����LKUa�H��yC��3^��o�F������c�D7� `�����6�r6S��]n?8Q�P#��I;ľ$�/��:d�˗�UN+1�N����X�:Bg�v�����msV���O���m��v$�<a�>9�[����8�I� m���=��	DSV�]3P��9�uD�4�(�����Px4n���5��w~˯8KES���e�1��T��O�n�9�p����:RtS�@����w�i�w�7���Fv��� �u��|=N�ٿ�Ƀ�=j�E$)�7�8uw�&���e���q�)e�@,$��V�n��͓�!ǾM��G��t�F��\�pE���_���b��d9��uZ�0�>9��<�WX]�?�K�D{W��VW�v�Z�`����)�Nf�®��7�{��˜���{�3jp��5���`����z)I����T<�qf�
��w��|�mw�<Fk@�7, ��îl�O�6\8n%��d`Ny�j�� RT�P!�WR㻦�o����K8ȭ}�	��\�uS�_�����Gm���n&���T^K(`�l�c��_S������d6b��F�n�@F~R�50�vW��AB
ԍ���ۂq��ɷX�o���Ft�U�w"?�or�5��:��׷`~� �`��o��6��&I\�S�A�����0!����ݞ��0geh�pT��w@]qp�	��8�S�*�:��g����1�u����&�JH^<���_j	�ѣ\��_�	a���t_ ���"����n��L�ڊ�rB�� �É�3GB�%@3ϸ��8l�x�{��@�=��F��9�
9�b�����@�-�s5?�<J�c���!Q�f ��i�,�2�E��{k:Ku2扎2�m�/&OI�,u�2�n�!��
g��y�>n��π(�h��e��_0i���G!���uk��R���[����N�]�8T��緟�QA@"7��ư��'�{�\ެM3�X���B.]��%`��A�����Op'ջ��8{��\��h���Yao�t�aW����m��WYw����]	��%*���/\����f���`"��,�aY��,wnm�]:��g�ʷ��q1��΄AeF�o��|�:�pg>�t�[�3I����MX���ʓ�p�x��YS��kL��_�kPf�x�<3˜kKKe���y�8��:�P�n��|8X$=-8ʬL���*��A^����\�{�'p#�
��J%��Mse�v�����̰��I�Ɠ���F��ڪiH�Y������&���e�*�v�x�����l�D�q������/Y~xw�m����plv:sjz���$rx�����d�'�gLh�8pcǃ5���㔛}N.��q��q��a�fX|{�0���mt�a�H}�Ӵo�r�Y�r׎�����X�)]��8An4�D�����n�����⬫暟���Ȋ����W�4^�O\rLNV(9�#w��Lݾ$̣a�!��!��E����D�����Qh��4Ç�&�x�Vxsh��Y��e��/`Ws�"1��aNW�0 ̤0Ͷ���8�?	
�tq~9�VR11����r��>Y����m~-�I��<�z����_�k��{�k�Gpb\���'����c��?~LH�9 1'�55�IKTw7��F�z)��~�>������Ж�=�Ҿ���ny,Gf��[�(��n��_��� ��T�� ��&�+,�Y�,�c��j����r|3w��x>�j�������H��q ���Y�
��MA�7C���:::�Z9����޵WC p����`�[��i._(G�vG����7�wG�농�ĎJ��`����������l�2�*��zX,XXX\��GB�X˘Dv�EvE<�t�'���%;�b1��"��YFg$"N����ب��y���W���.yf��?������1O~��aֻ8yx���9HD�l���_�?sY�k��OlO�<Z��a�U[�>�SQCbbbҸ�Y�l��\�s��a۟��0�Gke��2��h�׏s����,s���@tΦD���z��z��E産�t���#.�E���� �,ݿ���p��X���W��,ⶐװJ�B�3�W6;;{|����m��C�~ZZZ�L�Rb��;l�滻���
�����o��X$+ݴv�\��މ��{����@�%赛�����}��j��ՀK�ǖ��Ѓ�q�9%�3o>g�U��L�Vϒ��mW��O��cH�6����ډ�u���.3	>w�j(^k���s���<����9����QV~Bbs`���#�}�i�����=$�Օ��ڹ#�� �v�~���v[s5hD�������x�l|���P�ӧO�۵B���������57?�'I�f(~�>\'H�cN����}$>ߢ����Nd9XT:E����5�c�:J�BW�<9�����م_SܹM��q�����FFI�/� ]�c�G�1��K�:����L����B��{bv�#ㄸ]�%t;� �P%㫳
^��a�p�m�2���s�Ή��^�vi��[���)T�epp$l>��r��+[��s�v���4+�1��V��1�M�iZ����pq����鮮.N��<�Ł��x�i��$���2>i������ ��q������f-�I��r�����M����Qt娌��~!4�}����Q���e�]��}����f�`be�H!遲���ߌ��S�m��_��.�ϑ��|�#;�K�l _��5�jY_e���E0,$Bx-��u��\q�=�Nl�?� x��B����l�������W�Y���I���JK�L�Go�n�VŴ�8��L�j#Fw�U]x�)I�ʭKG҄��u�t�^s�t�jhnRyy�����ɝ��U� ۟��L?#�h֑(�_bkHAI	�����:T]/23�,c��H�ɕ�B��V�'E�k����Xcz�'�����E�ۉ���=���4��E���9�����򠠠 �wT�uT����c��{'7�swvgN�:����Şb�K�9�;}ee�x��/_��k�F�a��8��e����s�CwX�a����������;��$���
��)�Άl��aέ�pt4n���:%z���|�U]N��w��גۨ��Qv\��2i1T�G�Vjw����r��yb�JɁ�^T��XM^ja!w4�����Z�G}>R80dt�&�ݭP���N����:�X@Spc��$^w����ӘGz��c���b�Gph�L��t��;�[$���>fN}-�ăik�ͺ��"P[w�W��d���`�F���i�i��V4�o��w��� TMMM�~�V,������3��X�rkR�vW�s'ܫt��/��Y�*�Tnh
	�q�TQ:�����P�3�מp�Q�$AC�[%�#bâ]4�9'bm|�
�UH�Whis��(y,��RN��3�Y�J'�طq���=������f^�dp��Dm�HjU�����#�$�@T|Z���y,�og"x�#�ӡwd��k��}����)�I�EN3@m����̜��Z�[�/)�J����q�,��Xa{��
������ҍ^���M�/ȧd�w��v�����x�������Nw�p�]� �f^��Ǻp[y�C�xl�p�OTtql��A�����b8S���K�z��K��|��#���i�����^�X$	��+���A�ߝ'Hм���W��{+�*���1�^<�\�(�Ъ���a^�͏_���=37	������Y��OB��嵫P�*����h�x
Ҽ<�d�^��^}V��ӷ�A8,22R�e�d���|d�j��aܵ�h~nnu%�Kp5�)?��@IQ�,>�`d��9��}�.��8�� �e	/�S6����ݳ7<h]-D���@^W��sqA���m�°T�r�m�855U�Ό|;7�!��ڦ�p;�ջ�pE?�ԋs@ڴ@v��,�e��i4Fܚ�^��Z�k��՘M"�R�hUnߣ��c���g|$獭���������|t�x�t	��t�*�M��]�5�����i����*~Gǔog��g�d�EM̱g�  �v�ݪ���ٌ�ʍhW{Bυ���GUl)���@���/|�'�ːe���:^�����o��c`b0�LCƦ��@�@����c��cB�5v\k�H\����$e��M-Q�J=��	=u�p��"k�"ʍ�G������4O�����5у�lJ�c�v�m�f܎�݁�m�#���uWt{� ��������s271���pb)))`b������R� ��M9��W&���������l8>�b� "�@��M��n�6�&�]Kb�`l�N�oۄ1�Ekȍ�^����C���"�Q��^��Ғ��i�X��n`�b/t��0o�R��?n&Ђ��Н�{�_@2�Jr#���ݷo��|�������ɵ_nɄ����g�Of=��S��˴X1�U�ck�C�Q1\�<e�_;���^�5F��>*?;/�$��Jl�]-[+.�Yj�������{���+TO_&xƈ�~i��0�b�YdMdz.3��F��q����} X~G�)�'Lt "�bW��E��ҟ�P�&wpp0���]���-��%�����hN ]N�A^Hv[�ܩ�z�P��h�%@�����OT��+�BE��2_�a���(Q*Q;��;a�I�`���v;O.�gR�kC�x#�2Q���K�~2*�5����^r�Z,���;p��D�8u���� �M��>O������z#̵���� ��T��.�%�����>�G�5\`G}�.��"���[��0d��3k�1������,�\C��r4V3++V�'����h����I,_�\�0�����Z�ͬ��_	�Fjt���SJ��O�=L�X����_V�]Y��%���EO�aǞ6Ԛ�ǣ�\*s�d,�����f)��-��×h�,@L�ХE/�#����8;��uP�$Q�-�Fq�lnZ��������W���RT����B�MC��6�**I�?��ZXV0K^"���<;Q�(y�fS�i�Z}�D*�ʠhyJ��?|���B�
������ ��E/!iH��N=����)��^R�T��,;�H9Ȝ�i�_C��{���J��f�����#���'����Tם��!ͤ�a��C1ϝ��;{=�7\�PX@��}w�~��z�xd��c���n���.�k|�sKH�V�%�p�@LM
|OZ��Q~	`��0m��լ�87V�|5���t"�;���G��R{Ǡ��oH��	��եu��l5�J�bn�M�1��2ۘ�w?�J��ݏ�>�0�Q�^�%�w��X���ݷ�0�?���1**J�43�
.lU�XӦSl�c���-�SAج�m4�}¨�f	a�HN����|��Fc* ��|�.A()+�XJg3����Ks��7UZ�m�.b��2?���:����XXX�;��q^9E�.v��ʣ
`���!Lllȝ+벧Qt�S����#w7����?�@]��z�'���B?��=�!��,!�	>Mש����齈�(c_<����
E��ýG�n^�_hXzCt�������̷�8q��1b�Dי�'����?X�[����a���=�m7V���N�C�rss��p��B';i�G�Z�Q�L���U��^_�cV �|ϸ]C��wj�v��G�H�!�7Vr�F�E�G��5��]����7�E(�{��� �Σӟ�n�� ��8����yN��W�V��������k��)�l*�ţ��eL��=d�4,������N6�D��\�ӈ���u ��ƭ�̈O�?��ၭ-��k��jzs�\�Ǻ���M��-���6��k� `�.0T��s:z���@IQO�&44�7~�7�1��V��j�m��K�z����oݻ�i��r{o@�d O���^V{��}(&L�{3�x����G���� �6�*A���i��
�19Q<�ZC^�p�(S�ۂ��n-������|��R�f<�!A+'p��^�o�:���[@��=-v�h��u�H��F�&U��T=�N̽����,��4�IwI�d�
�^426��2�.�Z6i;=7^咽DM�Z�T2�dk�px�'�@�'�YK��T�"��5�˝,׮�:������D��
��?ϰ4#uNk�N�Dο~%�W'�P_�f0~4������P�Q�v"ĥK����}����� ���ڵ������#qmƤB�A������r��^�y?mP��*XU5S��?�P[y0� ���t�IL��9o<o��M�%��HP}c
5,���2��x:v����%P4��1���˯�Q�^;k/���3¿Vп�I���73=]��m~!�D�&�΢Jo�_�	sΉ4/�?ox"��^⍯P�jj �b#9^�X�v�JW��_��xK�s�am�K_)ƗS��^�w�L����֯m���[*2mbV�����p0�'(�~d�W��\�$�uШ�1~.P�}��ff�߳�S L��@X�_C�5�<�W\F�)?��������D[o)y��|'u4������n�k�*��(���c�ySʢjq�q�9�yl��ĳ�mU����/���hc�Ƿ݇�`ܢ$��^`����1qG�kׅo�^�E�h��@>�d�z��ݨ}���J�j����wr�<�>�#QMYlݫ�f�_��vR��.+�6yE�u2�25��I-Z�5���y������'�����u_��%W�]�N�,<���C�3���s��|k'��O�A;��+;���������μ�2�Z|uƫ��+z���8�`�����3{=�� �I8�a�[�>^ڎ8O���M����2�`R/�����9�I�HY�n1�\*@���vuZ�L(�E$:�`�x%�W�GS~/v�͜ ^vm�h��ƍ:)��L�\��O�[_��
L�}p�Yi���C0���
��k�ɧ�D-z�u:]���L��O
.�,����>���������8��(m���k ��1=}hBK�ӎY7o��f!�.[i��)�A������rt)���}�|����h nc��Y>|�]#{�x]o_�n����~� ���v�-x&�D���gԸJ�oϩ4y�as����N���ɠr�L����e�/=͎�	�oDv���ّ��k?��܇�5]�=
k�l	�Q�XX��]+�+�F����yȁ;����Н'�>LT遏(�0��TJ8aH���9� JBC��Q?���b{��+[�-�š���d[^5�f�s�?����b��9�܁#]���!On���nwǻ��9l����,o�.�>}w0��_���Ł��n5�C��ybv����,��F7���=<�9��}�뺝H�A�N���`4Uuu�jO̅�j㶨Ɓq��1�e�� Z�`F�}�Ҿ?lU���~w����'=f>w��2��x2�D�����B��
�l�m���#/|�O�w*�'!Ѳ�zd�6��J����o&��-���@#s�
�C{�n'�@N��S���i-�L���ȵ�M��}
��׼���(ľ��,��0�{���0 "�UD�D��̳dH�NTm[y�� Һ}$@�C�KG
'����n���i�.R`��`_R�zXM����8��������"�b|q��ദ��4� s����F�ڨ���A�mN7v�E����K�&J��ag侴�ueF���O�	Td^?�����/���>\���q��>�p�h���.�'�9=�����Q�omĖDN�֘�s1�8��P�J}r�s�v�����I�������L�c�����u�W�.iXy�1�+��M�0�Z5����c9�R�54�<e~�β�;�Ґ%�	W~zg��7�(�.Um���^l@lQ�8��'�t����/>���r_�~��Dӻ֛�V�͸7�i:����ً�2�ʦ�5��z���;�[e��,�U<��l#Ǘ�&j�E���Vz�R�1�Z�E�ͺH�q�}�b��p���T��'Hh��R������1�L����/~2S-[�A����ݽ�Nse��Q���+�'�6�^'(���з	xu�����9ר����n����F�'��T�i)Ǹ�	)ȩJ��!�޶��ab]eǭk>�`ڕ"njj:��g� ٽ7����<O�(�z��j�������>��HO2��7M�s,���,�	�I�}@��!�SIW��p�.�
M�q&b�nFù������&���~w��5l���)��`�c�M�S�o|��ds�R��u�~��	g]\��p���x����gU����J}��������	)lT���Ue��8HH�ֹ�X�W�������������}�N�6J_h���5�Ƶ�[�N��� tz�պ���PUU��ifn>�(�#E�\�'{BԹ���yG�~̫c��%�����С�4�O����2���$K�j�U�b�:$j���;�c-z����4�`qp�l�ݘ���ǾbR�>\��6H::;wV�455u\g�W���&��)���:�₯�A�!�OF#r��-܈\9��Rɬ��?ʾ:*��^P�c�@@�[���F��.��N��N�.�����;���{���}�}k�Z��{���~���9'����[>��K��R�
�7�R�{ɚ��pW�=�7kV����pe�����O1a4��yD"x�xY�ևih�'��b���-�C��� �Z���)��+~<9������N��6�c���3�o(���..��8�<.�诏9���j��?��H2�SST1;_b@E������y4���v�U��M=�QV��!�F1����V�����t\���=I�����(.�r�4���]���xiw�螟�%W��gH�?�~�;��ˉ#l���bY��H��
fm�=���t�~�X-������x�+Im����|�}�A���I36�F�y�`��
�J�Vܝ?�Չ$���yH�Eu�Ҁ��|����Z
>ĥ�	����Ӆ�#3��^�X�K�D�,!���WFqo�}zi�8^f���{��!L�Aco{F#��6@���=����a�DFu��m�n�9��XT�R�k����dE��?�D��<�T��X�=~���� �&>�r��L ��JB ������l*�8���]��~��Dk"~g[���w��8Ƚ�E�:�l��5~��68�#���C 9��䫴4㔯I��w~x�S�y�zF`o~i,���	}���	����'2f����}�py��΢#0�|��9r�맃0�x�]����(�s��)T�������
T@�{T�k�G���=�⧮�	�1�L��~��F���bki���s�����;ӹ�;--������y�MU�&&�N��K>�/�ͼF��`��bP]z�),n��1˦3�PL��������X����v��g�$ɝ ���K�v�oo+LQ��>�6����D>;��Q�W5��O�����Q���.C<N�%uKf�YG��I9l�_P�ݻ���Pb2�ǵU���NwjoW僕���nr�+V�{r
�b����q,��c�aRo\�_i�}�=IR��}򾡥�ݘ����e�ͳ�p�zʩP��׽t
�N�C��b~?11��q�tņ�Av�����D��`������I�f	n��B���(����49�!�����[���mQ�]ulz[iAH��s����mx�rh��h��Iw�U�9�0{8s�됖�n���X$|>��р׻�i�����V���$�-�h-w����lt78�B�	��{߳�qG�,BED;:��s��.P���߬��G����D��ݵ�v�s.\�GMș/D��azq!����-�ta�k��"�2�t��q�*/gs����yo8�Ӂ�Ũ$M��}'A\0��A�U��[�gjͱ��������oÁ빧_V󢃼ff6'�����U�ƣ��K�h�J۶��`d;��@v�1��q!b�h����xY��d1��;�y�[ M*�������x��L�8�2�GR�䎳�cx,���(���h���/u�� Y���H�k?a^U�� ]8Z	��Z�H��v��3�ǭ�
,��6�+�	.��dt:[%i��\�l=is �_��8:�32��V'�XQ���ӤN�tq7���sK����ċ�ۉ#@^^\d�w��A�?:qվo�256�+��h<^�'��<� ���ZA@z߸��0�v�a���b�Ӡ�[c���H
.HD��7��c��GաҜSxP
���L�/o���ޕ�����q����>ɼGR�ᴴ��U���/ͺ�OU&i��oog�cIR������[]����� ��������/�y���P�8���Rd�[��uk�?eg���a���h� +ڍ�	vW������ގ�9��d�β��fh�ֹ�]y�a�J<V���A'̩N	� )5�v��ao��ս�*u)A/\��5~�-�0(\?}�j�ύ�����P!7KH���4 �r��tooo��o���;K�� e D���?��B,�kd?g�ڈ�ѽ��-�+����Se�ZtKw�<��/��������@�@�մ�J;@N�/�Q��S��h��MCAR�l�  �*���9]�l�\��LCI�*􊖖�_�~�9�hۤ����]�6PN�Q��A�%����IR���g��x2	���X��/I���d���A�
呪�ת�P��(��
Y��~�ID>d��x����I$+I.x��*-��� z�U\��B-<;�������x1<���A$�@�)IŲ>�;E[��7U��G��΋qg�ʇ�\�*�����/��:���n����۪�s�9��X`Tm=�3db;EZ����hMSX�4/:�h�F5�J�Q5#� �_����^^���"��3C��*�8�SR��A[�1�k�Ӎ.-���CU�,$<[Kz~�s��Pr��&��sV��;5.�z��JG�uwu�7l�Y�^�����\O(o����hD'�P�Hb8Vl'm�b�m�<}��Ư�;/�ʜ(�k<PH��6Z璻z���7JN���?
X�O#��{��~���.�~����\�����oGNm�s"�B��8��Hnt0�R�gV�6�-�vB�����-�̫�8..��E�X��p�`����Fn �w�ޞ�KPq� /���E�����}�ţǫ�{�A��z�K�ޢ������C���80���8^����7� �8b�N�+e>�ď@�f��XB�GEK%�����`����C��W��k�o�6?M/j�]�ԡO)O��hL���t�R�����x�P�w��l�P�	�?!h��'���y;�LMM,=N&�?�3-��7���.mD�W�N��3$��Ƌ�{���p���j�-^R\�<�EY�|�6YM���eGǷ�l8�����D/P�LD����a5�<	��>�M�U���L-�D�n^�Ի�ܼ���A����

�y��{�K`�H�8`�L�3|j�C��K"V:��Ǿz���Z"ל��h����6Y+-eVF9+�üb�b����}����B���Zi�.�HIK�ԗ���f@�숞���5��a�j\?Z��ɩ׀��0pXo�s���[A�R�m�D��?��ҁ�K��3��Ӑi�T���'X�PQm�O�NW���(���pX�uGP�	U�;�#yJV;��Ў ҡ� ����Gs3@zy�� ���o���v�M&"2�� ;=�](�	����B��9��A�V���Ư����68*W\<�[u]|�Z��n���l�>$"��7ع>N%�8�X?����{�S]��;��w�;i�a_�FY8���ZYI�U{��/�OlxvA���Y����E�.�>�Sæ��X����A��M"�a��o&V���7	p����!��}j(T��ߞZ��K5��:k͡�\~���7
-8Q�d%���& �P�r!���K��O�����#;Dl�6��M�#!TƐ
�/�K��3 ��h{�f��v莟wq��<�t/t�D���l�����1c+��e)t��4L�>xLr �n�t4����:�.aY�oG�7�\��<���o�_�nOO�߄.������d����-	C5`�a����4��j$jΦ{�g	��*0�;e�yI=�BTH�wf�����޵�s l��Q�
�׾(8K�σ�S�$y�t�ϭAx���d����a�'ՠ'Q~\}����ka��~%zЎ6?ܡ���#.�$��g �@|2RE���#p�lY>d���[Ծȶ	�1X�r��W�ջ ȨC�[$S���;�SSfn�*xP�Pd� �|»"l�NAϫ��O��+����Tb�dS^��<,����~�=�à��à�@�[ݻ��?#{X�FU�s+���>����o��/�vi8L�c�2� 4���U�9jcT��&�Í&'�@u]�!ujE;(p���FaU��8���X�6 �k��C7�b5/�-&!7�~S�"l�����\#��7k�B����I���5�0ĩ�d>#����3-�dL���1�S<|�r�V�ͳt,��b~f�FM{غ�Vp1!���`W���7��Bg���w���R����-��x{L��/���`���fš]�5�k%�&���ˠ/)qh\�}�� �VCҜ�)���X �4	ؕ�}�޺�X;��T����_�ᯉ�����H�M��e��P���Ο4i>�ᨺj�	���s-��̓zL2.fW|Ff��˶���8��|g��A`M�� S^q�FY/ݥ���^�Y	�>���L+��%O���w�	�4v۾xsF����َ��HZh��6����A9h��?����w�P+���3�z�"����ݵA 9Z �E��p&�Q���f���#�u�j9�!��+����A��ܫ��<���� ��q~

$ҁ7E�l��%��fCn���A�̰/ �L%Ǡ,)�)�4��i���MH ����9�V_�\�x�9���. %8ںpa?��R�2�n�2�&p������g  ��x��I�� ���"w"֏�O]�Z��U�< �uJI�VN#B�8v�����������d5X"QTV�w�Lp�@'i�)�[�>|��`>cuh����ŵ��#'7�o𓗃�� |5)O��Ld�d�2 �/�Qs8� P�@P�d�p��a`�g����j��>I��^��W�.l���KYi�V�p���ǧ����b��$IMyz}a^^ޘ���h�hQ9�~��71��i��~oޘ��x�	,�������
�^����1B%=�4��'s6F�b�\� �bl���� ���>z�0�2LϐP9�1�-�Hb��P`<�;���,�w�Kp3P$ƅZM_��+#��,�^�������`D�t9�N��N:���������{��%6��N�d�&���AsXjt[�rԌ�&A�n�C����r�U80��F+� �q��猫�W«�'��J���B��[ �{���@Lu��������"�	���b��t��	����T�d%E�6 ���O_V��>M��7| c c�O��
2w���}��@�����jO������T�~!�Fc�U���kEܘ-��@�	ďd5��q�� 0��� ��>1qI��N�	���4��@e��V��%���``c\�������#���'88%;�@�AK���#�n4���.���f�~�����\:�5��iL�ڕ���I�
�������-�������Z���A	�f��V�'啛����� ��3S�~Aq 7-���~ e0H���5���*V�6ߣ��2��t�L��$�A���Rf�ƹH�O�nG&oe+-��'wf�:����{�.��)Y~�b�݃��>'k��������5����QLZIeN�*��Ta ���^n$���ട������Ӄ��i�M�u�њ��3�@���X�٧� � \��\�9�m �p��yW:M� �G�V+keƒB��[��J�^k��s����bj�Q��py%���i���gacի��POE��̠������r6�n���6�n���i:-E1�`왿me�	@�����	�\�� �*�i��o��,bV�$�ܩ��~�k�p����aF��L#��@���E��@n����T���`#���ģ��,�Z;L�O`@0�Ouڷ:㧛���
X�fq�_�R�Lu����dHQ a%=-�i�M�l29��'a�]��$gZr��P2�VZZ������>.* ?:s�N C�/h��ZM��8�Ef7,�������z�(�Q&d�c:��I�x�j�(Ꞿ�w�
�mh�����1��C��7�/4O����R����.�&&�wM��e
\g}�%6�CT��`"fm�^C-�����ۊ�K)X�yo���A�8k�� �8�E�PHKo%�ؒ~���&�f��� 0��Ɠ-�"%��dff� ��IDʡ��zzz �Z��tһ0Ǚծ1��1���D��s�{��-d.I�8 ;�_	��w��\m�x<�79waV�Ţ�H�ck�k��0e*���4-� ��h��tHC���U�hύ1Ў��, �C���#h�5�����``���w!Ц:k�̑��(��޼�,`���2."�?�� ��,z�U��N�R�Q�<��د=?^�sv�6�e�uRR�U<9�Q��ičLO��h:���~������߆�Z�����"�}��KQ�����2���@Е�}�C�@cjb��##ZM���z����c��y=��T6%j�E�Π�b��������gq�%���������{Xb�6ȵ��>f\O��� �`�Ӯ����z>�4�W��"��ȱ������ı�=C�k�߱/�	�".�SKJXz��AV�\�Bg����e��ӫW�#|c��� ���b'�>N��c�D�'|���B����G�GV$��#�b&�	����+�Ʃ�K��C2777�����ܘ����_癞ӆ��#��	SFGG����D^N%h���ʅ�6���E5�q4��2�2& �hj5`j�q:�4�r�������������(({41K���M��k<CXRs4�~pAT��q��nC[�������ʅ��#�� �����+Eīz���9���w�3 �ϣB:���H@�H@�9`3Tޘ�;�6�ZL��Ow�%�܇ ��a����M����M=��7�����x4��D���2����J������B$©D޿�z��5�uq����_��e�c@���t���D�dL$�J�����cs��?�@@�f���E�g8e��| �Է�
�̮�Mޠa���Ke�|���X	ҋ��	������Lǒ����?~��L�l���`S�V�QL̘sJ�d���t�� ���$���y	]Z��� ����y�Y�[hӠ0�Y]�����6��y��_	&ڽo�^��y�_ɩ��KF)������<����+��JE����L4����c���<�F���{n]�iJ����;�ED�8�i��Ñ(A � �W.�=0��\����s�Ü�ZI���FD��g}��Z6�j���|�]!�q��&~5����SDX�c��\��~��b���8'�Z���J������7��A:�%�c��[�yJq�,��&�M�5�G�3 ��S�r=���9E4��
�l���C��8����j=i��s�o:���1L]���V;l�wgA.ic
�zy=e@]{��c�)s!�H�L��m��������μ�(����W���&��_��=��ޘ�!�ٮ�ɯ�H��S������{2�m^�Zɋ꥖H�OS����3ӬE�������	��{GdA�"�7Ƞ�F��F��?�f/�x���_~���;*-�X�|Ҫ7s�'�{��f����z�Fڷ�N��TС��][F��a��~��Y�`���]/{�`�A�?/��0�~LmaڵBW(���k�����UeX۸�N�c:��p���2�^.�ذy)p�pnu����v�WO����o�]8��x� �⨴}#� F_d����,^�b��g��q��l���P!u|�z�b�!��~͞�W�o�����l�,��'RS i�߼SX�O*�\�&Y�ޮp�t���q𒔔�O��(�%O�i�<�5֐�����h[�7��1@�y��((��-=a��bŦ��խ'.m,cM`8�'\�+�/bu�`j�ze�UW�]H1M��%���ȃ������U΅���"��'�1����#��6�ye}!)�^Z�������â��A���i�����p��X�W[J�OM���	��f��]D��yV�|�T�����(�!�镞�9k�T�ǴRri�џ6�Qp�����W	(fm: �K�1|�W�7yRn��.�K�8u�<L/3]:p�$Y�i��T�`0O���B�%ý�k`̣��t�[�1����~b\�����m�jU	�j���̔O�;��&`f
���ꁁ9�Z+.�ԟ!;4���?!8�#�@�A�(�}/�j�r������Ɯ�,d�=Q�@�?6v�6�*�&+\�.Y}����k�Zί����8'fL�1l9C�N앶m��L��Z�]V< ��v���.����oRT��	V�dVm8@�Z��0��hȧ�
�R���I�=݇Z��9�Loy�_���OFd���[K`6:|ۏd��^��cvb#�w�5�*&2z��_����
.�#�'�@	g�P�Ӱ�|���ڪ,�spL�G����u�����6%���j��<e���B	GN��VdZM��;%����'�޶�d"��ģ����\��LPKr��5P4]���=��w;��Y�]럏��@rWj͋�OS*���O5g��m�_v�+���'��eny�AA� �,N�`=��Q6e������r8HSꏒb�7�oWh5�s��z���1[��+������Qҥ���|��+�}lB�p��z�����(!\�˖D�[ה��f/�
T�z��f=#�Z��j�pq�,D4(��p5ڼ�t���|��L	|!n'8���r>?�����A5��F�6���ťK�b<�ItG��A�j�����Rp�&����S��ت28u:6��J�
�[���<�mL���*j9�@D�:��po��2 ^��3b��� ��L<��;ӛ��/����4�L��)�k��k���!y�*���%�ɑ����^z��
W�Tᵏ�!um���w�8�jkK�cL*Ρ��*t��C����ccw��K�G�#c��/�>K	&�g��Cv���j�?�-��N:������tmv��zh��i����f��\��~~�qj�ᙦ}E�܁�ɏIA�_�8|��(�X�qk��N�+�f�P�yY���i<r�.�����&�o<}]����G� _�������Z�0��D"�>҄%��-�
&˭2��2��UE�"I�v��*T�D�\�h@�ݙ�JSuK��:�y����"����'P��7�M�iɤc"*wp�9�@{�~�mf�c��3N�Ze6��𯯇��<�1*ac�c~J�Sux{��kNzMԹfa\Y�	����ڏ�Q>��_�B�Aʹ�����5"��t,#6oS�CS_>sJ�9R	����	�%�k��=!�M�о��N�޴�:�nrr��V:�E5�!��1��7v��k��H���d)&�o39ݞ3z-�&R�Ѩ&�S�TBH�>�����V���mI��䍈��{�3���b7�8�uϔ�����F�sCmE�������ő�-��L!��Qb���#R7��C��&5nx��v��Z�â��kr�a"�`ơ��OFm���B�h��k�_�&�6�����~��r;�m����W\?���0��xም��i��Ӓo��ɍ���IS��i!�*���PV~R�JܕE{��M�:�O�#r�t��3a(�l�C��w�Z�>,`���`�gs�w[�������\����=���L4T�l<��b�������w&����1��:��qf�ЙC�xgfz������GG��%s�=�Vp���]����ckWW�t���o�Ml�+���>��(��m����b�j-o�+"|�QhF���/D91�=�1��VO���5M�{���{YH3�&\	!�����`���q��\���9��8; ��^���p؞H��j�;Zv��n�����.��Aa{�1�q�SF�m����c�Z�Oڠ�]3���U��>��p�ٝ�ug�ȪF�[�!�= � 9��PX^2}�%����D"���tul�����B�owKn�(�-���6H���9P��P�M��Xu�`l��7��凮�6�`*��g=�V��*��ay�ݎ��YR]�`ƫc��{�4?!���7��IxB���!��WC�mP�7-��f󿧕���9�KI,��j�u�L�
~�v��n��:��d�u 	��+�h}�?y�qg�__G�FѾ�@Ӫ���2��l_���2s�VbŎő�������$���ݽ�����&�����=�Z�c�o3�ZH�?JG�/0�?Xxb=''2z�wnsk��]���@�it��,�η��RWo�\2n��vq2�"ԌY�	�x�4u��ac@�b���[֝�AN��|���zn0F�S�V��+G�Z	l���˅I��17�R���e�勳�tH�{E��#b��8Α�*�����B�U�|u�h+����w~���������mGN0U�~����.��ʔ�2�7`�CY�$DD��ɵ�����n��G{ү��$��>3�N^�e'}/����p���wo�7��7�·^�-N �p%SAWڭ��俖�)�trσiyhЩ������{���k� ��>s%����?"0��Ƃ������G�i{�gv̇}�59����6tm��)ũ��:�m�pw�'_-�Xߕ9AF�]���5�מ�N���|}t�]�F��u2�}��*����<��0n'J@�ȉ��5gJWe�~ܨ	jH�<2®�����/�:�i7���x��m;�p}�	�U��E��|�ؒ󀑢Ì[�V�c�R��*��
u����2�~b��*�m�qQ��Q߉̚�l�`l���&�2���+�?-�1�/,�"���.Zo8���4?	=�����&�K�J<(ެ�xH��-�G�nc&:���Zؚ��Y��99���e���]�ځ=Cv0�� �Z#�"��m�mx�4���K0~��8i�S��>[*aO�JmH�;�}]5�ӌ�E�nHL��0��<�F�W]�9��z����!2⏱���s��JXH*�ۇ<	��Is6Woj��-�q�8��R�R�Ȗ���21q��#ǖ�����c˻����XXV��ٮ�����;��XN��$�͚;�-��U��X�Ol�-��<�2��3m�Fa.i-�3��^h�xO��K����z�/~����35gǖ!v�fqJs#��4��^�<r�Oj���o��
�ƍ�&Z�~X4�+�N�u���z@���K���N<9���\�?"k�38d%Mv��U���T�bg.��m��W������9âmE"e[lƢ�):�IX,;�g����d�Y-uy��V+WV��W6n{��8��:U+,,�E��W�m(wߙM���x����{RpR쳪p�p�Wr^6�lH\1�g�fƲ	9i��0��g|�fłԕ�g��?�r�U����@lǂ(��W˓�b�{[���C�1��W��Xj�D��Y���d36�Z��ڪ�3�Q�\�3s0D~n$3�v�>�QQ����怊,r�*=��q��]i�$%��k�)}6+�B'�#�PV<>��|��-ru�Yr�7�b�����n5�F-ֈ>���*�����V��F��m�GT���>����~���� �w��#r�r�k���^<g?N�D9�ؙ� G)����C\0��ؖ6���ki��fbFk�M*���D��8=}���Bn����՝V�H}6�P���,jרD����h�~���gu-�LE��%������08ߙ�Ht�k��M��=���HyIٱ� ��RHrH�[ t� �k����;���4խd�U��Aҟ,ז���b��G|�z�n/oߎ)xFJ-�r"B�O�3fe�:-vp|;Nd �8CIDk�k�k/2\�vb%��n00֘�+6D<�$�9��%�b���Dn�7��8T3��Σ�9��x������+���QO�O
�,�]xT;��+�a�]����ϵ���tC���!��8B$�����2#��o���,��lI]��0���Nn�dpj�F�R��(�O���ď�{���)>]���S۰�J���f_��,-���T����3���[�G	�� 7�^���v~��X�"4�,k�������`��@eT���M�#'.<?���k��N�oZ ���G.��1�b� ��j�c5�L
�v�o�Ww4�1W�#�5<���Yk�8������,��d�E������V�]�#g�e_Ѫ~�rti:�*�aT~Z�:Ms�|��`cb�`�h���}�������Ǉ$�O��B��S��uV-^�M~[ؠc�'����3[�l���;��	ɋ�vad���u?�-kb��S�jq�~[T����� ���4�p8-Y㖐��;���.@�ɲ��RT�t�\���/���4,�@�����]���D�%Q�^X�S�|w�E�����)�����EJD������^��}��|�!��Isz3G�W'����
�V�^T	�+��J߄��{bb!���y�3�@�$����������c�`���A�x��!���8��Ǩ�ݲV�&0��3Sɛ��&ngJK�Ԁw,��8�V�?����*F�X�����-ڗ>��U%t������9�k
M��n��Ԣ���c�L�D�ˢz���ɷ�|\��6\�� �Ӵ�zMǵ��7
y������GJR]�hu"����#o��!ڮ"���Jr�`K�K�"v��[��>��2޻���]�z���"�kL4�}�L���=�?I6�$�d%���
O~\�*@�"jc}������*6`4�c�����T��nV�

z��L �l���=�1�]�oHw����ɴ�e^z�s�A�����O�Ղ��P����+?c�E����.�Τ�����xS{��+�d1�����VU���s����0N��ه��j I��|�:T�ῑ�]+^l�����A�Rc���pt1�I�2�
T�|�wG��ihl�T�`���%e	����߿���Z:Y�?׎��uo7��d4���(�#�Vw��U��J�ER���0|�'�� �D�Eܼ�*��#�:in%|�tz���}r��
,���Z\"�w���v|���i�9=�{Sx�:�`8���{��99iZ=��b�^�L�x�p�&�����O&m�^�p�2�S'���D�[��,]� r��{�Y�XՔ]]�@�0�_�h��L�q��x�!���)�K��h�zݙ��
�������g s�Tnx�X��ײE0��|����/������������݊�V����P�HHe0Cy��x�	!�yٜu/c�r���%��ok��v�������r��ߵ��;*�o�6��U�5y�J�xR5q4���훨����Q�f�p��4����u�0�G �5k�7�(��EC]��)K)�d_�n�kB�y�ɤW�����Q?!���E��шOg����D�\���ŷ2��t��h{��80;Ns;�%�uޟ�}@t���R1�a�˨��r�t�̨[�bw������ok��Ω��U��1�t%��������:|*�BgC����O��n�<���v�<�I
����i� �1Wj [	5�a���O4�*|c��~�b�~~�ls���~�E��k�?rTK�l�3c����h���Z �U"$�8�lh�0j#K���т�}�B�a_Ử�#�1�ʽ�t&]��c�=��f��@A�&ڳ�۠�kG�m�B\ă�7�]�Tζ-�V�t!��O��t��f��`#��j��t��׽���(	���	z%�w!�3�����*86�Zit��f#q�ڕ�`�ė�y*3�����c������E����L���e��ʠC6���n��g�Ќ�l�������*ԝ�u=ph춬�u-�<MX�E��%�@�:h]7��F�f5[�s����ʢZ���o:|���z�%w���n446x���p��$*Sa08��To��k��4� �N�34��墪s�g�Oq]nt��,\4�����޳�C~;/O�T9߶(,�f���̤.�?�̠����Ĭm0%$e���42������;����\	�1&����I�D�	���*�Q�ho֜��{�D�$�N~p۞��_}�ϟ�r�q�W���uLME[�4�W6y�n�nt������� .���FOoE@�}/�EϬD��XҕD�O��\���]���uѝ��* �������B�ۛ6��>l���^���߁ ��C���a��Ʈ��*`)'�n��(��zOOC:W��ȵ�@	s��#}R?B�����jphJ�[��ivDN)M�0;lsg#���TR���sI�Ñ��k�miut)~W���чs~���	�4<˼������������[=P����A��I���ŏ�x��Dr�( 8�^%�,�{�TS��*�f:�${\�&�G��pI�ǕA�^Rz�Ŗq'ͤ\S��Z1A�j�ϩչ7�4^&�د�6q��l#��
�����U��G�[�t���5vr%���X�ǽi� a�y)ۃ�-�����??�v�����k��r�tw����?۴QB�H<����p(��,�]��ۮ��xrQq���1Ǔ��d���".�r1��^O� ��C�|v�IQ�q��&�Rc�'����^b3��?
��c�N&ȫ���¤�8�h Ⱥ���nC+~�A��Y{�ͳ���GvtnZ��5O�<��3�U��u�N�+= �� �*l��{.�e�l~��o�_��1�
	�]�1wv>P��Q7�x���� �Ѳ��(��!�S�f���.b������aċ�v���G�q����G�Y�� B��V�������6�'l��B.���}y�f�<)3�(6�Y'�����7!�U0k�F�v����Zd_	�����>�*b�y�����#i(�<Z�kY}�v$�!�;��CS��z��P��2��4}y��C����
�ے��,F20��Շ�^�<޷��)OH���'�������=kd�#Q1�}<J֬�>']��V��
7��xò�v+�,?�,9��?9G����)��)ү����s�,t"ˣ�5��T��w���iڵ�M�&��b2p�/���1?�A�/�����������l ]q�_|��*��N�C@��A�Sp8C�)�6�nx���oʆ�\���V�,|G��s_�(�j9d�`�_��=���n⇝��D@��k�D�s�d��i�����ݶs<^�Gϐ��|1S��t)�O�Oǅ��0w#�׸�s��Qd���v������A����c�?{����EThN�chm��3h���_��\E�Ҋ���7bցN~��������Y����(�8Q>�`͉QK�@�hw�����	�ӝ�O�M�OQ����i#����"�r����,������_�L�e����L�FaVAf��ʛ���0�&�]���f�G�v6�c�jզ����	ў� ��{�T�g�����Y�Ky!_B������z�z��w����`�ǝ��ć����
͜����,J�'��ǳ38.6}-3)vWd�Y��Yb�6��Vd�!Z����Op�9l��������m��/��o&�_��S��#���]���d�w��+���� mܟ�r��ȼv�����RUN�6ۈ��8�'�
|1�i���߯ �><��&���(���6��N�9'E<� ���_[y����~E�+�$]��vC^��h�]��S��c�Nm��b��⦊���.
�L쎔�i_p.�O�G!d}�VG����'O76
�r�ǆ�#.�֒��ZİfWOlq���Y�@v�0d{�y�O@,����h%Se��;����bM�l#���n[���ζ�!7�ۥ�P�u{mp��4,��lI���.�K�u%OB������J�!e��kM��z�]���+7����&Q��y����B�璂|������ﶬ@V��4̷1�ܰ�K��IU��b<��C���
�k���=6+�o�j��<B88����F���Unt�9��G��Z���ћD����/kd˸D�n�Ҕ���x`�,/v]�e�;�A�A ;�pV���������l�Q���V�Z����}���p6�̪��G�i(���?+XtI#���Q��`h�8܉r���yL���/m�����y�5)n������a�����UeQ�z���[L��m)����7BΦ�ˍõ�;��kp��!yZm3G�)���Z�^�g<3K?�%̓db����n9	�2��L���1a����c%Sd���J�4eƅ�n1�ȥ�1	'�0�~O���������r��=0n��� $-7�ſ�9����|R#Q�['�0�ʔ_[��!K�x��r�,P���]C��ɭF�[3[&�w�I�N��ii�*I�F&����<�y��'�3 CO�s�]5���3��ZIa}��69+�1bq�OB�5�'V��/��(B�yu���s��mO9��n~}ދ�����󙙊��3x;���_[��1����M1��:[k�H����̯�lU����>K�e�ˊ�F����A��<.�ض}�H^p�W��v�X�H�3+=	���f��k�tC�;Aɔ����V�g��E<��V�˒#�j�3Z֢��x�RةQ�k�Q��S���W�=m��\�j���~=W̓zf���p鬭'e���O�~�O{�73`�s�;>1��1�*g��/7��b��^��M�<yN	�/<�����祺�?�B�~h�g��Q%�����Ns�o�o�Q�(�~�!���/ːR�[:	'�=�`�(�r8Ӱ�:�(��I�͜]�C�QF�I�UM-Ua�M>���OJ]i���u*���I�Tp�d=	t�(Ő����G�$u �D��G���|���QX}�x�_�+��!��y����\!�0®(w�0�#.�-2qg��'�����%E�Li[3�>��t$� ��|~'ՄR����;�QlK^�u[:��5�ѭ�����P��GjZɓ�f�";}v�|�m�Pgt����)x�Cq;��w%�,��8��Gw%�q��8�zh�w����o��[u��1����e���ˁG�T�Ϧ6�G����"�]�y*M���y$��`l"wl��bϽ�t�J����L���d8�ia�!#3���=�'�?w��Mv����'z6=ƒɋ^�B%IH�8o�n�8)T��e
0)�E�C!`�^^UN(�?u#Ȍ5�
�_�rD	D���oJ����#���F�
�e_��4��3j峸������&��Djx�=#��p� pB�,��	f�_!����QXef.z3(C	��eD$�˴@֊ �,ZN��~�	6a�zh����������I>  ĕ������*40��Vi����?���f3�9�+KAG���ߣ>�Q}�6��~C}v<�J���U�����w,��������[�+J�H�/��o�Y[���kd_Y�/~��-�|���~dx=���U��W1c#n{�%
K$jE��9h�t<2Y'�WP��{�ﯡ����#A�)m��Eݲ-�-p��)a�X���f��|��	�/e�[�߁G�rt��Һ���E��y�{J��}~U[rw��hc��x�7~.����?��M�V��=��pM�����0e���l'T�<CH'h������u7F�<�W<�x��a��dҽ�㨫����*����T�IgED�J	J�AB��WE�.]:H�n�B�Dj� B%� ߹xyޟ�����br�̙s��:s��1}�4q�����C,1_.'���M<c�D2���Oπ��<�hae�)u����v ��IzL������F�4�)���_t��ȕD�}[�k�6�B!�T��&��/��;lQ�v�뗽�t�h�sS�ɯB�'���O\��7��&���������j�s6-A�Uo���u�7]Ώ�[a_�sq�:��d�8������Tu��W�&'��uՃ�Y�����m:�tr��w�:^�j���B��J}w$|���/O�c�����4t��� A���Fg�æGݻ��/���A�Y�B:���	?��Wsh�,���|�O����`���H���sv�ɨ$�$L����Zn�N�����H4�z�,WN�z �)�Yd��vEA؏gUg��ˍ-H��x7��tfp��$��_;qz�^�)��wS�[�rT��V�W	8"G�!��WF�w�(�@~�}�	�)����ʳ���Z ?O_�t�a'���e����*��1�c�-���.���r��}q2N|�}y~�(��Wq�Ni��Z����$#"�߼�0x�ks�i��F�0���^�T��]
*&\J�����he} �qif���K냫�d��f�.�.}�+�*k4ig�d*�l������ �VW�����M��k�E`7�l���h���S�	m'z~QTGN����]n�:���1r��@�@;���$�����_&ku�/���;�Π�ѽ���+�t�$oַ�����iD���c	�y��[�}x\	����瀃;+������K�����tWf?4��-�ҽ�YK��3�jc�x�s4�yo:��}�=�[W����E��l ��j`�:��W�a(:p���Rnя<��iW�*M6yi���MmE�;�n@�\� �H�q��\8K��S�C8l��U۷�Ǡ�z��ӉP��h�l���5��^�Y(r��F����Te]����K�0�Y?)m���^��率���9�i�ژ��뒮c�F������
^��sR�[iXOWX�Q0�b�/ϼ�p��G�l�?�Y\b������ �X����_�&��m�%H�����>+��}�jn�~V�~��F�3���(���D�C3��lu��$2խMER0AJ^+�ё�8o��U1t �`ݮa��:�穽�v�N�i�|e��閘���~�� �>�Ǌ���>�TK�T�����օ�t���s,Wi�.�ʯ�$�q0��o�����\W�n���1�?i�b����fg�Eq�!�����`��Ս�+\�::-δ�q���O��#k���v;�]t0�k�?������(l�0�O^����m��.�n���2864/�r�����TO�WM��Ik�w(���ۍ��[Zy�._���f��¡4�J��-��&�	��Y��������}��-a��{��,�T�`�ʶ�I?{��C�o�٫BNv_V���;A�}=l�%:w�`y3ñ��ŃJ��:���`g7���&���]gu����
v�>�+���F�j�<L�=�N�笛�lI��W�Rc�Е܃A�Zm��5B��v0��G��j� 8sY�x;t�%�������d��N@��.[���,0Q� �*�/�!��~���4��q��6úI��g�K��P�V���j/h���s=���^E�'���Z�GGc��gǬ)�/�F x|��_��馫�O��Ё�Og�o^�|�H�)+������2[1��D�i�;�0��J�*z���'���a,��	�{���0�m	c�[W���ͳ/𕚤�ؤ,-��cb8Ulg�Zk=}�%��,�N�n�����f	��Jo���\�ġ�@���0#�o}��/	^6��O
 r̚��V܂����#$�����ט�`�K�Jǎו^\��Y�rB��C�D��r�c��'���m�"�8�O�U�=��~ �#z���僸�o��@���8�;��d��&�^Ԋ�����=�᫝ʰ��G��v2k�[�9�� y����i�FBģf���(�����z}]��;r�X1阂ם�i�׀�!�*㈲���|�q�4"y�, l�����*����]LX�\~���m���N���_\����r@��p�}����`�HMǣ��M�J�*b�_��=F�+�%�Ux}��B��A �>JfGػ6ALJ�V��~��Ά�t��7TgGt͏�,�s�1)*]�\6��쫙 ̭���t��#�������A]Q4�8�W�Z[[u�k��ir��F�.�ww�$�;��a��e���l��w*�4�O��Rޕ���0-lQU��*?#�p����&��s�/5�^b��z�*3�K��w����
��T`�[��nV/ܧ�A� v�h��&��nv�U��Ȼ:�Up,`����k��
�Ba_]h=*�)���.~݀d��M�.�&|���Uu�\�����l���PX�����脌\���o��O�H��X\�Y���H<NCII	��y�^��5 8̚�����C�a7 ���u7�!���!7�zt���7�>�nf �y�+W#�3��rƭ�W/f's������'�åk�����uwC�p�~������)� 1���h�H�:�`�� �n�I"2�2~3������.#��I�����F�}�uٝ�q0�e����^<������g�3�4]��楤܄�v=~�a����d:L�c���$�R�%�;]G�p(!#�˥�pd31f�}�V��sY'�������L|X�j�z���ex��	�5-��&552}�m�tө@¼��6,�2q�M��b�~@�i�P�-;~�ڿx4�_F �M�������ć'��2,��f��=����O��[�׿�>x-CT7�������i2z�_8�z	�}%bB2Ew�7�y���/�B�����t@O���_�~7����/�k2�d=��=�dG�1�(@V6��T�f�B*an#��z9�/ߥ���K�v���l�G�\�"1��U�5*8.�3��r]��'��K:�W��Ƥ�>����S
�X4l�h�1�����1A;�g�\��<��7���߭ߍ����*�8��mᓓ���0y�\��*��ۛ�T+>(��(��Dy���,��o�%���/�U��]�p�x���L�G �x[������3"|�)"O�_�+�K{���8{�-�!)�"nk�����f*� h�f����@b��!mrL�srs�ʇ2���^��0�叽fݢ�4�)u��e���g"R�-f�~٫��/�X͔�|t��.�@��+j�#çt���l��wbw���l��]�56��2%��Zy��6��m+X�!�.8ő	 � ����T"3�U ����v�h���,D������3QQv���n`�{�v�Z�0�%�t���R���W9V.�V+x�Sz��h�nrҰhgsuvu2nX$�K[�c9,��左�Ʊ��u�ܟ�VR.�H���S���-f�'�.��-r!er�l��	���y��0��;��0���Μ��I�!7�̔�z�D�A77F�i
ރ�'��	�3��N���2�i�8�� �*Rw�������u���?���v��;�9�,��n<���3�#��}����M��������j5�����A9��=��C镕2j=&(����e�'O�퍔kv�P�[�w�JF�ok�yH^P*�땭�U˽��l�Y��V�TA���FJ�� �^���r�l��T��lݮnm�_Z�h��=��I=҄[F�� `��w}��t�J+@2#�~ -41�--
�X�U�T��=Y�Lqv6�ߧ�Ta��5B\�ș�����2���wGW�p�b����k6g�����]���q(B�Z@@@Tn��t�{ڠ�������]VTƴ^�7*��+6Rnkl/Hn����©]i�~Tn�=zר\���-�Q����+��Anm��!F:Z%��a��u�u]�y��jS��s���ع���>t7~��YZh�"��~�����ׂy�PƺI��(��|����S��Km^ړO-LML��X~!䀽�����cG^x�x~�I����b�6w}q��P�k��k��Ǐp�����|�W����p�P���A^ݼ�`����L�u�?�;������j�l_�җIN�oO�$|c����I4�8��SUHr�'��l�$��y��v�v��5�K+*��ߋ�PG��,�cW��_x��~�-�2¢�b([Օ�5�F�̸���W�a��sǋ�h����>hr,�U��=BO��oW`���S��<]���#��5�㘤��_��t�l =��,��}��GMb��^�_B�*(��j=�����jW`��l�;	]:t�s�V;&�J�Z@��}'�|E�T:������6��BH�|�h��H���s?cOz�i��1��N��!��R,? u�j@�w��uQ.�������yZ�Nۀٌ6�CF	����wc�nI�jvC�RK-�ε��w��Μ��9�̗�o���L5���|��<�4S��Wu�5�`e��
��VIl	������nܙ��cٴ����L�]��R F}�40�Rs���O�B~}1'ے*j���ZJ�=["W�Y����q�6n����v@u���s�����X ��ia�6�a��sNsC�}s��}������"l��=�	ٚ}���/�N�M�*���WӅ|��U�!��O^V��fp�&esR�������F�2����=,wLȯ���<�8mAI��H��B��V���w;0Dyg����D�ƣb����B�mo�pr&v�����q��
 zSb�A�5ͫ;<���z�5ވ�6�=x�?���[i����;v��Ы�S��(nA�o��: 7���I@�Mm��\����,����U���SG�Y)-�m[C��`��D���K�~0�4��^U�?���5����ra嚻�Q-�
�4��U*�����7��wxr䵝�+e���%1y�!�V\O����Q;��>v�baS}%ı,M`��c�ce��n|���o�K�fI��9+��|.�c��v�����M+G���d�Q���1����QMt���Px
���o��ǏM�q����	�����*/�R�J�M�x��@6�۰�%��Gq���3�'�YVM;5��LM��s��{.%�◫���m����7��ݎG;|��?����2v��������/ΛGZH>���K�3#ڪ��~lJjJ,��o�������M�p1�Ƿg��3��C�	N�Ya�jjj�%/�.��~l��b�7�����^iM����w������i�Q8=�� Μ0$^`��Z(��X��CIJH̛��ӓ�q���Č�dQ�)Uق������5�=��-i���KL T;�ʜR�;���>�V���1'i-?��9ױ���-�]�����f[48]�m��JI�KRF&a^k;@�«���3<%����Ro�����t�X\�{��i�A>1�O��>Й<�1�Lm�w{ǭ��-tAb\3ڄ�0��:�~��b�GI�j�d���+Ű��":���r$�&g�&���3����}_���c_�<������2�C^4Rhd��0Z�rH�YYΩW�d�6l�v�����k�}���V����[�W���݌d=wn*9lll�K����C�@7�,��PG �g����PKtu�ʞV�Yl!7MdD
(u"ѳ�I�M���YgX���H�L��I2������R����A�i����$�D�����O����=<u���rw��b��r�ތ�z�2b*	�	{	,p�|�WGKYU�����nŭ4�<Gk��j^�W��ѷ=,K�Okj�9�>!�7.Q�CZ��,&fI�)>5;�w��B&JT&g "�����8#m�ӥ90��߷z�����vR?�?��l�d��K̳H\2Z�j�튖p?��9�\�9�;#P�NK����D
b�(�v(t���O�GVo�^V1W\���l@Pv^�c*O�Y{H�����U��H��#+����&�v��?��{z"rz0�g�08_K�ʻ^ĳ�� u��z{���ߠ�$�
�Y[�Y��5T�*�}��5g:��1���{�т�ETy��m��X�$O,�آ%
*B������z��+�{=X�޸�5�@�#�]��9����1M֪��᠛}GϤf�_n���nOʳ|��Iq�-��Fջ��k��<�J�7q�
)�2_t^k�Q�u�L>��Qs7��c\N�0,;���궢�#!���#(I�p[o��Y()��Y����@�Ы.�x��{T�;�F�8��W��旡���H�J�b	�5�����V����沁)6�2W������Ħ]�e5R�K�����^�n	KHH zBtM|�%���פF��T�Y���E���%�B�0�����n�27b
�����D�!0I�h�O�[u,�ٻi��"��xc�ccxPni��t�Y:o���f��Uo��5�缵>��g?͡�\�8`�>Ojx1���>H�a6�[�e4��g�P3�0��JC�T&̆������n�qv���j[`�g�y6�|r�P�tn�v���c�o���F��mmm�-������<1�EV�D�q֑���D薾0�.6��w�	���9ۭ�`��;�nM���qF?=�g>��h�j�1�Y����yEb;��l�n�xתeE?�LtB�a�2�o�����<Gq)S��b�y�6�Ƹ�ZO�b�Ȩ_�ـ��SeQ�dM������kݏM��t�Y��L%Qk��M�?�8~B����x���M��}�._�������k=(��tmAtW�<������^�[��CԔm��ޞd�����p8�A~gɇ�Hj1���Xzmv���~9�<� ������*F�d�96�8&�ב�TΝ4J/�*/�7�>�E�V�U���m�Pߙ �U�TT��H��dG�F�m؂�h���짼��Uvf�^{[_��t��Z�7_-���O��������
�:����P�l%�J�����0�ø9]���dsP�p:p��� B[��sI�k��Q��ND�.����|\v�S<�p��� � �$3BC�aa�"O�dUеh��:Q�J��˞9�-��,�$B9��`c�a0z�;MU���j�jr�+��of��z/T�g���������'��j�8�2ǡX��������\��H��|%^v�)�����M��՟iF��f��C,���Ӥ�xd%W����D�(&9��_��qt��Y���#�n��R1��){v���g��g�%��<�;�ځ���%�[���LO�F�u����}�� ��I}L>�K��9�Y�0}&�>ǂ�p;��|��:;xHu[����e@9���{�,D0���
܈l*i��m��i�HGI���r8�6 �X�c���h%iQ�"U=q|&1z�ˑ*a�2�#��k#IP����*$Ȗ;+�K�pn�����X��$��T4��� W�����|@���H�=�"y 'ǥۅDs�>E�D��f�f� ��2����OU,d��* �	}4!9;^rh˾�v�0K��sń�2�)A����\�qn�:�dYru�n�����c����C�Y�'''�P1�<�����*Ae��^��:��^���IJ&	�M���w$\�&�%T�Z��^��K#V��oN�p��,�޾b��+�Br���5����1re���F.a�Rp��ׯ�'���}����.�c-�4ຘ�j�IbWӳjt[�J�0�;��T1Z�<���i�c�3���B#��%��g��6���b�61�D�]~Sk�����2T�c�<�������d��=��"4��Wi��R	؞X�<a�~�)l2�r�r���̝����»(�JR/���t�N&��3aD>t�`���}�*M�*L'���,4�"�y	~T�%Ҁ4��g��N���U��ER[[r��Ź�"��xi�F'H#ևܭ�k�}H���%�'�'�j}�L�G����.������Ġچ���\�o��b3x�X6z� Qߑ+if�~���sR���%:�[�+���M�g�JmZ��������3����h���pg��j�v~�r��'D�32�%���gڪ}��hI�����At�n�֤��eu�������f��sZ�:|Q�4�@��:{xH$3U�~�_�O&�15�����՜m���WϏ��;�����;��K��;�s�A����^�7��7����&T%
�j�7�6�%J�"e���l4�>W�\ (��a�!����nL?�U��/L%������e>��>Q&�{� �����j��lLgn\��E��*W�{6!�����Q]���\�P<;�F��ʫ���-����		�r�)�w�z������v޷���egr���928���Bvt�7�,l�����N��Α H�� 㪮����c(:�'�y�"L�xΐ��p��YU0�rdy>QhCE��c0��^t"���sۑ��)�tT�L�m�+qf�j�_f�G���v��_���u�z�D��I~H>�2����?Ҩ5`�N/����8�&����"g�;K��.!�kM�T�4Gls��u����B�l��T��lu5\���_��:m�d�"_S���>�qM�cKs�Q��۱�X|����J3��8�^Y����L��l$Q�`��؛?�R./;��������+r�y0~� �3�:Z�MK���e�>?|�p T�4��;U�WI���n��n'IH
U�����o���@ê�]NL?B�~�(Jd��s��_H�#�|=�B�%�v�Uk���?	'^Ř/�+����c�}�5���S��˟7dy�Xz�[���L<��1��GZ�>�%
�O����xK���/�;��2��{yRӲ�3��2�X�����x^nN"Ԭ3\�yˉ>��Xb�7%0��D��M��6���]i��V"z5T^znZ���^��k�I�┌�#�)�n��/p��m�>ݝ�6>$��iQ�~/�'��)�;��&�ؚ�qi���������Q��lZ��em���(�7����(��B=��zz윤����~	�r���n)����!m�1 �������$�wRs��R
��Z��J"W�&�g��� =���*KX񃒉�Dm�U�o�y�R�3����m5�zv����޳�4�4�U$}�=Z!��!T���N�$�7r��B,�Sv&J�J��́��ܩ~�uԽɉ��3���Lq9џ8|g0�9�3��9�_Bp��!��h�(�_��.�U�<� H�r#�̞0����Pl�Xt	�
��#� �Z(H������ezO۹@ �E�������/�=�F�w����d����=�3訛������,vR��i�~ߙ��CN1+J�oO �뻤]nX���@�n�q�AZ%PY����A�-:�v�{ڊ�x{�C�M!L��.i�
Kž6fä�
�o&�i�Ƨ��s�Y�`�p�\~�1�Y��iV�2��M�����!�"����hUM[��q���%�͇<�Q�.i�v��1]Q��!7*�����=�m���e��~Nq�����!cyL��*�e��p�DT���}�v�Dz�u4��Z�J��m�K�J�L>o/�	�V� ��1D[�t4��f�ϥ㻾ejm�+~��뗏B
�O��a�+J�<1[�i{��\d�揦����@�:�5܄ML������~@H�k� qpF�(
��i6t�w{7����C�M�1)��C�1�ZA�ҥ���i$Y	�e$����` ��3λ������F~v�E hb��B�8W&*8����ɛ|v�T��](99rR�n\zZf��*�2-������ĖIX]]��.x'9K5i0�i�2��DJ�D.m*��/Q0de���¯���`}��}v]X�Ў��'��Ǣ���͈�p��H�h�>]ZZ���Vjx��[�]�S��iI;q�hgυ"��O�~��_�
Z�z|��S��[�UhC���8OI9VD̸I�����_�]V*
D��Q �]<�p�����I����7P�o�#.Ck�@|� ����֖�9J�� �
.G���n��3��q��m�ȋ]�Qk�d�A5����~_�S;�h�_�'G�y�J�)���N�?��Bn&�K�}`�be)U�Bư�@�V&���[f�ʌ�p1��C�ǁ3%^s����PN�{��*�Xxi�j'��!�.��b7{��G��*ہf<�v4��`P����D��7���sϳǾf��v?��M�.K$:��5��,jbFn(J)�BR�J�&O<!ї۸�3t-�-dpQ� �ek!�`hf"j8=Չ�aQ׳�f��9����o�&�y��Y���&r7X���K6�ި�L6�;@���&	������eq �4��+�d(������=�j��9�u�%�r�}z쳆`K;���?�unv�k��t�s�kS�fu%jm	$�_�7��9��վ��JBpr[��.%�g@4�z���x���s��]���n�]������r���tc�12m��Y�M���74��툪7rq�A�慨@�)�mЂ@�k�� %
x%�����$�=l�R�-5��аˑ�Exࢷ'��^�	H1�5�rXڲhWwB�erҍX�a���nk���G�v[�(�"ۂ�fP��7��*�1R�~��1H��	�/��p�jB��� .�\o�z7��>&����GW�;��h���y�Ѿ��=Gk�����P/3s\����2 ��5�T�`'}����{�@��1~jƾ��0�*4?}��Q�u�\"d&X��;��{�C�N��,��a����4b��d��u���A�h �ZR��x�ڧ�<3LX0�L�`�{�D��� ��E~*M�G�4<�
ĵ) =6�T��ȹL]���z����v>��K���'�#��'�n���>��]ZU�K�Z�v��������ِ*�_�[1�t!�J� �W�r"�<�� �BYi�c
���� ��_Ly$�A�\���n�l���e�Ӫn���5Y0N�Ά�y��D;�Zk�C��`��p�Qe����	%e�0ݜ&�7��}>��վtJ_�mޜ5Zm�8�[s�����R�k��]����a��d�A���`�r[���W�\�P���k�K>6,.����h9KX������A���AG��lm��`��e%&�+�N�����M�_��k��= �	>���/��R�ݵkoM^;q�j�R�%� �A>�)��ùL}ِ�u`�Ì`zW�.�6LuxcP�O~�i��!����~gO�2�J_����_���}K=1�\FL�l��5q�p�bd�o����>;�n�~!��{�OM+����%@�^-Uh���OOl��VݏJm� � �)2�Fz��r�i��Z��@�2K��hW�#�I��׈(q&63�gg@��Ci8T�t�]_��"8ug l�"�W�	xD�f:Ż���3}����~���b鳪�$���8�f"�2N��	����g���þ�ЍA�P��]��i _- _���Y<��$ew�YŝWo���L���TG�ϖucD���d���1Q3�v�B��C��[�ò']��=K���2�r��0�ɐ��SjyL䄆(wWnGL��1u�� 1r�9�I%��3l�	{@)����A�ԎQ�/5��J�0��Y��#�!��p�Q���Hj���P��%i��#��v�y�v[��2dX�����1�S�%�T��7��ӏ�" [�nH���ڥ���^�pt,c�c�_,�`��Z�0�߳}y��`�;1w��������`K� �@�c��]9$J����7�`F���Wn�~m�"kl-���©�#hnY��#/�4�Ux�%��]S(���c -Or쬊��j��fE$��w�wŗY���A�&+>�,Rf�E�K�!���P�]�ҳ/xM�>'�F^�{�~�k��9uOɞ>�d]I4I؎o��x��9�V��ܮ�hS?|wd@�j�̶�k G}qB�8�Uj���L�q���#u�v�{\����C�˓�4P���ż����B�c����ӛ�x]h~.�`���J��2ွ��9$7�L�IL5��G��\�o���P��gj������z����l�c323�o�>����Jʒ\����˃��,��u��^�XN�W�K����?����h]S���x�Db(-K�ޡ�]<�=6�
�R�;52�ӚPB5�x��M�v�F�=�	�[I5(|��~o4��ȝ�Y�ԏ��.Yj��ww$��Y�?�>Z��Abqdgȑ+7o�z�r�ʩ�S�e�䆏Ys� �M�K&��ʇ唦Ծ�Lhn!ќ�y����~�5$	��a�Զ�x&//�e����ߗ�w�=e�K�f� ��S��1AMh�fPs`����f��~u�����,�>/ e`�U��5��S�3Fa\��wgg/���]���Dul�{~�X?�Ez�w�^����[E0�V����y8� �&X��DJ4�_1KF�ti==J� M{�յg�"�R^�V U���$lE��6�L
�>c~���H85=h1��[�'��*�v���t���n�z��)1 ) `R-��ٕ��^����Ԑ��Jנ��:hu}�_^�f1�BI91�m�x�0 CO���>U��^(��3lԽ��=����{ȄNCeee��l-�Ђ�;�b6X��J�O;[O��h�ĭ�<X^.S�'����&���E6p��ԑ.#�3&�s	��Op�g>-���~��a�("�;���9��Ώ/M��i{{o�����a;��ڑ�F��_���x�N�Ўd�e��U:��8�E�)��8������%����9���>D��L�є�&'>�ݰ�8�M�X���?��)���>��*.f���E�j�!�BU�۟��B�s1yh8��ں� ��i�y�~SR~z���lR�`���ZLڝ�/�����#- ���1���c�N�-�&nL��dк����\�>R5�g9<����Nd�]�:���	R���rMu�H�4,�s������q2^��#I�i�~�}�gM0�#������+��+����$ƍ���줌���$���$l$���i!@���#�� = 6��Q:r������^I��l�{��r�G���J�Ԥ5����[|�q���m�2���	���B�a�%�ZX(Q��٦�ZPe)��E�!��r3_�i9%U�Zj6�/)od3���`pw���X�^pl�	��]��Y�5#�6�E����S<w��w��I[��[�V���S72
�����ho�=�� ϗ3�:�>�\s��b󦰔T~�_Ϡ5$�"8�+�X�~���|�E�?����������~2^���3z��N�6�Ա��O��u��)����}Z�P�>��la�p��Z�m�_�֟b�e�h���i/���+���=�ӥ �ձb:#�,���j�{zM�<�������}��x.����������N�6����rˡ�Ko᭵�
�OlS���NF�Ğ�[���g'����w�����[VWW����T�P�ؼ�|���2C��93��b����j�)��//���_�K:_NMM�qtDC���\��_<����<�Vbr��X���1��y9�/9E�-.:%�u6���Pմ%b���ǖ�W�dWu���9M����*o1�U��x��2�fFʩ���5F�Ц�A��e�8!�;RiʯE��{�D� p>���Ǐ�~�r�$R���	�i��`���xt���ϗ1&o�~-t��z��I4�}6D~ǃ�¿��!�Q�2��3gơf�"�n_������x��:��%�� ͈s�j�&���Y�?/�'Y�S�b(���+p�o��bdG��J���]��,r�(>"��W�[|<Ж$��Bq�c�'�r��o�����6R�<)�V���DT����P�[z�`1�$~2���	,ԸE�W8MX��ʊ�@ٮ�<;D,��]#�`�������vh�yx��ٹ�i�{����}�:ٜ��!�C�6�
.��������x�w���#��j���!�nZ_��YS�{}_��Q0Ǧ�r��sz5�ݤr���u�}mv5�5,'�Wrsrr���������oZ&�d������]?ʺ�|���+!�T,���:��{i�s��暍:�=X�`)�Ơq����|�N%5Q��=[�3��[��1L� �);�V���_�
VI��[Db�-o��5hK�nN�ᄁ�������J�?��.l�&_�c���V�c|���^n��W+��S��|z�S�����O�Є?c�����7qD������y��ښ�c��K������A쟘c�Ρ	8e�lu�W'�*���P��B��FȢI���#��g�D���sFf ���l�v|�9O��6���W�!�����Ib���9&۶����-͏ݶ;��K|yy9vn��3�rC��{526>�׿�"F�RCz&����D�{�*�;y2�u���$˓�/���IzW���P6i��9�}WR$+�{�YZ	W�XZa��M��ua�w��ӱ�/~-t��kmU_#�~�ɨ��D��������:a?2�f���\�k��wM�ϐ�l�;%���6!���4T$XLRo_aE<�G�"ot�/_�E�Z�aº A9������2Qr?�������L����+�w�ݨ��_l��L��ƯV�Eb��}=8�x�=\����Ɩ�����? R��{��PNX|n��z_�	ԶV�t���3���}C�b8t�ѭ'�Sy��4�CD�o?��#���-�Ժ*�u��ω������=�^yJfF�X/g��s����3������@9\~Z'�����l�s�(;���g�r����n`u��]�=Z��gBR�v��">��;�ŋTA���l��9!v�0���������7����:㊀��+�@�J,C���o��e�c@Q#��������
���CX�tss{�Ƹ/t�@7��L��4�Ғ	moo
���6���
1����Dg��eA�_A�����M2��Aj�������j��&��}���`����6�&���)t�ٙ��N]�W��_u�x�S���N��ǹ�Mb��_���=5�.�����'롽� ��ȉ0(�����q���=�mT��l��`f�J�����������7�7��M-Sk)�a��O��&���L��(ݳc�I�܂G�����t��7(}�΍�3E�Q��V'�C��Vg��?�x�����߳�`>m`�������|�՝xƄ;��w����.�*��/}s:1�&�J[��C'���U&�-�|j����$���-4��.�&1j��$T��"~�Z���� h���ׯ��d��A�0��������à��\g��.`��J����x��s�j�c��v4swr���ޛ�:t���5�#Ф=������ç/�@�����m;-����ĝ���k��'55�������-����5�;_g�?�K����x�l��E�MGG��򣽯�
=A�D�|kLY�UR+���+���P|�W��v����m���,�@����s/r����KK�ߌ'�BB^���W��-$��Y��K�|���:��g��mq�/����;a�J�c0��7U 7bqm>i�z��V��m���Ǯw����Y����A%ї�0~��k��7W�L�X�����O��9wmVY~�tO�^jﶣ ����/���DT��� ��D��Ɍ��#��D��Ћ��u�Y:34Zl�A�r���M�IЇ5u�;ߡ\����C�l�������Dog���_/#PәI��,O�\�u'$�Ͳצ����\�4\b|��'3�.l�m����w8�]pCT	N��:��KKK�L�G�~��&bkg�&�3�*٦`��O���,|_e�5'g5W�E�z�U��v�%�x]��}P�K�_��.���@��zz&Eµ������dÉ���6��Z�^r��%op�6R(��|lx�LF�0��� ~�DO˹j2A��}_T�!�6S�1~@�/E21��zK.h�G���Q�|�c��@M �m�Y%�}��db��������3)�?�31�0!5�]�l�����?��ά�HWCD=�����x�����w��U��Id#]]�	~E�xori"\k��P_�+���`6ր� Iכֿ%I�,`f%++�|� /��{��	�,�)��\^^^�>CF����Yl�`�>��u5G�Y٪i���T��Y���+l`���'h6@����9���]���R��Ĺg����M��K_�C��?;=�Z�l��SK^{-��zŷ��Z8�bVʌ�~-�E�K�@\k����V##�y6������eα��Xz�$i�����h�]J9|�k5Z���=�}N�}��J���b�I���O�س�9�s�عf��3U����;5�kB'�6F���G|��A�6����-%&���A�8Yq��3�m�����X�ǻ{J�(��o1>�"�q����*�	��F�0�	d�����=~ iA�������n��l^QH{�T_6�����m����� �:߀l
����=ON^��4�<8������g��&�HRϙ�!��0�#/D��zoL}x���0�����`�����o�>�z��{�	�@g�]`�A5V`@����|f iu=�l
�R�
w]�������fw�@q^K��;e����ډʴ禪�N�8*�!�c8r��`�%��o,Z�pR������YqQ�Q���8�[�%��Z�3X�w�����2�����|m��%j���	m"S���o�� ��O��h)>&ÈY������к��f�/�:��F>�8
2����ӯ���,~1R��r�[�i�z�ީ�����RGs
�?�>�砼-��mA��:�/���Lp3�7��1��Cj1	�^���k� e�:66�����:�
�s�#~��`8��ܬ	�ZzA��������ռ��#~��Ǎ����	�>�9[ gyo��|�]�OS	wf{vq��օILR�,��ٽ*�z�T0^����>�c�~F�(|��އ(��	cu��\B����g ��r��l�^�v�)�\���б:#�-�դɍ~lux��<�&ծ��2+?��
LPI������o����+-{/�]���3p�Ԑ�Sb6>RFd��D�]Me��/Іn�����b{__�,��zVxP��j��c�ɞt<2�J�����u1V��r7�mbO���y�;�{�u(�j�w� Ғ�A���!P�	:?�E�F{���?����9(v������,o��Ю��dA�S1���o������rR�&Ɂo|4���c��Ӽ��Ҩ6vV+�k�H���
Y�.���"s��8	���@�[�B�g�
���{ �C��x�,�F�݋g��wQ=_����ZK)��D.���Q��� �@���)/��:h�@x��]ڮ��Af��-�^��؋�m��4��c�f>����.���l�!_���c�����F�������
L����l���W'u�2#���3^����Ϸ��_�5<�X�m���5v��w�3���".�Q�͡�I#����Ng��`/Pv�p&�����+�a�Q�sy/}N�i��������1R~��S�6���J~/r�VF�3Pô9
l�/K��8���j�b/R*��Z����BK���S�lu�v����]T7�2(-�{�0��J��g�9�ˑ.�A�������H��Zp��J�p)l��GL@�e�>��P�{���u4�8��B�ޛKX<l�'�u�������{�yAMT�ݺz��M���۳)E��#;�Y�x�u�z;���x���T�O3�zG���o���z2WP^��C�	��=�q���>�։��ڒ%�'��t��68 �u��e��rj��ݾה�
�Tʣ�6@���w����dojY������"�+����D����|�.u˫	K!�l�=�8�=�*9�����dT�9���Ç���l��AOG��m�W���i4�)i��S�W"�T�]M���������۬y�V��.��(�S]"��[(��8��޻���B��2��$I��BZ�Z+���JTō�����fi�T��I8��H���?I���P��Ɠ���c�-��Z��a�(�@DB�CZi�nPRZrhT��n�$��A%F�`e�a�n��������%�x�l�X�^������31BJ$���ƽ��Hg��������I[�7%�掸�`�_8��Ғ�#�� �r��4�	�b;�~x8(7)����Z��V�O��:�_s��!11W�>�Uu��l�c��t��;��*ãS<�Ӛ���5�'4��^�ϾS���'�f}��R
ibg��s���	vR�����L� 	�[!;��J��I
�Vήf��I�S_�ǝ�D�vUf���	��h�����j��u������h��6h���e���D��r�F[�C���5nv����J�%���)�p�(�2�8"��/M[?>�"Sd*q?_b{�,T�ض������ez�(H�>?��Y6��]�����r���O8?�� ���Kxjr�bǓ'߂�an�U����,����gv�4���q�~[R��R��q�����9wt n�܏�q����Z�6�֒��y�>�~ڸ����R�;+�{ �F�x�P�J�>2ho:[�2���f��ô�:��2c�E�F*	83�l{3��M���ن1&�u�7�WQ��E	Ѻ19� �v�׈F��%���'�[D��sz�ģN' |�ǛZt8:c��c�v���`�N?�;ڽvҢj�S����E�=���g= u�Je�8�Ѡ�&�Q�-�E��&�ə�o�{��;��QY�����������W��X��=׈#�X�L#F��L���0E:��������.���M�4���']ϩ��.or0<������(�!�c�-�m?���C�nh�{�6p	�y�?��Ъt��g������4�ӇL��O���ޙm����^,��zt�joNu[U�a1$��{+�uz�	)5�N{��(����M�<�ڐ���{�ȇLy� q��z��׿����UD�X�{L�"��JA��v%7�G��]��gk*�DM�Q��="%d
~���s��9�ۘ�e�п�����f`���O =$%##S��61�v�}�Ȇ�� � ����KQ�eq1bfo���v�}�~��4?[GvEF�~��`~n2B�9���`�8Uؓ�7�uDb��z�i ��	�KU_7-����\U����Y�|�y ڋdfa�ilBrqW9-t�6����qm]ݢХYc�L�}ι8R��@�`����a������|> 	*}�t����;.Bs;���c`t�ifؼq)�fv���(
���}bbuky�L,��)u��b�Pr9�Z��[��rN��iWTD^�A&ehhX�cf�4���̼�3���6�Z;vȸ<�N��Z���w���j���yh����V�O��P�r��)�)λ�)ej�^��Y{��$��S�z٭4�J�O���Ylqvm�m��� % 1Z�>���aIU!���U��8�L&����->�f�(�����ZV~�z���hl�]����n%��V�<p]Hl��W��o4xeh��P��{Tફn"���P�� ��g�g�j�K��-���3:�Z'P���[:�6y���T�2���[�D"����Y��e��T�yWtu1>��TB�H�Z3��x�"O��� Gy�:aZR�?8�
�ѫ��7��y ��Y!&��������>GGJ��陑E��	c�6��}	Q��C{��=ʢ A�@QeUK��t���9^�2A%O:����`��FL����/�	Z�h�͝�یfES'���rt ��G9��Xc��) .&�ieo_ ����n�b�'��9�~����sw8,~����O����@N�tG����x���Լ��\�cߓ��i����r�����e�|�h���5�&����?�F���<�Ydu�-bS�ڬR�yU�E�η�!��PY��^F���}s�~1�op:U���f-�c��Q�!�qYa/����(eb��_u0O��L_D}1��T2�ݑV@�-�MDI<�0d~���M�"?�Y
@��X�eȠb��C��a�H���I��;�>�bAL��d	_U�����k^�4h��ǁ��n���f~$��{�I��7լ8�ޚ�z�:����P�~E�=���[J�~�vb6P��dԘ���Ϙ̵�r:7���}`�흾F�(�_��8A�cp�QU�����[������U��-�j���!��0��m��$��<q�`���Y }��cP��sw���:y����1�i��nM60�'�+pA���@X��e5&^���[���(B��ZG�yQ��'�x�rRטXe������i�ǯ�r����ȁ�4w�g=��p=j��a8JC~d�kk�b���"���&��pj�%�r����;��1?֓��z�t�A�ᾊ�L]o:L&����K�1��22���"K�x$���� ��Xf����d�	����>.�|���39K�%>+W�&�����sG�9��]����b(Z��C�]�F��(R�C/�U_�W�wˤ�I�3}n�l��t~f���S��\[pCĥ�g���{2��:���Q�Q]2I"/gba����Δо���P}�qC2j���I�HE�e���_�ϳ'7Ż��͠��T�b@3jz�'_"��୮ep;3U@� ��;��o�+�l�]�sI2E�o��1-:�-Y�F�<����x��z�w���Y�����+�_-���0�$�2H�����SE���mk[\��k�Gշf�9�yл5u���' f����b�k�u��^ . �1�ǭ�t��}�Խ1��A���b����Z������x��aYCS��ȟ��IV�/�ml���K����+{��~�]���ѕ���%!�y>4~�T}�\���kZD�,�d������I UX��*a^�q8��}d$)����8e|�c�VYBO�g� �v�|'��t��s H\^�ZT0�G�FJ���gK��l���:��'�I�q��>����95���Z�4>�Lm��(U>�q��X����~8�rq�ā�q�ԉq��jE��bӠ�¿�}�Şd.����x�v��r�������DR����N_eϜ�b�������j/VVM_�X�X~�������8#�F�1}�楩��M�	��B�Yu�ɯ��@�ڢ�r�����s��6Ͷ_&��AV�Vվ�O�ݴ�k`�٤���)��X��A+��0z�Q�0P��^H1H.;�Ś�"����p�oT������2�,�%���3�p�			uI^�|sx����ŕ݌X��7��'��F��� *q��e/ʟu��$�)))�VK*h���Q�?��P���=|E �kf���[GK����&�oR��î�9⹶�|m7*�a; �J�9��n�z��"�3�/c!5�0-�j�c�®1���U�'{�P_|(5{��x�����r|�Q�[��H}R�A�jj���У�Y؋ч�ɴ�����J_E����+�Ȫ{�v�+@9���2@����^\��e�7_U�u�S�f��Alg�����G]Ǥ�4E�������3�{o��M����-���/%E�wVd5jGzƚ�9��~8,f n�*Z�/�`@�<ذ����	��N~{z��(z�}�<��$�z��>��%u���G���D�ywBi��#˳h�ޑ7�*�ɢ���T�%1�4�ш�׷_W�1�E�lQji#F����?M�R�S�ǡsr~<80p[��Usdl��5��	�7o΁�=V����U�®��8@
|���pK�%&�;�cR��j���w��ܷpʪWG��9�/�R�I�]�w��\4) `ғ).��:LTуY;�F���ր��Y�r%�N	7ܑ��D����<٥�P�i�J����R�Nzw��.�1�ҍ��ߜ�=�j���0�����Ӎ��z��7ڞU!��3Ծ�%�4��I���V1��N�SSt�bdL�F�s�װ�
�7@V�l`4���H77p|~���inV��r��jaYY�P�vE:R\p�����7�2�_�jip�U9�@�Q�� ���yʗs��=<1MN�#���e���<���_W}�ǘ��z���K��&�^"��
��;�Bd����JL��$
9M���὆g��p�n����l �)���t�� u����~�#���Y�E��'�%�PMs�S�u���$"b��tB��::�Vۘ��y��Wu��*sU�;��_Q�ٳU8�S���_�3?�:�LQ�w���f��[-�e����p�ˢ?�zs�?�	��kz<�vXR �jW��X����Z�=,--]�,v9�Ϫ������FZi��S�kԕ������i��8x�*�FOhb;o-�荎���f��	��n�7�X�Fu��,])J�)V��i:��{ї1��|�}:��f��$ <a:�͌n��h�Ff�"����~�L����d�+���`���@���T7��|H=7��ֹ��@����`���v��~&��{���Ily�7hSGً�b?K�u*7�js��b��ʷ��LMm�?�WP�'�����`���\�H�Rǟ�|x���69�J�a�E���u:��1��Rq�g}f��xy�F��ӷ������<W�����JJJ P8o#[�D���W:�=]j[H4���˫��
$��������:ӏ����s#�1P��!���/�6��y�X��D��u=��_���IUu�Zf��?�����F��z��X$2ڼ��쨸%b@^��V����*ւ3x���nP��Ou:�
���[�RǨjh��yN��@��Z���߳,��X���c;���*�?�:Ψ������*�������3F$sq���F&�@t�kfM(�*�s_�m0�ݏ�`���s��jȔ^���R�JEm?[����8���7��j�"��6,��!"�6ߊ�.�Gg���_�ڂ������kX� ii�$w�b������"OfpWW���&�}S��Q����,�������H����R9�r!�t�,Q�bH�!:�����K�M��4Īz�e����7������\G;��ҪY�B/�#p����jq!*-�z����΋H8�z3D��Xu���Q�+.޿n��X��
�°v��2hG���2��:6GT�$��n�����	�?;��r?F�1s�>� �Pr��9���V��'n*� �*����B��į�Ƴ~v��I��N��d��}�� ����G�m�L�x�* O����yI��⃃�$q?�1�}dP��F7,�=2��M5��BHKKwTG�,'�X*_*�qŸ��1��ҟ3/�S^޹�BJ���փb�'Rֲ[q�ס�Ii"���IjY�������@��2)g����mR��i���V�3�)F���ƿŢ?����,�8]�V��}����_D��[��n(����
W�\Q56������]�Z���� �*�F��&Ʉ�Hj�A�՚͞�p��>�ȵ�-|�U���>�R����NV�x��MC��ڳ0-~B\��Q3�5�a�3����-���O4��������^�"��g�* 8��{o��:P9������9�'��P0�>��n���7��8�I�[���5���W%vd� ��Y*�]�d�p�ٗ�R$�;=lr�1�c�3��d�&�	St!�@�/J[�#8���N�#��aSX���R�1�4"%$����OM^~��%���(Ak��H�R�=s�,�B��'���U��
RT�}y@�)h+�3�%�G���ְ�Cw�R��H���uy��؟���+�%��F^�y�;���:82ZVB�����{�}�M�q�}����{X��ֽ%�����ǋ�~��C^Z�݃��j<��	L��$��D:eV�}ܶ�5�E J"�I�A�w�GG�	����|��̌ ��:���)R�ݳ*jB`��G��!�<�Yt[2���S�i���`'/x���Ȳ�����Y�6#�FD\H�O�DO��r	=��Ron�J(:���l/^�fXXs?��%�mK��>-�P=aa
��)
/�g\��=��猈��X����)�̥�T_3��{{;�j�C+�-�QD�����*bɘ{W��� ʦ��V,�:�{1ϛ:��`s<!T0�N��{���A���¢W�����2̤g�E�$&���� �;���F���nX�F�'�7�8���y+�{`o��?0��Ŧ7�����uMG|�/2�NǾ/!y������F��Gg�, `4��(e�Ȯ���~g��͛;�U����6��<Ɵl:���T֑���S��H�x�9n�iX��JB�ɵ�E#R����}[! �v�--�ka�,�AJ\@��4$�C�����F����`QN��M���{���}11I��XQ5�Ð�^i W@�����:�����	��?�ݺn�a���rcnsӢ;:v��4����� #u:|�Y�H��I:Ea�7�5�K�|9��?(�2���,1J�J�#sy��,�@;i���g����6a7��<)N��bc��m��|A1׽�=��%0��,����qS�
;f4��:(����Q��=7b�M��M�s��ْ�J�r�g�6�y�=��R�6W}�ً_�זҎ��j�g�rr��{��AY�n#�N��wfj+�xn�1w]G�*�])�%O2饙�Z'�#��RO�_K,�?Ο����Z0yJ�3`�`6a����R���8&S� �T	�1��מ$�؉+	g!"���Az;�{[:��
׊ .�.�djsK�b�O��I<�6w�e�1&-q1�|.������"��E>G�g'�5�^��]�����q.M�mA� 
ԕ�'�O����s���>�2|����0pq���^&��(�����9��T�Qq_�V���ͳZ^�W���(�]����lu_{���T9���mC:��� LP�F>��ԸH��W����RP�i�RJ�^�tD�����o`7��0�Ŷ�`���i+�\٦�Ŗ����DT�"J�#��g�v
��~
FЬ��SO�7���i:z�'�����σn �-Q�L�/�UX�b�M>I�)F�m׎L�@)���N��{��(m�=�7��0������ �����{[���^�!����8����1�u���Z�!�J��׵�w�&�.bfo�:��ڂ����jĕH�x�td_�
�����\C}i`�D�Z
˘#n,��w�|+PE�"W��N�R�>a�o�:c ys�J��	����M��/A/ ���6�p�0JZ�>��H?	a,���hGy��N�c9B����W����>��QSˎ�ᘖ'�k�r�"��b ��Ɍf�E�޷`g�O�*�>z�LN؛RIhOY�f8޼=_%��V�����gw�<l1IÇA���#�=4l T�K�3)x̲�N��x���[�;�� 4w�v��Pg�$���:S��8�֍�ⲴB,�)�_K�Ư ]W��>/߭���aT�l��h{�9��]�|s�5��Զ�������Q�D��a2�}2�{#�8��a���Jwf��t�Xa̵c��X]Yi0x����M􈾰"���L�~��!X=��H���>ث��8���NO׎�iG��ζ�s��lz�~t��hO�q�x�dro�/#��c�|��v,vҋ�t�"�)��~�ˡ�co�~;@3M�"�2�pp]��wg�Z~]�[fs�m@�%S��Α�^� ;�p��ώ�7������H4]����O�*��OL���GKs�zp�PΦ��r_�����ѿ�H���h9����t;�ݏ�5�֚5��?N��Z,,�;�Y����`�A��`Tb��s���P(rr�H^ӹ��'��G���Ҍ����������!��	����|��}��[�Ǽ�ϭ���yr��/��S�g�hٙ���G��,D����x97D�r���9�h�R@����ʶ���D���d*�A���P�	�Ԫ�Ō;�J��NX��Jk��.h��Ѹ��G�4^�[SEWhK�ۨ�E�����Z��C���	jg��% ��46[�����="�(%M";�,��t�{��6�%��ԛ�
�Z�����SIS�� ;1u~n��L������|���v|�qYHmjL����c�yۥ�85�X���Ό�ω_��ƕ]�K����E��b�9B@��It�`�!J�3+�Z�٪���:��vr{=2�[_�}�gjUE&v��7=���`ԯ��Sw���m����5:��2�syQ`�@	.��چ�	�5b�S���|,.���dRn8�t����7T2�"�}lKM"�j�wR8h�ݜ�v��w�f|7������
�v�M� q�!C�ȦT�;G$�͞,�V6�g�xVV�B�����i��k�͡����- �p��=B�Q��mG�>�S�F���8-t=������q������Fjq�B&����=|�X{B��B;��C�(�v��L���]����Px�������R�/�:Bh��N���4��	B���|0`�<���-��p0����C��T���gU�_Y�8�T�[�GM��	� �q�5��R��e3�f�p�r0��K4�Mҝi��B�p(N#�6+���?:3J.���'�m�&x�`p"�`VW%�,n&oຑ&h��2��_v� ���sOXv~a�G�����P:26��[�c��>_��aQ�]��_2��T�`�iS �O�x�����ҥ�Xuf��[�뙢u�k�@@þ�����χ=��)S�Į��N��>z�ZQP$-7}���Hu�hB)v���_]C� �Hi.7��/T.�����7
*��{cWυ;w0�'����<��+�R�Z����+�=�7����Q"|'� )�Y��O�(�2М��3}����-ο{��N]'�=C���)�.H$m}��5U��k�N��G붎�W#:>Ɍ��~_��͸xo/�ģd� k�bu�F��&T��Os�2Q ��r���`тO���������
�6_�2K�bK�=nu�2���S�)�̣�P�N;���q��Tf��f��Ju57=�=�Z*  ���% �:8Hae<;�gt�&�������Ӯ�m��-2�����K�꣭"�Ƅ\�~�=)��N����+
��kt��� g�������_��֥�рI��H����V��t�c[���XQ��{>�r��so���"N{���A�~��`sZ�Gc���9+'��Wq{�p˵��⪤�l٫�?u����Rlp���R-�WC��.���gD�BnĲA!.��8"�ԶP��紜�c�
��k:L=�m2p
v#!�~�Gb�@0pਣ��9m)X����Խ��}Z�'7~eC�XD��N`�f�J�R�bRե�����d[�=�cj�<��sJ-Z p0m���[U��:��>5��Fn(~���s����(b�/�7�Yv�����ʆN�7}dŀ ��'��&��t1���́{��7�O`���ut��ć�ڤ�⯕���$��$��e�[�6Q�C 7v��h#�YR����C�X���J�^��[)'~��`q�閦�����$��qI�� �x��O6�l��ޞ��&����������$$P׭�rT�A���������£tܘ�OTٰ�h]�SQX�h_�k+�ŅJw%g��S��LAFe��j�L��r���;2+��_��������S[?�e�Jkz���z'� hd������?Ƅ	��6Oe�i�uVy����p�KPVZ:������5IB�(5�ٹ��X�]�Q,��O��82YC-�k�R�&�dɲ>�N2X�{��/eq�I��&��b�ٙ�ڮ����d��p/��)��1��Ȏ5���]j���������'pW�#�~�)m'��]s��QLg2$��E[D�Ţc�. ��'4�<CП~�d��� �$0e����%�P���.���������Z�4U�� v�l�P��y��
�H��zr����F���\��HM��������7����F@L^G𗋙���B�q��f���x]��1ѷ�������|*"%�	]�6�	�K�"�G�:n�$.m0F$�ߕ�4�r��'��a�����<ap	��M���B�>����!���n����g��om���6�o��c�=�u��ZХ���vR��m}��:���J�6��z{gG��
/r��IК�C��;�܇G'_��H]z:֑��}�"it�fi���w�)�=c7(K��>���E%�jLU�)j''��Lw:ĭ��`06f��A/����N����V�)���)+�-�$7LoK��>�~a�BWs�=zR����✱i�
Qy����[�u�u�j�U�+��ؘ����j�|?�T�p�}_"��~}���yqY�O5;썍G�_ŷ�Z�y��˥C�"���Љ\���&L�jXeǼ��� Z�e��O%��ً�)���4]M܄ogz��2��*��B^F�Q�GU���f&>y.;�F*nM=��8*j���\b��ܸ�`}�[%��M�K��*�����1m�0m��O��ѓ���;�:A����g9�����d:��G�� r�`�����]�[�4��U�������ħ.=>%*�R|lF�c2k�I1e(�`�Øۡ,O����W7��Kc+��BK�@6|�����c���d���o�Ag����^ǹ�y_=Q�Α�m�)��eC�=��rx��V@��'Y�����=GW���,]�/�Ƙ)�����t]�`;��<_��|��_G�h��B[=�/��8�y�h��ܢ��W�uq��<�R�*�}���c�$+�g�͸V�0�@�N�shDau\�6�8�
�?#fD���0ߋ�6�Rs��H�D΅*�T��G¼4��s���rBZ���ߍ)N�Q�ׇ�ifq�35Z(g(S�K�LT:p�P<��wh���ܨ������҅��,��{�s�������:�|b��YxOJG�l^���Pl'#�}�(�t�J_!n6�-��Қ]�0���Ⱥ`y�x��v�^����ʗm+�.�1b�2����������Q��K��ڋ?�j![?R���ew�/���s�q�,�e��-hZs�s~�*�t-��1�Â���O=�T{�|���7ښ���sA�7U�G�7y9�����:��}�}��8�f��3<j��ZE5���~-N��w�����&��$#s,[�,W�d��9!�/�7݊��&E�a��JM�Mff��V�q��R�X���骩Ň� ��\1O�Ǆ[nI�g��y�L�[��X�Y!��+����Ww�����tT��������u��s�Q��x��u�T��A4H�3�Y�(��=��o%l����_����<%�.nC����w��h"�B����t��۫�dl��\e�f��d�����ܙ�����sZ�=0����[�����|o2>T0�M��;��&�����M��F�<���[�,�7�K��Vo�U�2�|�]����l-֛��BP{�����ׅ��9y����uܺ���6wfz�)n�efw�Ruzmơ�i�Vj�t�` R�jd�~�:a��D>���O	�ͮ�3���Z�c�o�������ش�%ZD�!�y65�(ҙf;�,��r�����J��Ρ"k_^�k���F���u��빋~��s}�M�"q��r��	���M��-ɏTފ��Kb�\��IU!�������O�G�z_�����J�Z�V�!S��	`r8�r�t���&��>���Q�ⵆ1;H7�@��*�w��S?Ǩ�����I"{:����Uu�f1}�R�tM�j=�S3�Fh����yi�RC���K�};Aoܺ<|!����
��N���p)#%�ӰS|�IpפU'�z�;]�I���f�XEo���f���W��!N����$���m�;2q�,�!|o\z_0��k�>��c�tLR�����̠�U���E�xawi`~S����T�Db��X�]�Ӽ	Y��v��L�:wX���mw-���dɱCNQ�� 4�(��h�.�ޠL�W���O���z�+R�u����ǖN.!��"-����"l2�e�5����B��E����ۼ�k��-�G��+ۡ��9�:2+�3Sc��j�*�)�ft?ģq�|Ol�[2�on��߂���x�@�K4<��1��=z�l2~''��
����@�J����cv�o*^��7~��ϻ�8K=RE��z�+(�XN\�@�ȷD�^�]��E�O$�8χ��I���;@D���y�����4������u�e�8�8�xꕯ�u5��\����Z�1��q���\�-��Y`�-eZ2(U}����]$��~lU��ܑ���7�wN�F;�9�p�7L]���<=�l��3�J�8Y��Y%�)_@�v�'Ox�?x�b��{����c����P�t$��]���ꜚ��T\?kI��]�zv�m�E�<��T�P8�dd&�^r�` �χ���2M���6Ui���[�n���R6�e�ܓ�e�Þ�A��'�L	M���$h��m��l�D�_��;Z�q���\ȳ�͍g���A3ߏ|6��A��Oğ3_�;�n��IcT��a�k�:�C�a?���YxkY�����.����Է��*/����P,��p�w�n���TBq*�~�ˤ7��c���C�Zf)�)r�����g����i���{!��a{�Ÿl���E�v͕)��~8����Q6��7��>��j��IO�}�(��u��|�Q��wo�Qu �(��xu��lvi���2���������q/BϕV�O�#�� R-S3C+H�~�U	�X���3QT#��Z�P���������>�"؞h��V����n �R���$�[�����:�����92���yC"M��%�9C9U�rC ��ڹ��a�9�4�lyk� N�qB6W�	�'�E�x޹zMn���P�B�*+�k�ە�P$�(�i���2�>5iN��ԟ�"�t�9U���u�"��r v\�G�(���[cv��w,R\!N'�z]{� #ڸ�n}�V�Q�33��f�����S�.elќo2>`�e�����ə����RTh��Y#3���
 g@���D�l
�55���s�"j��(�t�՟��4�ҵ�����V���e��MIyZ|�SSn��>	H8��2�� �z��sv5^`+����E�}S.]��N8{��Tǖۃ17m&�1��Ѐ��������}����+i�d!t���A�[���?v����[���,�x>�w�x�OOƪ��|t���b@yRrI6�~�c��n�M��- W=��� �ql\y>�T(�X���R��zZUV|zAY֮D{�E-g�*� g%
2_9|�"MB1`�'87ѓ��:���:bn5�Ftճ.%���f���Dd(�m1��^a^S�F���?�a6���i���z���X7-_wo?�2Ά���<@���]����y������W�b@���s��K�+�@U`[�c�D��,P��z��&%L-o�>6Z�8}����Yf�����7|�|`K���Y ��o�1���Qr�9�/b�2<�۲?��_��rQTn��d�o��3��`���ӌ�ƲJdQ �n�(y�؄�?9���V�y8��RiCz>�#�3�����?����%Z�#���8��3*��i
xm�zz�P��� �z�I�j���Wj	-1$*+V~�����4���td�鸺�t����1�V��eX�@��^e�t��@1LX̨[~{�O�q���p�0Bw]�����IoojT�B�ғ��B~�?\�\����q�뫔�C�j���'Q�M���1�;x}��w瓹��e/dEռ�T��i��D�W+w�P����µ��־B���,m�^�McEf>ÏG/����� �LjX�@ؓ���	ݚ~���5����74R"��K�ȕ;ǚ�ɞ�һ:�7܀��ܲ����}�h�S������s��ϱ(;��\R��̉Afi7�(������W��(�D�5<����Ss�0����ׅL��е���q�a�����7&�.T�]z�h �p�o�-�j������D,�7��(W�JΟ�c��q�]��*�z${z���؆���DI!Sۀ�䂣��i~f��7
�K�=�}r�����e�9�P�'%�R�Yke�ZvCg&�4.�-�\����������9x�J�e�Y����q@aV� �+!T[�TX�e+ߜ̯}���2K* �����ȟ�UtO�8��ת��T��Z�{Cwé�F�.�zj�b� �y�����G����v��������H��u�-���/B4��|�4|�G���B�+0C����vQ6����ܗe`Wy���2t��?�"���ѫ��,0�|gz*�^��p�D�`r�nJ88���:�` �T�~lu��L�[B�1�D�!ܪ�聽��������3v�R��+~��4��9�;?�3+]&x����
2j@> 
:�~S 9���rC��n�K�q�	#9�S9n��t�XT0Sm7�%��I�i�<�y|��$��H�)��b���Xh�0�ve���cO�a��g��#&5!�6M����k4��Mo[�$E8{7���AӢҏ��3_h��H���s|@��[u��@�����Pj�K�P��Gi�60�}k,�k`�pϮ~{_�����{�7�U!&6��գ�' ^���%'�&������#9`au���Y���$Ǜq����o��4�?'(�L6^�Q�sa���A����3�d��������[�Y�To�,�`׆&���ũ0�2S~����B�=E �{���>�"|����IOh��,om����|x��l.��uG��t�R9S���N��
i
�%�
K<�D�ߡ����RQJϷ�i���3�=Fv���'��?v�̣�Ŭ��y�\��u{�>�(u���l|�+��P`|hݨ9:���mg��E<l��� ��kM�%',%�ׇ�By^r��-L�%���j�dʅ9�?�7���'����qrC=�+)���J���+���N۰@sE�F�/�<�ƗF�[}�����Y��W78e���`��T��-�,��6�&�󺺻 	eKT����U�ކ��N7.t>N�l+*Y��q�1V��$d靰�;���i/k0�����[l^D���C���۠A�gN�_�F�e��Z�h�a��p�T!�e�	��E�D�UF?��&�B5�XPє2
����8�k��?:�@w%{L��W75�@��q��?��w�\ 4��Jǂ�-yU���#����	���\1��"q���d����2-� [Q_cL�2u{[�t�����Dq�$�q$A2�!��vOO�r�gn�L���������5��������cŃR=�F����?��I�ī4�B�c ^��4�A� Ei���>��)�Қ퐖QQ���W0ƷZ�������M������� f�h[b��m%����w�M�k������}zk�8��[I��k���W�c�r�2l@�F�q��w/8v�������X&�`�@���3q'��9ҍ������bV��l��O��oё܈},qP�f�!�H0��\��ߦ-w�Fh�)��Ҩ\��F0�D �g3.3�.F�O{pyp}�	СʈK�#�~Ы˒s���vr9ic���Q�>פ�f+���9�Ԫ����b��br ���<;<C=�a\#�u��|${�5ɽ��B�AM�.��J���+ufz�\�t�u0�~�"�>��<_m�^j�g�2�ؑ�V �V�4�䗒�k���Ȏ�sPjzZ���%P�ގh�
��j�v����{|/�w۩����I���k�ۄ�����e5  .�s?���7�7����L�`�E�E)�I��r��?2򓥥^���.�\�ξp��x��FO����o0~��ܛ��[1��t�#1�Bؑj5 z����V����2.��e��=���i��.��%ߟ�7.@��RN����(E8�.�+&"r�r�zDg��u�Nl$��,�"L�Ƶ�� �i�k/��1�=2฼�T��O��ڃ��%|z�J9���a�K��7�Ζ�f��gh���7�Mí(��|��A.o���8%��u�EMN^#d�ϣ���=:��6ۅ��6;��p�P�n?���G��S��π��6U�9�P�8h�� ����3&ʧ_��lS��c�*�܍��;�]���	���No<8���3�1��l<�_�z����C������A�69�8[�@����HΪEŪ��ӡ��	�_�Ϭ�>u�sg��[�*@w�v?��*�^������E}"�6md\ɓ��=t�^�B:��=S�gvl�#c}-�^1���@�����W�J���jt�Zq��U��f_��s�画#.�l�V��G*���?UC��z0d��ǖb�
���&����w�H���u����pכ�~�o���	�q]�,�麲��f2�T|����.����غs����-���*����������m���U���*i�Ο���LD��T������ƌᬐ>�>�q7Ap�(�A�P�/����5p|9��o]8��eo7����SK`OI�1S(5��v����1��2���1D�4����� �.�}|:�_c�e�_�H7����DS�� ����2�������'����pՅ=�ٷW(y߼,5}�ܴ#l��cӄ������<+��~k�>�w����[���&�F����'3�����	y��`��&�f`�P	0D��?4�]
۸��eV=��uWOψ��4cu��X���~�NeނB��h`����� A��ϩ��j*i���x);�;�G�=��OD=P���uk�{�����Ï�;B� $��n���ҍ�ޖ)���G����o�@-[�A�r�����A�X{=%}����1����ܧ�%~~����3ݞ�B�V@� ��Y9��Z���[��y�#Ȩ����N��Z�4�s�"�n�T,�J���6����| %�3?���3��6$'����[�?29���B;1�&�j�C\�Ř�eu���w	;�6uJW(�}t�Do�`��آ�@}mN�BSq#���h�W��������N���/�\Ɋ���&}�,
J�F�5�-���9e�ۃ�/%%�ڴ����u������r�dM��/��m�ɭ�o�c���N�Ų9���+s+� ��{�Z��e��	)������p�v6��񁘦i{�?�XaIy�||||�!Atӯ *�vR�{Un��Fb�j���%������ /*�@+��Q��An�V&��؟���MT��&��"dk���XE�����{�a��/�����.�Z��TؠS��,ڔUb����ӜN��2�ku�:ES�̗׭5.+jOӕ%+�9,����3O4fOv������n]X�������U�w{���nt2ڬ�9	�0"@X�b��Ւ
~��W����6�!���3��O�ه��v�{�k�8����8�5����:�^99\G~�r㦮����S�2$�W7d�� ?�{�ӈ��?�O�H���5��,��!�*��ھ>*b!�((�t+
�4H��t���) !���]C����C�4CJ�P߽�}�7k�d-�{��g�o�i�,)-��ӄm�6V�Gr��ű�1�\ץ����ˆ��t�	9\.-� |2�����/J��?Q�d�#�����F��%��PJI,]<<&�x��[��-�r�������<��T!)�/M,u���	&Su	�6�QQII	f���6{�Nɉ�ބS!!������WU������9sٙ	K�kT�b�#˻��?{��o���Ԝ�ڌ���2?�
�	U�W������å��=��:�����sLn L�['����c��ʋ�x��"t�W�$CG�1����K�t��d��ڋ�ل��\�c�t�YL򠨐\�G�e�V��� Ҥ7�����T�ׯ_�l�h��#�ֺř��#���w��]c�� ��wV�����b^�xKP�j��pX$�����a	X�-�&{�uttȫ������
�{�U�.��Ω�B.�:W?��� )�U�;�LH�����n������"�D.o,�Ǻ�K��b��x����m�������}�a4r���e�8���Q�3_����#Li�c���=�GA��ʤ�Ä���D������g��8y� T�mVy��A7k�,�h�H�@�\��8��-�O���:%�iJ�KY���?Rz�\R�|�������o���A�F^OO#�?l��l�?'���SW�"�B�����{kj��8?�Қ���>	$K8�0�ak�AW�?T�(���@��
שj��53�<����"�����ic*:�˘h7����5ȌX��tu#��q�g� ��[c�v�kGB�э�+ Ϯ�� `7�m (7dTPR�\ޡeb��t�c���V��m��~�
�j�[�������������/�C|-��F�{0�
hl�B���I7͝�o�J�G���Փ�<�t�:�d���d�C��F���E�W�с3`� ���e"��R��


FM�w����\��&4�{� ������(��	G�9��7Y�L�9X��+�;ou�)Z�g��	��c����b|<P2��f����r��랍]�ȃc�q\2l�����4~PE	�!���[�>���:U�g��ʩU�8��־���yю�N]9�)��%%�bS��B��L�bؖ�O�f6�#�5��]A����  ��_
m%8�?V�Ee�R�K�&s@�_����Zk�b��Y��e���|�� ���%Ă�Ab�Y�k��(��"���z��66#X�.�I�j�D����A�V�t;/]e��jf 2��W�O�X1���g4����BC�?9X�L���_��7�A���;j��}�V��hpQ�,��4���aؘ�����JL�7񦚈W/�|�19��p��W�G��E�se�sE�z/bSJ�I�UrdH5ૻ"�����������!UJK���Y�>��$%�dʒ��!Zsω��Yc!}q�F�&�4�2�i��PI}�G�l�� �)����.W�Gݙa�)�$���U�E<�gv�|�k����x�����k6㷽^�c�,1ZIz@��u�����?���I�(��M�ҍ�q0&XA�|'�9lrA�{A�S�ESf��u�rʞ٦k�����9/(h:$K;���4�v|�Ǧ�� j�n��j�~pϮ�v�Nx(��P�NjǴ����7���dH���ތc���eXD���a���%`>ǈ&g�\�LI�V�\E�N($�}K%�_�ve����/��Y�}�1p�w3䤸(�N��qW��^��j��o�p̌���R�8_�[� ���!\��Y�x6F9��Ny���Ck��ё2mq��m�����0���눿��n�װ�����7&{e[#��}m\!�}|�l|��0��8�ɘ��)߾}�<�oZ�9����Om� `a-�H'���h	��ڰ�w�b[�宅�)T��P<����-6��x���o����pJ�C�S�5u�=Z�1��Y�cS�b)~A��I�lR2Q�t��(L�s�1�n]}x> ��{R#���Nq���_	�N���Iå���-�R� ���@��4�ZmQ���o��]�^���L������gP�	�I�������g�N��4��f�ډ�F�YhK��‿��|aE�5	�W��[�L>-g��1p1v����@���,@:��$�ϡ���i<��N*@����Xn{����WyUb^�%��'�k����T�����w���q�1e.(SӃ��>�V#��m�FX� ����( ��ץ�����k�3���0�l�+y��N��Ǽ!RB���2$yt��&W�cQ�KRv@��P�t婤����d����!��f�q+Y�/�f�j�?�[a�r�|ߢ����e_7��;�Ⱥ�����l���zx��>��c��<�����,���Q��X��x���[�P�f�L�f*�ƈ�Hjo�p�Ou�??�m).�@�ڻ�ʥ9�i�Ke�쉧�,���OKG�oVU	�6��2����@[�9� ��M4�WR1
ݺ��㟔E���䑪�7�&��.��ifw��^sK&؃:�v���F�f��5G��8t�7���$�(d�w�\EBİ��8N��`}�U��&����]�o	�~6�9R�a)�B�1���6@�;���K�\�;h�'D!�ҏS�\�y�Vm\��r� >���N��BY߫��V<��e6,ُ�t���bc�O�]pDiY��Sѥ�`uBL��9s'��z���|�W�Z��dE S-\����`.z7'q���$T�n�������kre�S�C�,���a"��|NmIrc� 7�v���QF�J���+�4�L��~)]ŗ��$;��9�qX��ɤ٢#�r�� 8���$�\Y@�x�� � x�����6�����j�IJ������S)��o��4&؂��;�����-D���,�OF�[x�dd���)4��α��$X� �@<�Dv��,3��V{��nػ�`��V��ɉj�\��s�\ik�r��n�L<��<���NI0���%_���~i�KC�3۸1�ы�����l��Lށ��Y�U��Ԙh����ޤ�tr��&�:'Sg��1�-��Ҝ0�MKή�7��t����d��X_1=����9��[h�a|�MYW	�S"�2Dn/�Ǜ9�2�+��2��ItD�����%�a�9�u����p�I�y3J�0�<��*�.N�|�9i��}��Y{Ԅ�@�yZ��:X�Y��n��e�-�z3*
�fxg�����:��0��	���yq�l����(ꍏ'� �p�$��2�g-�Ӄ[�km��0��$+6��)?�;u��b�"��?+�D��D��K~6y�B�Y��ȑ�W���cW�pm�`��>c�A��7EQ����-���f�����$��6Q�`
�� �H;y23(by�RLǈ}M�}����4%b��O�N͙E9��e#�%N>�e25`!a�Y��[��x���:�b
���5܍��|��=�"�[!^��{$�����	���zҨ�W���#����wR��(�X6mֲU�����{����~�P�1�r��{�����I$P�(�8���n@����2���9���T��O� s�m7���Erp������Bӈ�ΰ�&e��!�C �m�R�%��7'�Ʋ!T,k���v� �3�¤����ӏ<jLآ�[.�o�A~M��	�0R��8x�&� �f�P�k,��Ǖ~�X+��(�x�w��j�2�,{ӊ/����	�]�O�<��fШV�i Ɨj^0Z�5��a!�w�"��G]j�������O���BT�z;
�R�;8dU%����ZX�KBG�b��
�ȭ&�s���|��;D�櫤�/:�R.`��oQ��"
 h��>/3���~[_qg��Lz���E6pYI��(��$���kvF]R���=�!
�Y�uhΧ�����ۧF�8�C=u�S��Aۙ��)�~ݒ�3jW�γ�"箸�.����թM��l'���dn$�A�6�7��x�,��ߔx�c�Wn�esJǆ�q�Q�U84k�)0�����5�z��xy٢� u�&yו
�O:/�U2����)4\�Q:A�qJ�����
%c�$lt��<�v��
Q�{�����sBJ�._���N1�ϙL}��|�S�{Kv�K�O��;o��L�S��ce�W�v=�*�WZ�x���0�e�����u/���]ƍgf3Tl��q��JГ"������ |+�J�����G=�D�J��]Ж����rQ�N���Ǫ�1��\"?�2�۷s5����`�(���C�<\�s����Gtk�G6W	��S�މ��/1^�zn�T�9{�OJ�; ��播�����[%;�J~%�H�������_�8�?���O/[���/Č���};����yd;Dݺ|m�V��s_}Q/ J�$o���FL����v�u��Hߦ�6=��͞xr�q�i�%��^w���qg-� *�J��#m�R��
]�RZm5/u��ƍa�"��\�69��so �v��-�z#���FCArb���ˡ�A2�u�v�Y�lʫ)��q��.��t\jH(��9��B��̒��Fp!�ʗ��>���y�)i�IՉ�=�J�(jW�<k��y�x~�C�A o�#FUS�i���H�w&[m%^Otp: )1���=6(yS��>�SO�*4�f;v�Xa<�
�j%wu  (|����!�/�mY��av�b��-4���a�E?��	�3�V 3�+|s=���o��S����8�y>��u��?��'2�+��;?c0����>�*�ǝo��M���$4-1�_�e�·���W��c"ް�*4�5�Ù��x*>�F�x���C�?�9�c�k �|�2��s�t���-^_3U���"������`K��'Y1Sr�󛞌�7ӒΩ���a��-$���T<�'C�Y,7uH{Ow(Z}%���L��u���d��s%�%���k�7/��ci4M���C�&?��k�D�V�}"�'�^Ae,b|�n��o���;p_>8:�\$��d�H�Bߐ��Ҝ/�=unD���V9�x��qu<.���l0��/!��TQN���*�Tn�#�ψ#d-aɜ(�N�K���N	�~|�����*R<"�N�OW�q�~s1/�\���(f�qX�&��X�=���O��ݝ��K�"'.�K���G��7wt�Cm��u�ׄvl��YXXX��7����nQ`y�$�05���� �ɑ��:��U�䱙Gl^������5�d�X�7�V�&�3 �uW�b/�^�6J�G��.Jp��G�cL��@<ϴ��o�ב{��S���ף}���U�M�����zg.u%��=�f ĩV�Q";T�12."T�o.k|���Kc-�"ԭ=0���*"�!G��+�ǯxx�K�^{�e�k{$�8~=������������ܕ��)K�&�z��+o�\(�}���,��S3灁�A�޼���8��jc����j�3λ���3� G���9�]21Ͳ�KpX���E� �q�:��Lҿ!:a�>.ǠDB��1.�aP yv����ʀ�y�~l�]f���������O������`uJ��f��^���˻	�/O"��}��ƻ�Qi��V�ջ�.�68{�%�8��-*�"+�\�,+:`�vS���8�dN�(ބIv�)LI��9���'^���~����@�� �Аgs��t{N��x�{�U�]��5_@�����f�$��E������R�z�-��Q���֥�ƺ�f�;�Ā�In�B=W�#͛��rpm�����ȇ'�dp�Ro��5�v��z�P�5G<��^|a6�W��׺�~���E>�Y4��1U� p��VeU�bY6���
��to��iU��
��s�����@_�9�I�9!LE�$)ve>��&v����˨���p*	�$�� ��x-�n+�@��݊���Y�Vx����/���}��Q�'nO�l�7��jG.�h�)?5��V"��ƣ�|2�x�����_p�N�ȓ���ol���~�3Q�#�2yp���:CN�% EN����7E&��+��f�fP�r�Y�+���_��"C.��T�T�+̡�/?�2�Bk���S�פ��pr�h�:6y�ytt����H�����eء����D�ź*�3��_%�+!����4�aA�o�&�
c}<x~q�qP��p���}�/�~YfbTi�m���~���qR���,ߵ.n�����[��ѱD�]4��)�ٞ<N()Y�[i�yc�P,#�k���C��cr�nI��� Z�*�N�C���;ȡ+�緈ZZ�UY֜���
��!\�R�����P���.cS�~?*0Vn2��_9�LDp3��'��H�QGw����7�H�6���)|���7L��ll45�mqQ)��gdy(��H��N�Fp���&�R��!�7$n��H@��X�L�S֔���!7�Oo������!�?�o�o�c3�������d��3����a��`?}���e��>�=66x���H�p�?{�HK�����l��������Љ�ZX8�{̢�U�������S33���gQp��d�G��z�ផ�ryv�#�z|�OP�^'�s��o��;m{ݘS��.c8���ɢ'��mć0��hNB,��U2��*^!W�d����):U��ED�,!h��}��.ԡFZ��T#�ñݏRV��L��u�Y�yëJr8cZ�V�e�45���B���*��S�9wc�L����"a4թ�t����p:������5;#�߽".�|qw�UZ#�&iYvS�.����l)m{��Y������_�b�^Φ.�L��r꾃�ѿtΊ���]�R%ا�CGO�)�姨+�)+g�uFа��`��m��Lq8�w#��I$b��Չ;%���+�{ꃛF�w�a���J�����/����X��Ka�������R�11��'t#���(g��� ����?+�b�D��������/��#Ww�ɞ��1}ݯ����@q�֚0��L��oI���N���EF�U���b��l�b{��zm�!d�w�Y9��Q�*��09���턜�z���?��e���Ӱ�{�x��w�f�7��l�ě\5�n\*e��\�VC=t�ed|drA?-S |ٰT42�@��7������|�ω���2Fv�d�uL�捂�g��dvaAd��G�.}�l`��+	���vi5=�5½|���B�է,m��td����^�%�/S�ꨕ�w�%�u�@Q9�D��@^�Y�N�)��x&{��Ң�U6�1��}�3Ipd$^�5�Ϊeo�1��h5���INJJJh9Zi!��s����;��]�p�4"v��<@���[����z+�8auf�.���j�9�;ZK��Iy�^5�c��t7�zh3��;� 2U�+���}꣐��=�;�б�,���)7F���j|�H�Q�q��\�̾b�y0dҺ��h����}|�$�`,������b/���(���(��4�Yr>���'טkvK��+gn���ǝSN]�h����^Y����.�q˗G��\�$%%�^���p$��TY��5���_�GY6��X�<=���{���O"�� �51����lш���r��7jrI� d4�x2�FX�Iq�[��$}�)L��x~+��,�o��Q�O�t(���������`��Y�϶�t����m|�9'&�4��Th�3�g6�
�z�br��*g,!6������^y�=��c�/XU�kh�sc�cYZ^��{��#z%G��.���ԓ�Dn��zG'ώ�*�8�]�4��B�=��jF�o�6���EqL��,���\�OINV%,|Nd�b�;���D��R��i�A�֭Ӵ�x�)~m��k
8������J�~��������G�2þg�v�.�s�J�jp?��־dЬ�3��ͷ/PX�2��wٹ�t&��o�4�A�#$k�F�)(�W�Ŧ�t��Wl�;Hֿu\�����v,�Ȅ�Z�ڐ���Ͻ��������w��(]��#	a�΢9��nL�g�,O�R
�U~��^|k�^Y����wcvn��Z����Z���R�V��q�ꧬ|�?Ku���zz��1�}��`?e�|��:NK���N�gAX�cwm�_�jNmQ�"9�i��z<���,3>�鯬98��"9��;8�x���ĕ3H�۟^���XASM�*6z�;ȍD<���&ώ.��v�K�F|6���nF1�C�A�}�A�+���7�p����T��UIX�6��.Q��.��a�g����r8��.+��nR�1�t��F|J*ۻ�sq��1<c�L"lW���PW��677ˬ�:�"F)� +�&��P��4E��k�+��u�J�$#T���U�K24�e cQ�v���U�]��7����!��Rj���� R����P�9P:GM����Ɨ�}	]�,V�2<����V[�g'7�6�7�j��ؗ�g�1�+:�H�v��+&!�L�~����=�ͤ�Q�r��g̗��j��������E9n��Z�P����8!���=��t4�_^u���"��TK�iU)ZsPB��d�@	�$�\F�KX��f[�"?�S�阱����T��:�3��z��|أ��	�h�������m�+���y@Ġ�Ln�%�����YP[[�U�&'�
��}Bdu���n�V�tj�XʥU��h��6d���,���8�u��Yz��Nu%�9,��cϢ�v�P�<�]�;3�6K��?�N�O���G=_!�6"o
S?�:B�Y��K��qq�0BR���c�� '��ӳ"�$��R� ��N��HKZ5L�K)!v,��J:�K�V5����*d�.�ua�8��|���CC-���B��������
��-� &wY��*\ǳE��~o"��ǰvw���O����w�k�g�-Kv��&9p�]���&����:�f�]Ч\��v\0����⋩�I�1��Մboԝ����ۋ�A�f�>Mɟ��1��GDFf$8P.��6V=Rj �?�fv{�*��7E�S��7<�>���%���I�_;�����-��@&Ջ����՚��V���a��O����6qo���Xq�ԫ�RW�|8Z��e~�NBpP�T���	#?�������e*��������TJ�Nv
S+ ��a�4�*�=��촯�l�Y� [�4��j|�/x�r��_:���ȸ}ÿ$�lѧ%�^� &���pS�G�t!Ŕ��C����@�B���A}1"��-+�g���Jpx���jOA�\�/]�|X|Z5L}p�.�|>v�H�O��X���	����ş�C��hT�j��0~���m[QG3:�g��k���N�V�wV�H;Q�^�X�ˡ-��O2YM�o"�ꁦ��07����S�B*ji�T%#��(���roDڬ���侫�A����8|qqdv�a����H��%1F�B���J_�Q��L���Ys����T^/��y��-�)�
�qy��2�S�%u�k2J0�����$�pO�6��sd���N��Y�!8hҺJ�����hE/X7���T������D�W.@�B;��&~��/kB$�,ȃ���mN!Cp����bӱw����]�
�L0J�b�uR�+����-�t�����u��"a3&�˝�"�2�1����uUn�1���-�!|U�[(�-�L܃/x���w����?�Yes��
��_�d�q�h�ڳ�q���e͓�<i3r���.��k�;W�_5F�����\�w�^�`�}�qE��,�R-՗����g�ǵ�X��J<%g�+�^�l��oVОx�����N�}����4�h�Z
�D�mo��ֳ��k�0q$厖����䢪D�&|�*=$����$�U[�|����n�Y��nv�i?N,&���R٢-n=Zì'y� ~:���$�ls�n��PA�����@�]�� �~�@xK
��r�6���褴�B�>�Sԍ������W$���$Q�m�O����B��%	��9�T\�3{�5;ē�bj�u�8TR�K���o�a��U��S���G�Ʀ �w�@ހ����c	���o�&��,����ܭE�LI�K}�x�x|����I�OIc�Wʫ�YUޘ]-��M�T-��-�r�Y6�����x}�+��dn�:>eo?� �E�ʸ9��*p����T���PX�����ܣ�=��	�j��l³G��c�uEȪ�|�����}{���o���@o�SiơvFm4k��jO�OO�c^:�D0�e477g�!��q���K)�Ԏm��My��j:��l��h�5��f�k&tN�|Vf�$�V��nǠ��ѓS-�՞[�褣��`_M9{� ���
`l0�f�����d���9>�2��$E^��s,�l1�?B5}UZ�\�^b��>��[����k�;���u�4��3�sϤ���>aau;q6��ck��V�E��W:l�e��X���ly}�T �I���G Ϩ��|�`o��a���W^�q=a1���O����8,�2�7o�X�:��+R[NR�v��ұ��Q{���a�&�Xl
��_&�Y�I���ٙ)a��yi3�`�Tp�ʠI�u���r�ol��(�,\��d���*F��v��d&���a4V�q��EA���A�h�i��ā���
w�������F���D%C�n< ��)���y�\$�P��^X���
8�x���>.{�	��ìS�V6[z\��X.�R��Q����)q�r�놃. 'R���֭�H��K�#���ꂂqC~�D��]��`r�#۱ҍ�Ý��5|����S�e�F%Tg&�$)X�:���fj���M���Ig�8��d��� K,�.uĵ�oU���k]c~������2)�f;بx�;^s3�,,�˴��3ȳ^��`c��qYC ��Q��֋{	8*Nf���wm�.�� ӑ�Z�hw��`K�/�37��d�"g{1+����ͪ�j�p����g�<C���}��\ER��5�+l�;�z��0�׈3�e�\�8UK Cs�Tj��S����-I3W�N��o޳6Lw߭��n��ݕa��_�6)���;g���b���)���l�B��\�B��_~���v�b
6��{��jI��`��r��$��@6Lf×G�Sؓ�3�ձ�v��qyvR�V
�*�ļʹl2}a�/C:gTB�ʳ���TM�<�z9R5�إh)��FM������@#%&�W?)��T��J@�&��x��6���k�7��`���t?*����N���� �,$-Rӕ�x�Y�7擔6b'	QQ���q��ޤ[��+J�f�>�LMJ��7�������+G	
 n�YEg8���j4D$�ҪǼC²�3A͆���uX��1�,�V`g��Sg��P�|	�E A@�[�5���a$�����Sžj�7r��[H�$�v����
XE���m7w��� ;N�֕xq"!��܆�z����Ϫ5#y�����4���� �G����2�ֺ���JO�j��"L����|���½��ŝջ#.E
����0 ���\��j�>4�@*��y��g:>'���d�W��m{�w�s�ԛl|���H�u��<�9`ᴕ�ZӾ�HT����aJ��vNbib��(� 	"�߄s�l��� �c�Y���闳�L�;�(��f�(T*l8q�x��g`���LT��\�!�׻��+((��D�A��^�����))��-��о��7��E�:7�;���P�7d7�ش��������^m`M��L.��`
�UGc�.?[��HU�'|���J�7^����C

H�[�Ei�
c�t�Q�*��(*�嫼������f\�����&B,փ?�7<rr���|��4�̶s�yI��0'���0!q��[˱Y%q�wW"�բ�a�!�BL.��^R�!��x����7
l_I�)7ۓ ��{,�ux��Uk�1��t�x3*']G�P���S%"}gy06�
�
p���<����FO�.G��������>4���I�w���ci/�E����07�p<��[�I���=1� Z^n��Vs���+�,7L~<�k�9�<���E�"�d43�4���q���W�Q�^����޵;2�ٰ%ʱLv
d����DC���s LC���
5�p̷���k�y>�{�n.ݯ��k�<�y}3�|����g���t��R����҅������MVɂ>��2��EAuV��}�.Q�2��\}�@��b�$ ao�e�@b1�o�G�F�����2s�=�qMB@�⫹<%�}{����]�^�D����[�@� %�4B��C;XH��o�WK��vE�n�"���dŤo�G�؍�鏗��d�c�Z�jHٱ@��'���GgRWt�W���=��O���9D(i��ٰ�J��h��w25�){���KFdu����_���	���Z:u�e�3�����ܒj�lT�7)D٨FvZ�[�x3�W�c�Dh�R��x|��r}����;���^�RI�jZ��������~B���v���Y�����&��{7�c�T�����|����w~C�5yR��T��M�]�\O�+�S����������žTY���˙ ��6������$0\8�#�t�y~��㞠�3�f�NDw	�t<���Tc�:B3�2�on!�}���H-�9>�� �-4S���X9	9�I��0ޜmW��J''�ZS��,��|��q�!��� ���ޘuP&����I�5����Xs5O��~�nd*c����8e��S���w�ư�k~�n!`ܳk��v��<�#�4�v}"?[.sɏ*!x�<hi��`�H M�(ߘk")T)�o�/}����&ù�����zU���^��o�Y��#�F�F��O2��=`���*�_ʛ��]�<&'��;j��. jS��C�tz�����t�h�6�a��/k�t�,�U�Ӹ�D����$]\�N��m���oV�眒�ⰰ���AFi��JCkP�f�7 ߞ}q1�� �T�յ޼�`>���|o����`Ô��$[����8ظw��1��
ߣ�&�/k�_�Ҕ�C
��Ў�R[k)�[�	�Ր�I����X�И�6���<�}�w,#�;�q��z���T����vG�
�T"���D�����6��j��<�"���hP����k����^=���;XS�0�o3�Ϸgҭ}��NA�P�{��r��������?Ȁn���5���PV���x$YbO�����c����
��ޤW�̬ 2��u+'7�%�
�S~��/����71Q Ji��Q�g�}�?X9�
v�=x��v�I�Y1lz���ai#�3\�V椅"��i�Bخz�(�)+H���$[tm�u����.}��h��7xO:r��e�m���rNK���SJ�eED��-�YkDB'��0�����v��z^�o+))Vxd�	 }��u����*�݇6[]]E�;^@�Y����1�^&��D 4�1�UC�t�[�SԬ�~շ������&�rO8�Y��?���צ��ԡ��,|{�O���?4^U�����fQ��e=�X���,w��:�zpU�����#�_m���N(d��Q�*l�)��L>�w7*$$��P�uf�d,eä�5G��qq�) k����=`s\���x	>ܿ2\��]��h�s��|��F�t"_+3 y���*���c.�	�V���u$��&zYjǣy�=�г ��|^��ǝT"�{�-\�b[����H$ *�777��qڮD�W���'�u6���>�լ96e�6$_h����߿����Lk�dd�*c@��X�y�nݺ�8�MD^QQ�^��h,iﬦ��N���,�G��v��8�AB�RJ��Ʌc�Ō��<�T�}X]��u��jfHDkC6���hU[�+K7@�@��i��dd��6sݿ�^(---d!��dW�[�4[�Ϯ���'9c�ӓC@.���˫������{�,'���fA�k�N�a������Հ�)�n����{L���`'9s��ԏώ�;� ǯ�[�E3�s8o�ˤ�_��r�9�Rб���!�kT<x�d�_�-�	v?(��$B���c�,���`[Yx�i�s-�>��H��B�c��'�<g��,`pD����$5ł��'Ǉ˭��B'�;o��m��� /1����e�05u�6�U\~|�@���K�U�S��a>����s��"-բ�Vl�Řu;�m����6�y�j�ބS�ˡm*�t����rVf��Xvvv+��P� <C2tr�#�J�� 8S ��vNN�a�=}��ꨒx���bD1�G�b8-SFFF��	8'��m38���5�M\�u�73
G�å��SR��<161a�����Ύ����?��Ossr`�v4Am:�>  �u�L<i7|+��mo��.�]"�~e�J�;=';�Eĕ���4�"�Ѱ��.}��Ԥ*L�S���S߻��K�r!��!� �R�.���L����1�F!����צ�� K�Ml*12|�E8����\2�Z�n��U����R�����k��E!�������>@��� �gȍVGʅK���v�� ��B}�gJF0��T�I��8l5��/(��ʋM�N<�E��/�!d��㫝�YN)����C�����G�������#����|H�EP�n��O�t� �y�r���w���G������~�ip����)cO_�7a��p@�G�n��H�zhՖw�W�dt��1�m�}*�z-�л�oٮ�0��W��R�}뢼�-:c`�4HI�߹ ݏ�S�X�}� �X�~w �LIX||�l��.�3�-�[2�тg�d�ƕ���v���Y?6�B�da�!��tTk �e��^�[e����}`�*�����<K��kԩ����n����j*�8�zxu
�1����w���\�O3T>|@S�D/	���b��v{�J���_<Z��ݻ���SIu=F=����<o`L�����h�7<f�û�s}�����ܫ������d�M�/p��ڱ�����������A|D�T��:�(��KE%����c��p�l�zhR��{�
�n@o�@_�����-e�
��5;����H�8Ȓ�A|��%_����.�+4/���{�V�����5��&�;�Ik_�K�޺����A����~��eٴ��x4�t�k�b#Bm�������f��,�?g�l��꠶��,.�<�%�6��_t���o���$*+�/�"W@8���XG!Wт?Tf'i 5	+�p��,Л��Zz�� �#�,7e���'1�/	�K4���\���/�%^� J����4-~
�a��$�J]��K���)�/B�j���a�2Ia��J3]l���v|���E��n	���
�65gT��R�n���YA�X�&gk[�aU��v�lBXX��S��#�޻�8ᴎ����o^���g�DoU	D]&"C+���+�X�Q쪲|X:6���͘@t�V�4n֚��%ͅh�6�t�m���"͐��sa�tc��5�,��|~�Z$g���9�`���]j���5l�+̂��u�`�2�[�ט������8.�Yl��t�)��w�1��j^�b_�ÂJ.<L3�0���Q�������D�;H�V�(�=3�k���4���g�@�Ʈ}r�p���7��:`;eն$���B�S�!����n��!��a�X1r	#��v�4"�?�&s�4�j�꠆&������-�?���_6,gV(Wm�R+q�S')���+'r�L���� �*�[��%yYV��i�J�o��@�z.�w�9?�p��_UG��Wp�;P:�M!�)b�J#��~-�4;�-����*�/~:��k�e���*Jp3|%��sf������V��g!��	���F�QI'�-��F�ᕓ�j 
fP�?s)��aq�F��_Z�Ӎ�T����'<t��u�+jʖ?�ֺ�[]󕎐��<0��<�歾�X��i��\�f��3�xO�ioQfߞ��0���	9���#9�o��e�u�Kw��)6_��UسY��u��d[	�� ��j�H�ؽ��a�h�C��z�Mc��0��=��.N�gV��* �@��kT�3��=0.J)y{��'��F�r�6VUM-`��e�fi�������*1��4��G�1r�Hǲj0[����"t�T��۔�𹂎��r�Ɂ������p���_�X��y&g�0"����C��c?#9��]\�1.���>-x�59���l���ݒ�+�#Y���7g�v�f7�%D���|9��&�ͳ�=W��ښr;��X3f%:;[ҥz���ڗ ���H}�Rk�E��r�����98��Vm�+F����ҁ�(]��R�W��R�(���E�6azc[�&�=����@v{Ip-��!��!@N�h$�UW^��oJ�V�6�,g���y4&�����>�	#9C�"��b�D���=B���(��&�3�����ǝh������m�ćP0�[,�s�4N��|>Ȍ����HwY ��<ŕf*��r]�I�4�ˡ�x�a�~�	F����r>������"Ξ�ѵ�e�F�Zn��D�;0m-|���eg&�����A�kv�����1Wi/�������}�^�*K�Q�U��H�a��C�%5�Jok)��ֵ�;�=O�:8?�1��26�\n��3FRJD%�����B(�FW=�j[��B�� )ɨ`dd�w���\>XH� tٲ�݀O)�^4����(ۓ�^��8��<�=�<Ӹ,#W�s���A�8Z@�ى�� �Uת�v������3��'<��'�����TUc�N� pPH�"5]ă�~�����Z��0�x��F�����Vs9yeZ��#=9�y[dz�s�vHZ�7b@,�0�Zo�GF��U�o�Ef���>`ym+��[&��B'IVLd�Y��g���L�9��u<G� V(c�-��U"8'�E����I�/�����&������,_�=R�!S���@�ՅG����9	�䨖gת���eW����4ߖz���X�
%0�o¤�
�6&&�F�T۶�ɵ�?+��GL�a��e���O}� ��L��ϟ?�iy����������a���j��:S�rT�k_�ٿ�X?TMp�"&$�O޺��@Z�I�B��u÷W}�m;3J�� �Tb��qr�o�o���C%o�/�#�!�T�vt�,��	����[ 2BR��w�� w�!�S���=��-��x�MO!���*�A-��"��X�����g�r����KbqHa�ƚN��Af���*�Fdy�Ob�����͹�p ��W5B¢p11ج�%���zݽ�(����M���i�� ��EdL[���>�LB�9���Q21tɣ������?�)�����"+#�C���#[B���J���$+�d�B��Ce{��{��p���������Ox�_㺞����%L2{���Q+�/oe{������g��%:�I��>_�/�2-/.�J��D��}A�P�@��-�
DB�9/N�n.�&jpW��A�����z�B��5��@dٴ��.g&����YW���O���:�k2Mۣb�k�O�]&?C���|⽤�m>+$����s�F��"����S*-��>+�+qH�;pܠX��G�=a�`��H��}ҍ�"z�Ϗ�������|�d�����3ƚ��΂i\�����������	��w�*�����"�O}��ج|���Vg��5r������T��;�����ȉk�`�3]�~hbz�wu{g~=ñ��JN��N�Z�!����o����� ��������=�!�-�z��x71����aULX��,�ӗY��Z:�im�n'��Y ���"`�4;;�M���b�kHYYY^��#����,Gj2Ra�p{o��:���jl�(�/��Gq�'�}�l=R�a>��ʌ���)�8���o`� ��x>��3�juk?<��<#��8�a�50{����vk�bY4�@a���`P��~_�*;�[`W�]nCxs;��X�x�va_�c>ctz@�-����:[�w�0�2��00��H*ݲ���bJ&�&�*S�V�4 V~Na�o����\� C���\��/�����a�2�ĕ��� �*�7GQ�J�"�:��������E�1�ʅ�u��W�[t3欏dv���j�х��=Jh[����վ3���p
�E+x�<װ�@����&�,�>�����<�*�9`n��� ��-AA-A�s8�U�ik���%Fz��q�b���[;���J0�����7�p���������4`�tB ��Q�A���@���Y�O7�/߇6� י���=�I��f�ǼD<lſ<}�8��tU`Xϡ��3��UJJ�3�ev�qx}�y��~@�"�[C�WW���� ev�4=p�Xe�N�bh�~b��G�s:z�B�,S��b�9m�Tm�r-���z�%�x�=F;E@��O�zb��V�+����s ���ϣ�P`$���\LFJ?�H<��`�ң QXBs�Lz�E����}��!����q���ϝ�����,�l`�qz�q=���qH�Bp�;W͒��F���t^t�-?Yo��0��XD�^�N�,�f#C}[�L���ɭ0�o�V~��<�<��a�y�� vWvN�c�מ�C�Ik&ֈ���`�VIÜ?O ���l����{���D!��P�)�=��	�v�SC֚(�b���ᮉ�9�5����&��Mb[��������P�̂�Lz��AM�B&��/87!>�=�� 9�y�5;��|o]��7��5���"Y9_:T�8!���LA��� E�(� ���C0�����	�i�Q<�>qY|������V�����$�2��u�q�@$֦��	t�-g+�_%�h}A���̑�8n^����d��硸J�r,D���P��ù���fg��?th�����KM���Do؋�)�0��6Ő���5��y�B���~-r����:�Ϋ�N�6���T$���R)G��v���d���S5BW�q�1'�ө�����w+��,�wi�î����'�b�+��lzlF�$M.��K����e�����_g}���Fύ�B)��
!��Y�<�ߒ��
?؅o���A	�/���l�|�[�"��W*Q���
/d2��;1U��Yέ�]�=M�f����#�Qz&"��[��17$BZ�ʲ���r��BG6è{����t����"ց��xڄ����՟Յ�
��^�\���g3��-�i)��"��.N�!�g�9������vW�Ӕ"���_� l��������XJh�4��-s\�K��z����4M��Ϲ]����Jo��*�ś�
(2R�����<�%
#d����]����뼪)�oF���+���zR���OK�CI�����j\��~h�p"I�^��jio[���sM댋l�k<����e�=˸����鄪�:;�No�W���s��m�#ƃ��Yj3J�)�����dHl��z�u�Z�3h8�7 ����8��=L��
	��Z?��5�鱈/U�w~cK�R%%f��8u%w���:�.7�����UN�z�+�r����-6�Sn���0�R:{CJ���1�p���2�z�����I=R�H����Gr+�S��aO'w����ON�cS�΀�o���N�l�_��t��e�~��+�&ë��:�L��>Y�)��/�|�d}�M9�D>X���M\#F�i�hY齡,Ów��ev��]4��'oEۖA�{��cA�VV|�ǩ[��g{_GI���*v����Y��M�1W�[���Υ3�=���2�f"Vx՜��\���� C�1xsd$����������M�[2&Bme���P�ld� )�r���C��s�o~@�@j}�����q 1�Ǽ��0�_�r�(ի;�0��g��N+��$B���L��|j �T�˿Q�ѺҀ���S�{�lٟ��+���jc��"9��'�H���^�a8�M����ٹ9�Y1��߽�S3�̌��5Uݻ
*rCW�ߚK������?L���x?j"�!sG�c�uGw�2����w�e�V�b��|fJq$RǏ�˘�<b.��l�\�,/��_g��S��zU)�������Z�ܷgY�+�x��G@C���I;�$�3Y�Z��ڨ�a�5B���D�'Ӿ�癶ju<û�J�:h����`�*7�\�~ޱ��������PV[�w�'Y�w�v���J���;���g _�<�3�8zp����mKz��/��ٝf>�,~�ok�i�R�{dᖓ.6*�G�oEp���cޝ�)	Ģ���T���TB�L_΅�_־�u�(I����-�^�+qn�$�hVi���cd�7R�#��[���'=��ai�b�%�U��~����(�3��hͳ�ҔO��`)"�Σ(3О�S�WįH@��Cȝ��jdl[܌�������]�3�������M<�~�b��OT��w0�\�B6"v��T'�IOV�Mm~/u�a������m"=���Ԩ�Q���d�D�R@~�ku�:��?�xN(ׁ�,��ғ|v�m~�F�5`O*��uKƤ ��l(x�P�V]W7Cg�˃�ub.] ���"w�y�Z���fTAEҮ�ˁڪh(��h*���e��S[M��T��l�i�u�\T���5-.K�-�:36������8	�t���w@�� �}JW��9��SV�r&�a��ye���n�WIz���v��S|�N3 c
G/<uSz��B�ҁ(�|��IA��ʚM��a���z7M��#;-���V�r�[�D�����A{Oׅ�,��j��h��Vn�t*q�ׁ��cn�KٺA(Z_�`;/�~^�����������W�b�~��ZjwO��W�+�bq�B��L����&V�Va�Ǔ�We�J���3~8�Q?��x	ߵ�����7>(qj[���d�,v_~9}�τ]~�D�0�v�ѕP�n�l����/�G�ϖ^�r�aC�#�:��ٞ�E��?bDu��l8:���$�f��-!�s�,�����aBtt;8;;�y�(�n���$9����������k��u���!wk��4w�$ux�R�0��C��4K��%��c�%���Ș,���/D�|����dO�#��y��+H2�W,�e��B�W�36����Q��F ���[����b̮�sC ���мN���e"r��Q���WT��ԙ�z3�����L?��ˬ��_���1-�Ztʺ1�f�5�����GL���#���<6���C<N�]j�P��)�G3ї��2�� ˬd&����zL��NOtm����;�;�X�}�g���j�E�ZTO��ﲔsB��ܔ����?�B�8��#�h:Pq����b	햳��ۜ-���m�huo�v�ie�wX(*y�e&`G��w��&Rr,�0R��`�����L��:��v��s�@��k 8�:88(?;I����f���u�����  9�n�&�1�d�����^v��D6��M}�%�&;G��)[��2�z��z-S*�	n^u�RȎ��"��@22���	� ���)'���Lh� 11��45� �j�,�93?ϟx��o-`�1`�~}L�FJF���DL��Y�%=�ff[���-���F����N����r�6�yxW<,�z�J�:��T:|�V�M wblX���\K ��T|��p�4J]	`���7����݆�����DFD ���ӯ����W�H�ae �ee^ �\h�km�1�ѕ��/n����K�9x�o��x�%��
�񥮭c�9����Aw�Z�$�N��l~�TQ��Ȕ��@oW�|��/<��a�H÷��%ϊ1U�mjRq�z-THc�{#,f��JJJ<�
Znz���HU8e2<]�C/��͈`��K=O�OzN��R��.����U$0dc=��lN�:��={&?5b?�bt�v���W� �Q;�7�����?�q�_�b�6��@�o��z��Ib�e��U����(��]����
�u�������*�Z:��"q� � �9���TO�8��Y��Xʷ3%N?o�GJ��Dw�n!
P�څ�7@]t��T�(K��ΰ��(yæ^F����?t���}��5{�
=[���\2P,;�v�r���z����N�Y9����ɓ�!�y�ZCKk6�ed�~�1g �e[�m�elY%,������[�;���.4�6:�p��!���w M���=���;4��"o
�s���-'uT��?&q��9(�Z�?�䕏9cR��g�Ie��֚����AZ�{��c�1|�kYl�Y��8|*���D��ї{���y������9�Od�nӼ���dX�����5i`c��&8,�`lS!+�-���b28̼"-�w	�H��o�.j+��`�*('X��L��u�������3���0�@Rf)=�M�����^rQ�9t�[B��X��!r���ϽC�7�31{� ����{�n'�\b���L�y�.�����T�*�f-֟}��'��];b�ya�#�=���yQȚo��y����**)$�O�]�*�펏��%��m�J��ws1�	aY���fE�����h��q�����X��L��.�s
�x�h�(�W��,����~��aǅ�\`����V�9���S� �w!�*霿��p,��JV��O`/���.��O�o�C*�y��w$ͨ�\|5��&��~h�)�Ce�[�c@,�q떲��ّ �t&{{�xl�g��8��͊^� 9��f�x9�y^��4g;�%�% ��S2} OEYݩ�Y�L�g�]Y{��7g�sF;��[Zx1����ފ���gB�gvf�a��V1�����Mp�+6�AU5�/���"�3�fm��(!;��&^�,��Z���f�K�����������A���6�5� jd�z�T��K�d��B��)��!x;��j��.�ٱ��8+��bCy�'�P����ٝ�S�U���aΪ�K�	-��q)KD'/�� �D�� 
��\�g��G����Ml\�)׼���������� .B-@y�A��?�V�.V7F"U�)��F�0F�ʘ��ˈ�Tl'���V���D�,W�T��
�ǀz�H��)�I=�I���.>�'ru.�:�˪��W����r�y#����d���w�B��X���	>?6 ����U���Gd��і���)6�`	+�T�[Ұm���,�n���墓����h�u���Di��}�������E�h���T}����آ=�<i5 �����r�"n 	QF<OD�Xe� q�t���ۡ�^�̀��>��q�����ωS5��ru@Lk
2br_
��q��	hO���0b�I	ߢ�z��U��##�L"��Y�Z�y�ށx���o�{#O��j�1'��p�b4PVY��C g����Eh����wS�R R{8�Y�)����s.�w`S�~��r�l\�I(�uQ�����=��*���S~ĉ�d��]9�},ਗ��|j�?��2oe�y��W2jkG��׿��jI쟋4j��Ѷ�l�f��<�rL�}�c'A��k�*=i���Zg����1�c��Et�B�xGcm�����_�z>�����X��P���;0`!B�؄�VꚚ�p`�}���E��*���*�uB2���Gm<H&��a瘝de{#8*T ���">��zWbs��`�z�JWR���E%Kp�'�{FQ���3�r9���_���)\8 �tr�,�?m�8X�D����-c�Ȝ �F��Rd�4�y3�3J�	��@`ݕoed�1���*�dK~6}�5�Im�>��3�%�����s�F�5q�wh�}����g�<�*++��6m�4�I��ϐaUL��K/����u�iSm�^�NK��Uj���Y�~���pҀ�v�1B�Uu%�v�r}�cH�Q��@�K ����/Nk!ߌ<�nQ�KJ1Y��@g�982a�'B�Tn1&>3~�E�{���V"�jڍ!Z���IO6w���)8$w�)��9e���T�:��	Ł  �wfx��'m��H�x�;ʴ���b�t����)3�[L��b/��,,�<R�����f��`%:��`wB++E�����e����«��x�퉒ף'F�דn��_r��7,;W��R��I���9�p�RK�UU��I*}�+,���3�t�f���J\�o�����}��p�
�a�,��yW�����w�=q�Ny��+�������v^w1�!}b"q�����%Zú.�5�����NCA%6��U�/v��E�����'4����;(ȕb�?�Qc��/_L���V�`D��n�r0�� �����m��,ws,����`��R���ի�����e�U�����y���̠�i�����>���V�r��/:��aVB� r:_(8����8�y`@�BZ֛(��/�m����xxT�o��pLzo�g�����̨F7f�NFX���7�����g��-ʰ9����h�v3?��z���|�`���	ۄ��(�ͬo)�}~��ou�d�	*n���_=�<��1��y3��W�c����@�4J���k�?�㯜�Α���>��6P`Qd9hp��*�A�w&�ܠHb'����RZE��S��j�O�*�����pv��sX�y�8o��Eg5Y,\"��'T\�0_��а�u�$��]3�%�+�g��9@Q�g���A'1��*�X�Y��4[�>��#ȕ(ޚNb��}譌�[�'2Zk�DzzN��Y��MH��?�8���e����M� ��½��It�-@�h�.\����?�k�N�|��QF�_�,����C� �����fx9s�-U*��h�3 �L��3�,ޱ:�cu9\�D~��	����]�z�b�_܈{�ϴU=R	�-�,�Ɛ�W�
�-���UZ�EɛJ�n���SH���P�{ҩ]]\v�'� ���Gu���? k|�e�}.��ا"!dC�(d���|�V?��`L��4=�S�L��z!�b�<�F���0g��'�a���Z>К�\�i{]/�S@�%�@��D�l�v�ۮ��k2\���ˏ9�IД�\���e�N,�����E�!����wXXi��z�0��NS���w[˩H5�\��P����ɒ�4��Fj���(�)`	�хo���7+^)�j�q!�l��#u���T1	�1�{vL������BH�Ӊe���r^�l�%zw�c�)ʈ8����3Կb�5���`g�����c1�Ghr7(8C^���DCQ���h�&RK�o��\.�M�F*��P����q�� �":ь�:{yE�k�R;w��T�BN���|��o�K����w��*�M9=I��P랤�q�e����8Յ���� �'VT�V��|���m���C�$(5WH��:�+6���5����:����7Cq�p�;%5]��eu������a��v^�k��(k�K���0�.:�%.��{�^^��<�?�;�(��z�2�)E�3ݙ�c�o4�bt�'zlL׆G��ʤd��n�h��}��Z�QOgvuY7]�;0��
I,{�l��w�s�0ǻ��6!FmB`p�����*����v� 2�g�p�τ��v>���^4�K~\6��Mf�����3�Cy88h*BR"ZvjPM��&f�������Z��O|�S��P-c��P�>p���r%k���A���	���Aɇ{S+�5��U��`?�l���WR+;���u�w���C��X3{=��5��p�]�����T����[59��W�Adt4Th˗��S�6�����⽿u6q�r��(��ɒx��zF�>C��͇>�~|��Gva��P���pq�]X��QK�%<oؾ�5�d�&��YG�O�ݐ�줺Ȉ�3!D�;����YU��쪻�qI��r��-_rz���n��H[5�\O
=ձ���R,*Q�cM)��-x�5R3A%��r6V7u�hފ�b�b���� ,Tc%O�3�0���=�x���oԅ�y��@�ؓ�fv���^����V��SI�OzP���aH���k�Ū#�&׻�U7��!�w�2�� Z�MI��T�h힎$����NX�+)�9|5�U�[U':6Pk�Խ�Yu�7�;t%��O�kbx> �)��#�����;���{kY���⁉�o��D�A��,V�*��2�ku��%��]�h��mˬ�)�rC3�鼿K�v��)�>�|��׮�����>K���Lo�<{ȪQ�C���2#4�9�ڣV'�A�����ah���ǀ���^ס޻p�B\��bML���1o��-���a�;�;��֗�Dֺ��N�Rw~-"ߒP��<v����h���8�R�r���E�;�N��>��iZ��T��wN?��w���c.���ٌ2+T�ߓ.���X��:�.���J>�9+q��B�p����"0�F�d2�;s�9S�>��.�h7�?�H�$ͮ�p����g.A�x-�Y$���`u��f�F,��XJBM8;��M�s���ֻcM�)�HY����������.T���{vʻ^^U���1g��"j*h�[��h!��U]���;�����������#�����+_cc�*E=`*��c���'ۥQ�T+v�#ʱ�(�E[���<�����S$�>Ć�ͻ��%��}�j�~��%���Ӛ<؜Z@�X�D�n���1���]��\��,�Xhcq�� ���h)��ai##P���no�S-t��qƭ��rx�*��Jm��=�El̆'��J K�7�^��������l�LD���%�Fh�s����lBǻ�6<���������oB�՜��ϕ�]p��u��Iiw���X���=���+�@� q(8�t��̏����U��ij�yR�����\v"������B�+��٩]�
bO~�]-5�W��K��ڬ;��;u�sr6VVH+D� ���~*�����wH�K;Eٲѝ�9�(}^��g	q�:؄RNzc�6� aN���P��@}��>At��!|��.Z��o�}}���B��S��)�>1�2���	]<�tL���V�n�F�������Sח��(7	1�Q]��<�)T����o!��͢�ػ� �U�k_ϸ��9���1so
�CbB$%-x&sb{*5Wgwi�}�������J���!g��y���ꮞ���֝���<F�|?�ɥ1]��Mu�`C�pxv&�E�]rz��tVfRO ��qgWW���`�]r�HubG� �[t����SI��5^����7��u�e]0߸����X����	������BH�d�A�&�'k:v����6��B�-,��P{�32�.\�03;�fe�s��7��Or��H��ܢΞ�,5~����f��H�.��m|f,3P!$>�el��-����Sd�WN�(^@	������$1/ys��������[l�S
�b�f�}��2Y]B�%R���^Cؤ��:f���LJ
B5�u�t�A��C��Dq8j��N��b3�PR�w(�>��u���ԯ�Q��=KD�����<ۄb���obUu��j�.����´ֵh��kGO���',-��z/xGo�F�q�������b�z�f���L��WF҈>����DHrÌ>�n
�\�"Q7����1��>�7la�����d.�a��^��tIH��x�G��V�����eG�?��e����3S2����Md/	nt�E>��|n���?�4w	3�6��F}ԟ�Z�-G*��R�N�����CX�3u�i�`��d��|2Г53ە����JҍL��QUU�B�����KO�n�X\�v83U����ח��6��;�iiD�B:9��	��U<��p����	oJ`;�u�jQ���[���~�mиw�=��Y��)HgR���ֹ0�j�K
N!d�FM�	��_�K�^ M�D�Hf"舢.u�4X�&{.�ѯ�79�i��掿���rc�K<�Pp�:�|�� �ŝ�@{ߏ��5Y�M�kw�AkJy��<���^�����p����|��[Ӧȵ�[� ��v�?��B���4�h*�j�?�,��9������P���e�%T�{}�����GKf����!�Tm[ՙ��m��r`�U�(���4O�J�Q�ۙ�[�C��P�����b���}w��+��<y8����w�⺫9$Jn�篣(���S|����;9_��s�y
U����:���6 =~��^�޾v�S�=M|	�h��*n)�Z��5v9^�ﺙ�K�C\1�>4mţ� G�o����{�X��S�D���m�7t��U:����Qe�L&�/�*��.��>w.} <آ/��v��W�O|�'1<����G��� �����Ҁ�`����&�;�)����ڋ��������h�R=h����Js��JO ���E��e��3F��?��v3��U�����pC��[�*_��D�O�wۉKh�E���"i�_,YCE-��^az�T�h���Q��eT�"��6^@��sor�c��@��'�1��쏇�W.�(��/j�x�$?��}�V��9X�2&����jv�o1ﺑH$�G�S���^Ȣ:Q])��/�a�|�⑈� _��� E���*�i��<���M�+v$N�{u�<Bt��48I����n�@;@�I  �E9:E+���,�(_,���5�����HO�����ϓ%^bQ�KK��
���CT���C�{u���m/!�^�R�h Eh��\_�?Y�����s�<G~\��2���-�]��z���)@�Aiii��_C����ō������o��>6�<����8�D7��V"d�.��kc�3(���U������z∫h��[��P��P aL�y�� U�o�tU��˖;Lј{��+,�6�p��6�����������򙁯/ٖ߁����8��^u��?�^���[Z��"���m�{�x�$���p�H��b)��Q��A7`OP��e��d���Q�v��o ���[&��A���+�gQ��y�D�G���
|�(�o�K�NļI]C�bgj�4��ֶv%��:p��x����a���ۭ�v���q�:���'��${,4B�.��?T�ڟ���;���ݟ��[|usf�Rl��";?� �p�^h���V���i�`/Y��호��|�S9�(6��ϝ���*��
ȱ)��`���7�y��������l��b��^��ӯ�g�V
��C�yh[T���\Q{|G�]�<����<���.3Yp�$"�G16t6������Qr"��є[-ŏ�'	�i�q�@M�~��-K_v_��E&<]��6���<�@tdDD��fDDtgfn���صޝ򿔚�@�fs��qs{��[j	\,��ߑ�7+�S8{�>|]�9D���
Sg�X$�e�^
C���=��s2���
���N�bI��:�O����W�� � W��7��{Ac��I]vx��4*���'���Ipk�e?e�\P����JL�E��ܟ��65�B��96 @hv�ڵ�ƹ텤�UwY��� H�̬Z��m��'Ђjl��ӫW�b;ө�C��ml;nu9!>{c3��<�N:�rrP��Y�E�.�'w�Z���A� ���H{>�:���ּ�Yڎ��\��T6(�/֓y\:� ��,ߩ�E/��'��nw�?�vtqq����OV���Sc�����j�3��+}��(�A��"��H�R���Ƃ��0�z�X�+ �wp�0=�_���`� ��E�2����}�o�|�!嚹��BE�P˄y;]��N�>��.	R}�zݾjo]2K�����@�0b����"�6[�!��o)�*e�e��Z��mI�aߋ���n��aw=v))����!E@]�s4�z��}1	��ceS�8�K�R콿sL;{�ꍚ��Z;�S��M���۝U>��(N�մ��0D�%|���ahz������Fɇ�\&##өr͓��`~I.�z7tR��{�m�TK��tL��s�/�[PP�b*	Y�9"jv��xP��]��T��L`�T�r�y��9B�*�<R���g��@w^�bB{��SX�|��U%"��:�a��ں��q�5�O(� ��t+��]�wsg�(�7����E�b��'^�1 ���`��0+�+Deq̰`vd�D,?s$%v1`�C]�P3��`���躛+;�
Z��m�]�� ��.]5�X$v3x
�f\)H_�yU�,ɋ��o������2��f���hp,eT�xVb�^>ߡ�����D�7;T���G��s�.�"L�����_�I^"��@w�@���R(���O�c��hm}Ü��2�X������^dԏ�(�Ϊ����D�R��G�n~����YH]���Wd�c�F�!=&���r٨�n���L��$�E:�!_6�'��qOp��ODT���p��u����KLO:_g�"4>}}}���_i��9�`V��? � m��.~�F�P��v���h�?�����!f6ڠ��P=s6�u�eg�H�K���}8`]j�%i����aI�.<��$Յ��Er�&l� ���e���W咥jl��F[5\A�4m6�X\Ϧ��=���S�I����l���<ݲ�*�]����S��dg�P�U@o��F���x�NbF�G;݇�dӝ�l�0�Zlʸ0�XK��T�G����JIF�� �}���n�@����0�0�hɒ�eJ$af�����E�"���;��R��b��a[���,���[F�U ��Ӓ��[N�D�g���w$�&�w����~z��m��0]\��Cx�^���!`��Ȫ�R�Q��P��xC?�I{,�(������%�F�4���"P���Y�(J��������] d�\���mFkk���g�s����e�`<�#C��u���|a�$j`��I�;mU��	���%?��i�qý�B2�������>���{>�j�+;�v6'ͬ�̬¯aj��K�{�C�����G�z��9c�sz��tR$�Ɣ����ܦzVZL��,Ӧ�Z�g���&ɠ��'������N����Nv�#S�.�ZP�����2�������j��Uk�N�P�D�L�BX߱���ή�}�9Z�C|��p�o��T��m���h�2v:#�b�zM:�
��*�kS_nn��ϕ����|��I�?z�^��iw~s܍��]��zz�6F$�^�W���������;�%y��*��U�Jm�V�Ӈ���M�W-���(��/����<?�ǳ�O?��Gw�QM�M�e�OP�F�s�q��%Jҗ���]\0r�;aؓNf|�!�AAA�ۓ�%ƍ���ŝ.Uh(��1`6�@���ٲ�}:�6�1�%����n�F�7���Jɪ<�bM� �������^;͂��m٣�v�`+�I�4��/�}O�6���n��i����%�̴�{[g���j�����w�M�Ug7m����
���Y���7�ܺ7���+�7��7�ݒ��I
�~k���Io9����\����X�)"5`��0���]�]C�7�N�ul�肐ڔ�'&���
	I3a������R ���Ɏx�*��9�W�И����'��/&m�P����:iMp]�����4j�Qt_�Z��9�
��3Ԅ�a��S\&I�o�Sۡ˹А8�Y)y�zh���<��f3�ÇϽ(C�(��e�1a+�o[5/�����1�	JPpa�0�����D�<�9��D�R���1�]�q��A�V���s��,�\�$S�<=noTt-��/��[��3��B��d���s[5�"#�o����)L׽�2D�ա#�|�S
�-�R��#k�(�!�N����gTxyUq��9���;�oO{ҭ��$A���d��0��}vYM#�+�ڽ�{muw��ʭ޾~�켼;6��sH$���y_A����ଜ��w56C�.}j��Z�5ka �.	X�,�a�.P��6��Y;:_���ŭ��-+�J�g���J�ī�f��ҁ�Aے�B�3�vRCKW�
��-���4␰��3tʮє�dJP^}�>n��`����_1}�+��
e�(�M۩l~|����u�5j7�p�,tL�%�9,�	���⽖Z9�_�$%5����ɹg�n�*�g� /���w�JcK������<�����CZ��[��b�>N M��x�nܹ8+���/v��ʫ���F,�^�� ��cϜ��*�A['S��֚v��|�� T���?��9Tf��\ǹ�~F==}���*�.�8@L�ڙ��2�]��˚3%b}տj9Y�_���%��y�hO�4AG��=4��ϭ�,�?������~�5�`��q�F������c�`�}�:��s�{"�k����xl�^z��2��!z��zP�f����Ay�>alY�<ٕ�]7B�r������CϵCP�~Q��Ss"�;& z����O��\K��M�\-nF�v�6��J]έi�A!u�����F�UyYB�1�Y��.�����P8:�`�G�}`�	�f/��_i[t��s�ٴ[>Y���	�� ��uɒ�����rPx�R1dh�h���婏��ξ�4���}%�6�Y��{���gfg�W��~��6M����#/��\l�U
�T��n?�w�ۓ��o����&���t��p3��k�/h�y M���������%�c3g��`jǠ��u��C����-����Bwj8>1��v1Z�^zpX1^1�.�'CPfq&_��=��3�5~��~��b�WJ&��<ֿۓ��Z�4�����n��GA���Ÿc/��\�ը)�N��~�l�3����-J�M#����Sn*���6�o/N�`��2Uy��P�bb(J�zSQ�2&;[N_�{i�}���i�Q�kw��>��==3�O�2U&��>�>��' ���%�[�j;3Zu����wԩ�˯7-�:�a>���%��2�z4؆s���������?s(������H��A����ý26vg-L�_�����������q�5�0,h3�����iY����?�gZ�%_�.����R�[a�&]�@��3�>s�ʤ���ͤ��*�?|#���ڼ�#7�]N:�Xk��11��$}��t+��TZ��g&o�{�e:r]�;a��]���� )�"�v�?��^O�{�x䢯�Wr-ᘤ�S^�M:�l�ӊ{��<?�0xb��f�ǥ}�L��K{�+"��ν�y�m P[��6�h�A}԰�&��0�/y>84�ު�z�j�#����-6�+Wh%[�.��?+�j�z�.^h[��6�'ok���z��-�*��%?C�<���XS�\]_�S����ש�;D��<޸���<���C@Ƈ^ر����>�*�.&[W�{�E�oy��W�vT�_9󸿓hFӈ{+ii�y(�r<$L|�r�(-�������0Z��9>�6���ћ�#��]ö�]"֤�ڂB��}��Mڣ�K[�
�^{��9Co8�2�:k>���r���=��wf��ݫ9�5��}����*�����OB813��b����dʋ�2hƓp�����װ����@���$���@ww��{LD�x�1#��]J"vix37)����s���P�N��03��;&D{>��r��If���`���,��6��󔠹cW�Swݪ�%�����/#��cC�{l#s'�?{ !-.��'��y��g����v��]:vt�*r��d���S�����仉h6�J�Hb��$:et>����ȘH~��x@������u���RbJ:z�kaD�EJ;�n��LU6�}#�[�eͅV߻��#)���MT��%����k�C�q�0[�l�lrgr�X)Rd�����OfnL�C�Ю����'�V�X���Hf~�+5����ݿR�6��plog_����vxp�؉㚩�_f���#UA'�8�+Q+��L�+8����ֻ�͕�|��t��s��j7ۆ�eWKkY�^�Go�%�U�,�Ƨ��E�_QN՜$H:1��_/���'CB�'�8!���b��]����Ȩ�'�/�Gk�$��w_Oo|\�V{�m������Ì�?�f!��U�f�U��R���p0��KZ*��üu��%'n��u@���9UB�2��c�-��A�Ж�]u5�C٣[k+�Q��%��*:S�3^�v��I3ݩ~�?mV*�*��_v��/_���2�^su�������+g�/�
q�b���J��|�j���:l��X��4t�WmJM�K�Q`www.�p2>��0���u���jd�Aى�����Z�ɦz��M��`(��n8T�^����p�XDf�:Y5¹�0�TP$�D�y�{���ܪ�1p�-��,}_�>���L��_���	�
6&���������@T�1ol	
�P(��U��EW�n*;���l��8������5�t�6w4�:T���!���ަ�%~p��Ю�Ҏ�-i\V�e�3�������\O���'�ő�D�Njj��X�� ����\�_=�5aD����#�b�<]t-��?Qi[O@#߭�2.�缮�
�.o���<��SN7a�X���dI��D������B�(X����fՒw"����ɠj�<��;�����ӳ�]���4fz���C��Y��������t9;����W�Ӟ��=�S�h]t�Xo����m���'yJo�v�]�S^x������\j�zp[|Ջ^G�����nv�ޗ�� yN*]�T��<���C���򊉄�}��	���YN`[�}ZU�6�B���QWos7�y�xd�(z�y!��=�o���
n4.�*�I�{�2�g	��}L2�a��jJe�p���y�~2�q���.��q`H���ԝ�C���'�v�f��<i��N��ޮb$����k��w��(k̯�I���#;�C��o��yL%B���oN,)�k�d��k͊�����agƤt�C�}AI���Y0g���������l�Χng����A�T���a��o�M��XS�^���+'1¬��L����y,��}�a�i`����ca͎[�=�t��s6�4�`�6\��R	�6��`��E� �W��^}������z�ݜ��Gl2J��=�J�ʯ��|��)�W��}^�?H�X����M ������r�qs@o�ۍ�Gg�!m�Q6e"�xcU��z�\O׾�u�)뗽���u����f��8*IL*���ۆ,��kDV�}9=7<=ʸ���>��Fte0�`���Ƹ�6=�ホY@��G��'?��ﭼ-�eV���r�a��P6�v�d�;?�?3֔A#�\�gJS����y-0�]�+�C���?y���yI������|Ծ���;a�s�����i��ժW_Reb��s&�{��M�|T����k�vP8�9��]�xR�4N��x���R�'�0��6sa�� �I$3Y��fC��8��4@O�SO����~siD�ˏe��{����/"VYQ�[J�|���:Rk-6~�G+!�I�s���#4�H�R�K4����$���_���|�I�-ł�e@@�t�s5�/x�mQ�y&����#�!+�U��iaw[�N$�Q2w�\�ZV��p�1 �ڦ/?j�p��'X"��N���[����>����{�*��}�xDiRB��PA�D�tw7"-� ��{�Hwwl�κA|y�q�:g�1���ϡc��{͹f\�k��֣DE��f�3�eRp��l��nM�OAzx��P_ʓ�+������|���� �E�f�ա{�&5���Q�5p�dP)���ݽ��R���,�*ׁj(�@�}��c�sq.�zx�>f8��8[�ᢾځ��oV�fR=^�C���4�7��B��?�m��V�7Sor -,�*H��	��{���P+*�Q��Z8�_�E�����>+*���H�	�ߦxJ��O�]Y��7� &���{�D2��N��&��;��ٳ�/�"FC����>Ɵ�N�'�$N]u�xZ~�q[ߖ���(mS�ӕ���F��Lh��٠Uwö~����ڒ���V.���?���̹؟�r�� �N��W(����4w�����A�TE#�}�|����qO���n�k(�濂r����$g�K%�����P�[)n�t��8;��!q�3�&�A�j^3������*��˾�݊-bV�I���d��r�(G�q�X��З*m!��J�P���{vP��-�P]��j�d��dH����I#z�P<��[;��J�ޥ�u��j|�y�+\q�Ml�_o�?>�P-��*�ai�8�����="9?@��$�mI���R4!�b�4���VۇV]��{�O/���:f����)����T�d�8��[����*M��O(7���2m��mt9�h�R�D�� 9q
 |>�xd�C<6!Qv#΃J�|�i#Մ}'��k@ۼ������ǰa�|'�*J��L7F��|k���;Ʌ;^4=�蠖��������I�&�����&'Z��ҥ�|)$�z��U~ h�=ܮ\�8�r~s���5ߖ����W�x+]oA��,��.ETs%(��O�9���H�)�
�-�۹%��1%�rBZch_�{͕8�Yˡ���-��3� ��s���� �mo��._�Ů �� ��݅�R�G�����ғR�(D��(z���>���%Q��X&F�8��#�|�� I�����G�}����U���][��R�i7Y4��?�T�%n�s�z`%��_%I����p��6
jm�/�����
�ՙ�mDH*�2�y{R��QP�`��=��(�9+�1��^d��u\s���/p�׫�0�*n�6������C��g�+���й���@d�a��@���:-�>q�~1>O�n�vm�ɚ`��@�:��Tv��7:Q>��&B�~�����S&Ꮋ�1������OC�xr.diՊ�O ҕ�� l���!.��+�|�8xԸ�zl��3���ťϧ"L 'T����̡21c�� �=��0o����[wvϖ`RW:��� �G���4�Eq������K��˨>�)5�����F�n�ҽR53燖����]^���M�w�#����zH�-O>A��m� z<N�T��4�L|�T�]T�)]R��MC����q^^��~8(+�ֹ����u�D�k.�����l�'��>"��@N�o��"�d�-ǖqlW�2�A���n���h�^�!Ʌ݅X%���{1�R������FO�wv_
��5l���o7�]qZ�	�4�s��`o�TI��U��w�|5�*w^>61����>���	���C��^�9��Jw+����d�t�u�"8ˠ\�`��@Vf�Չ��^�"ǽ��w�`�#FFϝt2���K��|���l�r[�Z8��;��ڮ���s���4�0�١��W� daD�W[jU M������:����NB��Zg����k/������'Gpb]����z1�� �����u���=@k<m��kC�d�A#Yv�κ��O��Vsa^�ɒ�����_E�� �㪖�)
�E�\��R��a/`Im�̛T�e-�X�KUrj�G$жg��M<�4�#���Egz�J�KOLL<���*��d����xĭ�80�u��T	��e=�Y�ό�/�"Lr>��%ut����y���yl�w]�ߔ]�K�Qq"�1ҝx��E�={�{Л$��^e��^'ͦ�T��Y#�/���FW�cG�+��]�zI��2�,�@݀D��Kw�w�w�L��<�ЏWo�&��SY�9�d���R�D��Ǡ��q�:�7�������������B:���`���6��Q�`I_٧�7�ˑ9,#Kj=l,[Lj���E�wP.�g�����`�M�N�!��l�xضg2����@�"�g��A�:�"(%M�M+W(���cM�(x�⹇��ꤔ�ƥd<��e��r{ƺ~������s�
j�nv��	ٽ���sƺEF0w���,�W���*l�ل�/h.�����ʎ6[��gC����@ߑ��6�j�U!�`�����ׁw�
y�g�~���'�B���GOL�1<?!�_BVeu�=4��7���ZDA�yD��Ź^����gӮ �޼�js��s��d�ˑ���:w���|ҭ�r���`v�I9�]8���r�FV��������QL�>�P�G�h��,�c�u��{(6K�{/}���O����>]uZV��^,�UQ�}�����5t�1*�(��5q3_V��D.��;��Y6�4�Ԙ�ta?��Xf�:d�W���>�4�|�~C�Fg�3�4��ڼ=S�Ł�4Vץ�Q��:.���z*����!��~���.����}P��t5k��$�
]��3���8_I*�.��"��ѿl�K/F�>ܾ-��9����JwI������oee���DZo~���92�pKū0��ن�v${qc��[>'��nC�@���ݱ��l{�a�k܄�<d�W�r�=�wz�G��8�x9	#�����G�^+)E�2����dE�zd��[	�
4'���W��+�(2�^��>��t���M	�T��n�4:�Դ�ļ�#��O���	w6N�չ��_i��ƋNSo�#z��e:^�g��-ah�_G�=�-wZ�\r���:��S�]!ϊb</r+��Iѱ)��K��h�/�姊w��_��"aru+��Bկ���9�\�ey>3����%��re�.A�蕷-Ж����U��u����0�K��B����W=l/&��yv�u��N��}&�p�٠aw�kB��h:B
�%��Hz�og0�mm+*�>�:jE[��L�&F��Q3<X@��M�Sg�U�n��t�p%:��r��i=ZV��?�=�C���E{�Ɖ:��xQލ[T����5� -�u�'��4��!T
��\�����M8�w��?�1y6���Xn�_0#ͳ�k?P���]��|��DD1���t|�5w���"��_n}r^�G����F���B=��Z�t�4�d�g<�t1�זw`)J��N���MT�ろ����$�Z�u('��A+*���3�~J�:��G��{����*F���0��'>�{�������F��l�ѥ����֫]>D\ }�D���2�F0R��`��E$��̱���ɸ\[b7m����8��.�r�m���\Nt�o�we���P�ؽ1��;��1/糩��r�bw=��ֆ_R�/�o/�*�Ď_��f���=##Y���#�Uf8�5t�:�F�U��]F���˩K4�u�6��Ҁ�j����ȿm5��RC��e)��t�+���	2�!�R��"��s���B��$n#���b:��?�]�}dr~�	�k�p�Z��")�&= �}��cATis�\�6N�p�M�#�Q��-1��1��T��c��D�S9 �~��Z���[n����-�D�t�.�rT�\.��8W�3�?�x���GZOP���=�hn�3�kW&N�Wx�mf��|��̰L��s��,,�V^/�=��%'t��K��`��!C;k��1��T�ݳx�bޮĐ������g���������I����N����Җ��B-���-٬5a7��?WϿ������[$�H��y+=��>4UL*3�[�V��Ͼ����f\+���WX��</(�Xb���	>45R.�-'-/��7�&x�Ԡ�x_��#*/e`�1�\o`���]ά�_K��uqxQZe�&�������S$�f:�֊v{/���#��ʗ�A>�)�"���jŋ��k�s!�B?oYa40z�J�3K���bQ
G �Z�db�c����D�7�Z�}K�X!�	����WAi�f����~����1u�A��t�lJwJ���[�^��z!�z2��F��;q��J}ͦ�-�JV&�����_l�|̀�^��x�P�:�/i�U��Z!�j2��O7?�*$	�-��d��/�抓8�:ԋ	-*������æ���B{=<�Z��rWM�}Y��q�[
& ca�����u��~�c\+Lf�8vb��~_�f����nW�{� xG4%�ٜT`e��/�����,(�7�����@�z8�����yt�r~봹C���o5c
�͝TvmiNM�?�@4����-}{�U+�~7n��%+W�`F���i
G�\h� ���_��B����䟥���=���F}Ez�H﮾���]��d�j�d:���1Y�I���h����ʬ��+���/�\�l5��؝�k�o��knk�Y�O��&���C����{mk����x���r�hn��vQ��Q��������Ğ�A͆����!J�:��%=%�_ȌjZ�%Z�>��hQ��u�����Z�x��:P�����T������J���6���I4�Y�ae��7��7���"�����ԭ�5�:
4y��hWf*���z/�����s.P�˅u�$�DK}����%2Z%�aB���8H�\���M��EɽP�e�4�Ӝ.����[�;�\������]��6$g���X�)�U�S����?J}�9���[����G��֜�h���9]+�ټf�f+��=R��~����[��.J��t�(�΂�]����vL3֛x7K�td��ʨV�Hs����ʧ-��\�<1�v�߲�|�ꂯx�g���*�|�IG��J�;^� ��uP#�K�]�쮔6�;W�F�u�uIE/tz���~�hjhm�u;,�xI*�n���L�|Ht3MC��'ԝ�bb]���)Y'��ģ��Y?��;t�R�I���]�^�
�{�G+ŧum�޿`k2���U��6�_Oߙ�K�I�c���2v��EaJ,���|�8�6�|�+]��+�<zQ�����'"	4/�M�C3+S�O�+�d>Wv��@'q)F��p�l�$jQ|��%��x���;�n�Y��VϨT[��KO�>�+�\1�5co�����>�Z�A;-D]���\�9�&)��5�lP�5̼0���6�&`L~6b���M�Y�ڷ��o�Ǭ��*�����a �ڥ/��F�?.�sm
/
�"PK��ӐeC�N����P�XD>J)�� �HVv(�9x�k��B���[�w�=��ȏ�Z���B5�W^dF��8�����S���~[RekS�yЭ�tL"�-zX{�4{;��,����t�[�pX���Ո�1G�h�:{�o���<I��2��{+z��9J�G�ǼZ>���M�jw�
���O��	�d�ɴر��B%�.�v��:u�\���4��m���w��G���Y�:�?n���_f^�7�MGU����W(�댻�����^1���J�������~LN{:��E���g�� Pnt/ⳇ�`�u�>���[�e��^���ֽ{�V�����������F�QYHȆ����K�T��yC�Q�[hQ'�)�{��)�x�h���{S��T@�R�q�[yB�J�����J��D��4�W/N���k�Vӳ>꾚�)S������:����PKTJ�����Gۡ�Q�n*�;$�+��Oqt�W���:���V��+�j�9n�OLm�������!b���Z+=@�Sl���D �ќ�_O�r�`�b�����3�{l
L���v��E�j����Kȕi����I+��Ϟ��v5���wI\֚��Q�+ӽ`���6�zG���F�㳫����H�3ϋ��G�h�=��G޽�c�7�E�P*<H�A���6�/�;����՗ȝ9���fg����
Pg���&�65���6�t9��y��W}~�?�� ~�{��`�4?�y_
E���4J������Џ�/���Pgs�-��O϶�d��E�s�s,+�u�Ie�����~cR�N�1��!yx�1�a>�?v��>�CR��D_�=!xQfd�oG�2���2���Z�A�������c�D�櫚�]Wq�	��xSI�k.�c��)����b6�v%?#
f�7�#�2e�k`n�/�5��2�_KG��";P�)�עB<X)r5�,��9ʘ�_�,^�Ę�#Mi�G�r�����:���}E?�1��G��%:�c]Yo]��5S�89Mb@ܬ�?S.���_d�^�����b���P���9/����uТyJ��0�8�h0f���F@����n+,�NQ��cT����?	_l1~4��Aρ&۞��gI��p��c�16wi���n���\��#���5VX��9{�d����-�P�,�]]^�$�T�T�`z��Ov�CD ��3�՜t�\����] ����5�E�t��ѿ�<�S��*��ʿ�a��A��y�'���5k(5הvuTй]$J�V$�j�{Ǽ�n�hnHԘ{�p�]S�)f���elq���_f��w�hk9���1��6Q�����gM�E�8�m���an����b����w�Jnהܖl=�����Dk.d6�;7�M��V��-c"�2ܺ4�v>=C��m���B/�6������u��mّ���s��LS�T��㱊�p����G!��B�����E�HeI�'.s!Y��߹��&?	�愈�+w��%_o��ů��b�/�Ɂ��GY����5f2o���L�9�M�a7��,��w�F�W�ȏ����:�ws��>g���Oyʢ⳼�&�o�����VU��ֲy6�s�_']r�[L��.l&ˌN��]�y�͡��p��	в2\�e�������O^�܅d[n���.��XI�J�>�noP�W:�F���8v�0eT8Z�L��&�|��f��Q�w}���?�\�Յ"#������:���<㿘���5`�_�V$Q��a}��N~�x�u���%0!�5��ȳ�;n^�d��GH.��?R�&�w'�1��^��U;�يDWP�&3Q�~'����,��O�I�R����J�ճϥ����>�ndxu;26e��)]l'3�q�������*��a ����X�s�\���l�U����i��\�>y}�Q�u�[<}�)[r!Z���2�gv���Ꮎ{�CKp̩a����g���-��Z�X/�Q��ǵ�_�&n��6.8d=)g�p��/F���9�8��b������|��,!|M���)hY�����x��<�u�	��z���gA�X��R|/�Bwd/�$׮p(b��{��㋥N��lY<��ao��N��{-���;��v��q�D��x�f��"{x��-���qՃOvz殺��p�1PD�}��g��ʣ�lo\�����]����8��TD����]��'�J_���H��H��Ϧ�Zs�����-�+XF�+C�e��{��̥<6��=���o/�����%��t �����	�#���OU~���@EA�*3�J�ǃ(&���rK=I�K�'msGGW��|����O��p�K�<�n �^&q��c.�8DN��|�r�o����R��pq��x�>:p��N|��H��t\�>�����i#�?��x�"��n ��!J:���˺^�N?�P�2:������1L]�(�q[��Ӗ�o�\���ϡ?d��e:t�%"��2#�f�U�|_7�?Yu�5r�c�����H��9vKr���^��AYxV�0]@��NM-w�^��nUݴ�f��YW��'���q�����+st��p�����{4sn�к�&A]q�J�<�R�B���ZC5���^����M�;Iנ�Y��Ĳ�O��7�5B���r̠���b����� � ���fg�J5q���Q���Ox�,h�� ��jq�%��;Ʀ�$^�8�1\�C�h<����_���f�bJ�6)������g�X[M�l|:t^��v~��w��%'ǹ�2:<�N�q��֯�&_�}Ǹ�_��b/�\��җE_+��6m���?Q�_�[��2P3{�J#<�o��m���5���W3��I^�#}��p�i&K�U�㏶�����s�$����5CG���*�l��r�a;��*�� Ԑ�:�)w��S�&:٠��!�g��lH�^w��m�rF�v�Pٟ���!}�H��*�S�8F�=����˿�9�Y&�:"�^�����{��p��p͵��:�I����7X]?�
G�Yu�Z��$ߔm&�Q��A*q��A�t��4�g�K�k�ی�S��-d0(j�+����//�T��J�F�nR h�(����&�@ި��Mb>#T{o�2K��6�1~�w22s��K���2 ���_��})p��ŭ+��&{�ĪݍWm�Z�,'�a*FC��F�����蛕m��t?���F���v���x������-wǅ]W��hu�u?��.�����G.c>��mC�`��|����D�bǌ��ZZ���<q�|���<�B����O��WH�d��Y�HA��2e풊0Q�j튷w4e�l@��շ�#�+u�k�z[����tkSP�	4g0v�o3ߩ8����M�=�Op�~D�
�ct�)��1�ISOG�8l�ՂS��i5A"_\���@�Jo�2��( u��}�~P���M���g"'���&���OƢ!U)�ChWԾ�}��owq�ߏ����?$
B����A[�!_�؎:�c�J�����$u��������y
'q\4lw&z��bR}/^��E���2�馅�Э����O{!l�<c�����Rs����1�����f���9#GU�)������{c#|�g�"w: �|���m������zL[G�KI<��:F)�3���?2Tc�T��Y�f^��x\��$|k��Ỗ�>I �p2
|�v��	cg�cy�sP��;q�;��~S�o,E����a��NN>DL�"t��W�x��*܈�q�~t|�m�6�����.�A\6�M�6���.��ŇD���������%;���YHn\��Ҁ�,ϑݝ!�� �Pi�$���ѽa#�zL��YvÇk���-���0���~A��>i�-S�V���jP��ȓG�c$a#[���1)�5�گ�?i���.-e�~;n[1?M�����ƌ�0�Å��{�wFg����H�x� ]�X�>f&TW�UjSm`ypT�?zͲ�oӶ�J�7��K��Cou������y��3wT���'�&G��Vq���𴟮.2��V��x�����$���W3�w�4�@L<W�b;��~�mD���DJ����]!I����`��|�M�F}�����,�����ʠŢ�[�Ю,�̀'J<A�|��%
��I��'hǉ���W��D:|`ǵ�+v���|�_��/*N��5�'�	�?|�K-��?���{{h ���D4y��������9�y�Q�걀��=�X�M.'G��j���#��4K���|L����p�rxr����145-� ��V�;��JV7���%�|�"&~zե��d���]���>��?h5��A����J����Q_�нD�*��.���^�H�B����W�ߩ[�M����\8y�l��uT�5��6�H�I،���0M�ci�7|�x\u�YO�N,&mR�0��m��U~��
��E�)S��zU'�����E.><�y����>���x.��w0X\�f��:`\lY㇩o�흓��h��O�	�բ�7��G�����qc�E���@aܯ1��!ݼ��������ezh��-#J~��l��mRKL*>��Z�ڦ�4c6�%�<�8s�H��*
%j9�''��*��(�Wsbb�X9|P�i�ҚX��wb+N�z|2��ʕj�ڤI:v2��73�0]����q�s!�Wz�yU�8�K"�S��uVz���|�c�E�R�
j�4y\|�cG�[յ���P�����BGR�p��� 3fp�d�t&u��,�;c�@[J\��,<q��ۍx��]�|�]�{�λM�����
 r+7fR=���
��I��������v�'�}�p��=����)�I��}�S�����&�D-UM�ӪvڲZdR��Ω��H׻��u�A����'�"����̑��t+��e����P�lΩw@����v/�.�����ֿq	JV})�
�4�r�
ް���LR.Y/T���M�-I[{�e̺W�my뭞1��)_�*�>����a�����\��4ڲ��G�llq�|R>���<��O ��M��d%-`���k�o���ިD�/��������E��p��s� $S��T{���+��!e��,�콡��oD�|������Gl���+v�}�y���)yw|�y�W���r
�zK6��;P��7�j��3�(zhD�E���r,���y���qc�i�*&f�!�C�r�p���.�?k�U��;کQ �����pp� �xo�;�=ض0�]�w����9�� @���;Ӎ��7�M�T���Y�n��r#{���˥���N�<���:利��Mۑ�̱�P���e��oR<#�տ���;ڶn�䯷�S�r�h=G��7�L�k҅��ި!3���	T�c%O%.U<MXIO�h�7&d��x��h����6�*es�%&q`��H�<:���!�f3A;ejF�^՟�<����a��Qg%��T�kUȬ.d�mS���d��l .ž��!�+ĵ@�B��҇$����o޳�2��J���0DF��R=�a^z��a���v��.#��������6���q�{FK}�����aLiNM�p���Y���n���+�gAA�����B�ܞվC�ո�m���p�⺫�G3���2��?g�<V�ғR���[��!;��xE��q�T�Kt�ם���7ji˪����3�Ucm�����B_��:g\=�S�������)�z8�i�I�;O�v:��˂lc�צ~"%`X1Z[���>j�[�a�X���]��|c�{�ޯy�iO��������0U����n����Ķ�	��v��Z�s�_���jx�]l?��KB�m^q�7u�p��Q��L�VZ'HW��}�0� >ݿƉP�����r�l��2�2`��O��g[6,�������i�Z�~�s��-�ga�\���x0y�Cts��/	�/1�]o��)x�ϝ'?i��` �������mn�	M>=_�3e�v����)���jۧU[H�����������6��w�U��-^&V��B��Q�m���q��S�7�x��^��;��Zx{�� �h�y\���čGR�.�%U��X^<��k�^��wX��t�M��ȳ�t�a讅��<���b7\׈�]�r�t-wo*���J�nV�Ǧ����%�V"*�Us⧣iX:rF��1T��ָ����rZq�Wg�Б  ��2{���7)��:��hat��zݣf�d���{�~:�8CJ6��1�>�=�����-� :	���g���AB�q��K�Ҵ0`�8[�W��IDJ��d=��a������	��\��r�D���J.���v���i�������3ri����g$C�R]>��ε�K?L��_B��,���.�#�aa�6U[Q"Zڣ�B����@⵵���sL1"��v�U������
u�L�������~0~OJj�e3'�j#\���7��!�'C�u��t�H���{?��τ�-�_2a��H�|��j���t����+SAm���g�������L��B�?��
�]'���HsK������z�۸ꆆt���{�C�C΃���ĄUYY)�qI:=���Ͳ���/�)�O2��
�_��+���?�
/��������쬠������+�z$�R\J������~�f�J&N�&��?��L����ה������<񎋋{����ϟ?�K�Q������o��_��צMFJ��Ƿ��54�588���������������I���ӭ���Y����< D�P_600P@Mmr�hݵT���W1Zfcaَ�Zw��۳}_fI�T�����t���W
�	��%%젢�gdЉ��A/���q��_d������d�s��`//���Fa/8xy_b��+!�韮�����CU�1M��6��~Pp����V,��蘒���ؙ�h�qy>GI.�oMk5�H����*�������tu��u%�u���3ps�|�z������y���̧��J�iii=�)��%��]�U�m1}����11$,,,o��dee������ζ�x;�'&T�ܽ+hbb���n��۴+����67���h����8�2�����BBB��RR�_�^�AG����#�����QZ/'��䥥��������5���NKK�i4g���srr����G�к,�UޠaOO����20b�Ѐ,���Ǡ)�Hll,����l�	��EES�kkt\�ƣe���߆��RRR���yx�PQQ��FJ�v!�Z[��)ıa���v��RC��㨵�,�Y¬�#@kA---Mư�'�����yxx�vV���K���=Ʉ�cXJZ��ׯ_�����{�!/���!;v��=���S��i�t�I�lXX =��Z�ÝU��	ٙY��4}�.����ڭ���k�<���1|1�;�?RR�{���\Y���n+���65�:<<\}u���	Z��Ey�O@�v������2k�N'L�90���ۻ�ׯ{ E�������_}}��������A���(�2���u_�nD�VP-�Uxll�#���BV�?*ŕh�v1��@�pNo H��Ϸ�l}oӎ��e��T���HK�#p�]3a��#yX9���W��QIe��\]]s��J�42��ۣ��e�@��:�@����^�@=���>h����N��U��!!�
ڐ��!��!�l���E�,����o���	�?�3����T�56����{HB�����n��iim_Y1���OD��{�g�HYEZ_Ldfa���Y.�/++��ۘ6;@�Q���+�3V�oml�C!~ [r�B����|H��A��H�.��2������ /C!��5,,,0�"�󑭥��@� �)-�FK�ή����:�u�+,d����}������������Tj�d��JK9��G����n߆F��j	.��P'�s�v>X|HD$a��Y%0;?�8�^�OL�XZ^&h"�q,��^�t�y�r��kbb�|qv+
�Ȗ��l���`���>��� <6�qŕ�s��ǿ\��gDD �PAA���E>���x���E��$vƪ�틽 '��ň����q����!111��<
`��h@8 �)q��w�����yX%(�����S9`>DT֫C8DDDf3�~��%�\�_��ZY�h���x���V1].�#��nկ���l��������5Q���7"�4շ�zE:�n5ut�������B*W��N����--��L��6Pd����L��FA�$ �
�.�Ä\�t�����֬�zto�ژSF��Y��cqY�|�M�� ���nܸ1o��=3����A�PL���c\�3x��|G�or�3g��\Xht4���WM�u�!��~��^A8�l��
�t��ƈEǭѿ\b��Sd4���z �08���r���Bө���˘t�4��y󦠨��:|�nZY���-&�Z�@gg=���Elq G�4
�Aap)(��:R+�d>�<���Xe[i���&�Tl�}gu�=�� 1�nSMT1^����Q�����ά���~�Fo�Ӊ���X-�yT�[�����Mf9�uk�T�ah�AA!I(W
t��\�~����2�ؖ�!0�Fo�,�W%�+��lE&��B>��;;֙$�_j��Z4s���JN���/r�&M���Q2�d98<��"vK���5]�8%���h�����b�ń  )�UN:�";�����"R��$�����B�Ķ�l��o��l�5�v�OH]S�|Q�o�xB�ݸd�kJz��=ZEpc�j�0�����?���g����@$vhHRR�s�~dB��挗�倨^?���p���\��j;��i	{�Hv3Rt"Nl0��6*oX#�W������f��xnf	� �")��Ҕ;U�����%.e�F�x�J��,�rR(��C �@����{P�82B����$�AzȐ?|�TT�P�E��G <�!#$d7��s�9��.g��4��c�� X�sA���6�92B�˽)��
�"��|��?AWf��}�J3�1;�cd�ƀ�oCO�ۮ����K^W�
�/�W�@b7����#V�ǉ�$#�}��l�+@����S+P"8�l|�\	� 33�⇻�YYY�Q�=�bttcQ����7zT�i�v��κo���ϔ�$Ν1ӗ]L����l�<���jH�m��s���Ў$IDLA�|SSS	�����@ ��J.b�t>Z���'����@�b>�q��l!�.D�i����]�S�B$���D������*do��������{�g���K�߉m졋E" ��^�����.�a��}�X!-PMVN��H� Y(x�?��x�q�-�l�0qJw��%٦�rA\�_�Ft.<7�o�䪀J*Z����nj�@�ؔzG4hB�Q��@��ç}���x�߶��C��+�V� ��I�����x�?%�}J�۹.�'��^6�' *�*�e)���h	/@<W:��A���I��K�Ni
�r�B�d�Z����f����B��t��E+q�����%�u��*ޱ��������zw,�3Wn�ȇB�-&E�ƵH�]�y���bD��:�GXX�%4� ��W��@�DbC ��0�=�N�~/  @DJ��?#�����{O�qŏ���D=}}pT�{��H]2@k/��'�#�A[�5P������7��A`6o��O̿��?i:���RYB��oee5b7A29��c%�@H��\ۨ�;���.�
ظ�Ȧ �qK�����Gj\�Z���!Q�c�q��|G����eJO��>%�������r�U�Oۉ�7�@�%"5��^넧�<�Ӕ�?p����Y�BSj3q�/!z��,��722 f�>�8�5`w�]�=^>�9+oee"ƐI9j/�d�q�4�f}�*تjץ�,���"�DW�|R��J��������7��{g��7�R;4�UQ�O�+ǋI�
Λk��Jh��f���%�\�Դ�I��O����Q("�'�Rח�%!�S}����\��{҉�W�.W�~;*1�ˉ�b�s%��d=*>>�ǔa|.U�h_�?:�755���5Ά����>2�?vV,�zo7tT~�}�엪!��V�1O��~^���.�Ls0O+�|VԌP��&usz� 5-m �."�����u q�$@���A����4L. p߽�dɞc�{��#�:!�	ӌ1������OT=��?$��`�?"ff��}z�u��Ua�e�PJޫ��f�+/Z �F�Y�
� �zB*����X�u��펂*<�����$�������ԏ�bN���;b�5<����g�RXs�~�-!e��(����'''��2�UX��&6�AL'g"4r����>c� �kl,�:���4��A���^E[KG�c��X����P���R��~����K�+8v2���kn!i��Y���2�?n3�q�{q�{q�g��{�IQ���d;���8�*_��`���TV�iR�P��(r�Yx�"��7�Hʨ$��Ր�����:*a�y�{wFx�������v���^y��f����< �H����7�*출��Q������ޘ>_�t) �Hӵ��NN��й�t����0������H/_�g��&rvP'&�;Y�`��&l����Xd��8�����`�` ������d�+IIY��&`�SҨ�n�&���r��IS���k�V�1KG��hV�l�+�9��M���,t�q�����:��8���Ef��������ꪓ���D"�30���GԛSCF������!:\���'��9}Osb�\�����@�ܗ9��_�sO�{1@6��$�p.���=?%�Ӻ�[�RR���+a�0v�5\?��ݟ.Χǻ���]��־����A6��@�Q	Z��FЖP}������Jx�<ռ��\P�������c�m���`�.��������+ww�m�ݶ�v�[0R�M7�=�|����11.�pZ��4��q�&<���p&H^��������l�C���1D�8������o����AÁ����j������QRR�MR5���9d2h'~{OKJ����ȷ��۷�Н V�Ag�FC�6f��l�_(�d���u�=w�0��d��h��f��o�'��߂m�b8��v%��bc;�?�������l��縒�o\���xy�_��ۃ�t��������&g�//.�1��<L������;-\�2h�~C�P!o��in_�=L^R�д�t
���k��C��P-��S��Kq5Ȑ�	WTVg��d~�ǠR�d�����؆|q:;��:є���}�`�5�)��k��#~4�>}����퍍���l�QX��p�I�ËA
ak]��ޯw	�nvo��ת�Df�E}ct�l���9R�sZ��XvKl�2u����Mp��I��xZ2�jWP6(�m1�n��t�rw����h/i��7�)�������o�6yBOS7�+�,������TT�!�˪��!L�U�lnm�T��T�d��������׊�HI%H�,���<��( p�;nǯ���8�J�=9�^�=�'=*`�a����Vb�Je��ὸ�#>�A!�܁qh؀-1 �����f,H��h<=<N�DNTA����HquRJ����;��v㛱Ľ��w8�Z�eV�!!ɀ��n�� bCU7i���q����hI��Օ~�W��=t OQ�W�	�V�����cqQ�3��~ Yє&��e8υ� ���:zqee$,(h���������xu�������&�.Q�_�vy�� gV��t՝�0�����ifE�0@�_�����;�L�W��<?i�>�Lp�bu$I�ˢ�9����;��o����́(t�B��`jT@�Ò�0��ls��ՁSY��"� �f�u:�V�
�W��w�|	�������C�t������恶�Ʒ}	WWW�6�-L��
�S�Ӈ v�m|�_�,^s�$�X���xy�!,������PP�4��hֵIsS�oHʣ�|�Y���-(¸L*�z��M�Rʆcvy���p�䒯�r �����Nz�{�n�D'�f�6Yi��i��R��[dÙ-��gp��>�/\���1��;��c�1\��y,jb�>l�F�y��nk��5i�g�v��j��f�u����N�P��Y~��U�Г��N�<̉ezg����Ymllܬ�F�K�1����Pu�Y�u�ǂ��y]�r���&(�������_� ͏����O��I7K�<���G��N��H	�$,8R4���h�ٴw%}|�y��3��b������q��[I�2��P��4Y*!D��k�2kc�ne�HDbH��%c+ً��3�g�>_���3���׽1�<�sy<�s^�3�w~D�4��h�ĭz}M�x�2�����4�8f���w���8��3a���m�H�F��t�_����xtz(JK�͍H�P��e�ίc�`�?�w �,��'�̘T�\I+�Ǳ�w�Z�N���>��m�R�`^�4k�hR�Vi�R4��"�4�6�[�B�RHܞDD�=�kRXmS�Y�������8����d5�/�u�%�Ƕ}7�_�\�$��>�ӽ8�|e4�\S#j�R�A��)�� ��6]s1Zk�֪��^y����&&eQ�\<O�H{��F�R_ig��Nt���Q�w�H�-@^*��OZjϐG13U��˔���4"_"����τ�M�G�s9�J��R���:s���M�D��r����=87��\���g��������pj���r8]�5�=��=�3g���IV*�F筥T�\m�SD ̮A�����T<���\�[�=�*
~���1�V}��D%Y��g�
獩(��lCb��H�~��2S�H��Щ�����]�����)
Y�Vtз��e~���B�$� +�7��w�r�[�|���?�̷�	�.��F�2� �3+Ay&&&��q�*W�F"�uv��ފ�e�D_H�,IE��^�����\���'�\��k�O���N}`omkK�Gz���a���9�X��ˆes�ː];k�{Y�0�w�'�ϸ�~��*�L�nQSW�^u�lŀ�;�+�����%���>�8����y�E<���O���=�Z�m��NM�T0jeśM��4�*���a����H���x'�>��f��BU��B�1��4W�����o/oc��g��
]F�Y��4^�J�o�l�������g'7z�TKSp����O�\cD�mj+}�'����)c��q�J;���CƆ�0h�c��!����L$R�.R@�|}i<7�_^�C�N�M�H���n{WL/��@�d���s��f[��FN�CG6عkW���kFJ�K�l.`���_}f���~�W���ȼ��0��uH�/�qp�$SO׷��)�}(�w���z�
?�}��#M�fb��<�g��`�2jaϚ�}2DY�d��1I����s�o�&�K=�T�7&���`]�<��S����� �.��@�z(���U�<4���F�71C��鈴O��� i�?�������o�6��'���<��s a�6�k���A�e��D9C��{6�T�c�#���Z#:�`�onv��SO
������L�|	�y���(^a��v����1��������(
U��
���*QΫ�5�Y�Dk��F1���<����;���5<;�F�7k�R�eJ~��* vuuU���=��i��i�������UK��J1v2���cTMM����ЇE#�)��*���%�� �ԩ/�L�˛
P	��t����6a���p;7O��533�rqz���~�f��k2�|#�J����ޞ������5�pQ0�"��{�9�G>N��l@��1��V��??�J�;�Nմ��">��׶�$�;�{6�o���kvo��G	E}k7 �@ΰn��hr:�.y����vi�P99��Q���-rqȞ�8���|�����o̽B ����:�rKF�����>�&��s�A�7�.!n|��N�Q\g3+]� )A���� lP3k� Y��$��Ԣ�.ʂօ��lq|(�`�4ȸ�J��p��:ُ!۩�Nmmm�>��_�e�n��P�~l���g#(Q�O�>�k
��eo!T��*��z���(��G/^�S��\��i�q�*��<e�R56�d\�o}E�6QSS�kM#sn��|��5�t�$V3I��<�%�Gzz�
���w��V&������ˁ���G���I����F���Ȝ�c�N}D�>�  Ѥ0�P�!+j��5ccљ�殦�Ǚh�6��b)����0'��'�so�
����/�]Ϟ=+����և�!��%j���F1�e�;��!Z8߲��6E�C1�m��C� �����̑��h�r�#_\��xV]�*��jm���E�j���S���u��Y�H�W�5�秉������X]0a�P����8<4T\��7u�f*۶��Q�l��՚�A�"G=����Y�������(�I����OB2�q|�k�7m��45�=#Z����ː�x ��vv;K���_% j\�P'=��tܸ�:=*�<^�dّyc쌼}a�X��טV�-�l;�rY��]����s�t��'�O��ݼ�m�j�d�왟�fU��A+v˵ �h���O���b�a?~��I[����.�x��D��⳶�������ަz�.4|��0�B�|���v
��0,���X#����&���f���p�ib1��B=`V�P�_-)*�?�>�+��2������a�w8��	�g}hf��۫��m��O�2I���sJ�����QBZ�M?��h/���rJ~�E[�κ�4��������'�m>�^v}�kԛ^^u��隚:�yz�H�IeK,����ok�Q��`Ȣ���Z9��_���>�H� :�M-�B�WV������W�DЮ�8�Kt�X��G��/��5�>h�Ħ��$�oBK���(���N�|������BX���DWwa��tB{�e�CC����Os�^�O�� ($��'�!��o��O�U�����{Ё`蟷�%(e�����r�6���S��{��%�3#����5a��ZJ���v�!f���1T�PU�U�u]�Əq��F�(1���x���.^vm�qvaA( 8�7��OMW2�酟��0���3�9VWW�ἜsW�z��{�Jۻ�����Y� fEc�c��j�ܫ",$��-\��FK�tuq( \
t���A�%s��/<�rT�<�����z@�j���V�lcmpo�O�>>�7�|�|Ｌ���v��ɽO�r�榦k|�����:9�uwq�y�}����/PTB}���^ qOV`ۖ� ���	�����퍌G&3Fo{z T��X_����漕U��s�a2gNu��>��l:�P������<h�uC�Omv��m�ܜ�X���ma���1��y��/jX���R0_qL�(�t
�!��ý��au���X�1.�:s����vq�����h#n�˔��bc8Z~T�j�+�x��-���y�`�	% <�I|�O=G�1���	���2�#5�t�f�m�3��W�@IG�d�+��~�W��"�<�Z�e/K��S�|��. ����*,.��D����K�姌��)MrB̇��d�q`��ƴ<;e��㳓��;�*S/EY���2gJ'T���,,gȢ���S� ]H������#��{6M��1:6VHaKjW��;(m��JQ�����7�� ��@���被n�ɳD�&�H~^����u�p��e-["����|P�S��Ah��t��Y�q�B��
\��Ŭ>���,w�������<]?�/	���8fD�Ѿ|�!�k�����w���O����O~�����hoWur�O�$�o5'������#˫KKK��C��>*J�G����<E��h���@W��/��h#��^:�<�9y��{?��^ڸ��R	B�s(��L8�e����x��~q����\74\���6��b����yR��"19��ܵ-�N0Ѫ;n�z�m���*Y�.2��������S���|1��%�����	";�y���y[�J_����{�,N �~�.���3?&�����ud�x��s4ٰ � nkg�D��o4�ܠ�xf�4�W �]�i�o �t�Y��`(��`o]�ZT4�vW�^;�$��:tC%��V��EE��([ܯB6�#̔+D��,*����j#_�f*�^����_cS��S�;"��[�@%��_��ŸFU��6���3�$$`������H�v�f��5pc�����g��
E�h+O<����Pm�4�H�7F[�`ᴐ' g����Ϧ��+J��İ�R��T�:��~ƅC�`z�U���9��|� �C���g?�"˵u�z]ʁ��H@��)a3k�� 9y��g	�\��uc���H��W-䷉��'h���y1�DU,��a�?��m?5<23'g~V���]gOլ\����Q,y����|��V��Ͽb<����Ν;� n�.r��Ç{l���ss.��	)��;�O%݂�=nR�N+7��%�����@Z��$���Lz%�򎓝k���c��S�~d��&�PX���]��fy��#��h��;�����O2<�+rL��j�=����kܶG9ܵ�Ԍ4,�O��Rn4#*�~�^���
���D�ieS�����܅`�n��5���Yߛ�7�7Ҕ��;��^�����_�d��O�<R�?�R	�P�}c�&ƅP=H:�A:P4R��v���т��J�1&��]�%M��jb"��E�K#\��c<>/�v	C����k&���BC��?-�,g���rbGm���c�w���v\\���=��v�<#C$��-��U��y<�;��ˊ�����m�>77��qc��߷s5*x���
aF��,Ot�X�:1�x�:R刬��
ޭ����_dѪ����q�e����׎#�ra��eD��U1���qy�l*E����Xk��L�ɫ׮���[�x<��Q��l��֯UA�I6�ϛ��ǘ���w��#���,��㾇�i���
"�������%�"�Ǹc'l��JI��2��n��q�BU�V�Y%�E�7]d޸ߙ�����Y�N�b�	�/_��d:PDH��u���e�����@���w~���� ^�G�l���E���ۜcn�P ߄~h��2�
g���NX��H�%���M��rU��s,-�T&�"�C&�?�lQ�lN������_���m�!EX��Y��rb��rK�E��k�V�����=J��)n��e�1Kii��89�B\͛��&�������o�v!��sc�J�5���M�\�ĭ�ׇ�^5,<������DWi���S5\�X��w���.�}I͆��111nn_�2`�~�}O�MI-<!+3�1��鴐� �O�2j��%-�f]� �ʩ�f��D�Dʛ7W�/�m����
�V���|�*��`��<k��ړ�и	sp�xG�-�x�%�5�V���WG#��J�����0
��K>��7��i�ܘ{/"����ҁã-){&�ʖ3`_bCC�:1%%E�dq�3Xݖ�y���P�׌���F���m�����k��'����=<�7��a|E^SJ��3�I���2����~�WKu��ڬ��wbI�B��vz��+���`%�`~����d�]��8ت.ޡ���TpL�uI�v�5,Z3<T5���{`P�!s��JS��o2E�{f����?�������K�z��4����k�N�e��",�%��~��2�`��7���V$1*�A�������_��Nbb���ai�{d,ha��p�G� �q���kVa�3��%�a�Ex�P��|MQ�������S:P o�I7,/�+i��&K�Ƒ5�f���_�� �m&md�Y��W�N �J��X�N��l�v�����@�,p�$�VVV׮]{A��ຉ�Փk��*�����[+"ҭ� (�
��ajf����r��ګ�إ@�ځ��T*������d?r� ��Nt�[U��"����C>C\��L��Y_=�ptQݗ�eЪ�[�
���:��l��[��<I�-4������,�:�;a�W�x���x';2A:d���09�	PT!k����T]��&��$� �?�<:���7�8�ک���6?��2�#���ES�/����5�k#e��];w�� ӑS�h����Wd�����<��u��:�yt+??����j�����t6b�5�� %�$0���x!�a�O"~��k^Q��j�%ٺ1�������)� .��Ǐ���g����:��r�F�s��d ��E&%m<��iql��V���/Rn�ğ)�B��FZ�*�����'y�N�U����Pc'K�spT��.ZƂٷ>=K�K�Ka䡫
=��I����CV~�4�
:��E=꛵C�#�f���'s��Q��P���ty;�%�ԛ�6����� Rlͳ���un���P�یx<~vUO�hZZ}뫓����)�e��8��M7�}�|�E�S[�����	42�� ��򭦄W���6'�RZF��̓)0�9ҡ&gP�6��?;��I�=ʥ@�Ʌ�S������%e7 �1m�c�V2�����G2�� ���̝���2IH
����̈�T$���,|$��G�y��='����C�$�yT-+�8dE�UF�܄Q5A�ֶ��X�Z���	o��wfW���sP��g8n�CI�,�DyV�i;V����k7n��%�H���EB6�Y��̙�kE���������� 1z�/����Xc0�<[̼�����dJ���	���q�^��jb�hJ�[֧21:���ڃ[1��jVonc����M$��A#���$Q���mp����W�n F����n����=`�e7�|g�:ۂ�������y���x��Űz���s� 	5(�d��y.8q� Td�%�8�t���}�T��W��UTT ��eff6�ã��W���HÅ (G{z��� �}�i�L��ɕ+/^�H��v��~���	^�m� �Mo����[�����<��2
�kG�s�G��iy�� #Ҟ\��T|�F�2@���S�13�Z�VZj�l9�����ya��|+��0^�n�I�y_&Y]\\��я1���~=�G�b�(]]^pC�F����l���?�!�4UC$o�xjPZ������N�w��r 	����d�djNN���v� ����:w�X��ٟ����T���G��3�L�{��J�H��uXm��G���V&m�O����B�9zR��,���?�]������(#��]r��n�-�V�}��:�!~���fr:�,���`>��4����8)i2�Bu󘕆�o��Y��Gɻ\9-x;���#Qj�0V���ham{`{Gǝ���)(�OOOZ'D�C~'�]߷�٦Rq��O��e�p��0[Ȥ`T�K\���9�� /�p�j�W))����K8*y�V�(�t��5���5�����/o%����6l�[ ���ȏ�Թ�2H�_w�;�LM�G��.X[�T��0W�j��u�*�h��+�XYQtW��Uj`2����E����@��[�M��j��i����?R=w.�?�x�˩)�f����Ic�k�.��s8*LRy�$�m�ޫ�H�~��8#��߱���ׯ�+�����ǭ�q��5�������,�<�S��5#3�d��̞���!�޹S�N��'~�t3���Y��2�����uq��J�,#�s׶4���]:q�D�ZW�J���toy3Ԝ��ߠ���1�PZ͈EI��0"r��-?���L7�_<�������J��/�vP�d!@�q�D��"D��9���<g�����U��]�1Ӣ�?��5㮍|����zO ��A[��,tW��i~��?
��8F�{�}���ȸdm�t�I���
]2K���g�x���R�S�+[�к�d$���r`�0����{�E1�I{x=��b�E˫�]�.rJ�W��rB�hok{{�d~�d��(
�9:�^*2�<$znv��u�C�szQ���K��	(m��ã�h�� ��.n�S��_�t��khx����u�P��" �ko�B3i�O"�˼٣�2��R�H�Ѵɻ��`��v���|YZ\]*���<�ӷm�[~���0�vf��V�"���֠6��Q~%:�*)q�z� y��]��u��̼L�pe��z�X7'� /��E����#.G絠�P��'D����0I\S �4<?B�J�TRP�K�������F(��5^�tY�����|�m��/�_O�P�TR�0�ͼ/�������cq�HkE�Z���z/���T(�5��'�4�]���޿q���Ƿ0u�!ވu%��V�ʬ����"�D�S���q�K�J��]a���]~8ܼ��(22���w۶n�oj�lR�'����9�=��އ�y|Pt?mN,%A���V3nm6�ҧ���� [���O�Z'�2���j�r2.��lkk�joo�'p�G�E@W�6?"�y��Z�F%~�7 :��!�����ф��I"US�h��0�t�wX��T$It�	��s�Nt�dbb
�ˢ�L珁����8B��@�Ώ��H���EFFƊv,� ���Js�ː/Z5c��Y�
j32���.%*���#���_/E|�"
����*��33�3�nRG�|8N����V��Ĩ(�ߡ�ӛ�u����׊E��w5A���K�VI�{�:�|F��������rH��Y��D�L&$�C�rJ���;��X<^������� �_�5.�z��S<���Uh���y����ge�N_�.�}���d����JC f��8�VV����*�z�E��Z�f��[�?'dG����WRS�dr�?kֳe�H�э�t�B� ��C�E@�Vg
���l��^�"[D��-�#��#�7��
"+YOWIiIA\.��l�6�n^R�G ��"�{���S��Cm��a�ho$����Uc�=��j���d^'o'�'!J������Ĉw܅�r7�9A�D��Ob��7�S��b�r�`�!����߄�����*u�B�-X��<����[3��_�p$A�-���%���T����߿�wm�N4R�P��̽%�T:u�X!�Z(���4�}D|�0�����[��I�3���n���g����؜ȁ<"��&���������v��0�k�{�؛kt+���L�O%�-6 �n��v��MD�$��+�=2��\n�<�XeS(�(Z\\�Gy����)�$pӤڑ���/lI��&tD�"����7����tGv�/��!��-'��?��ӕr�.񗾾~o��0=&c��>ܔ�:l�8�N�8Jb��L��H���;;�3wU�t�p���,��L�q�c2��b�*'3�Tme�?��o�F*�����~b��|t���׬�	]��~����\]�}�zK�W�Nxj�ߣ�O#����e���������t�>�*�:���pi���į�`�j��w+�>�l�y���=_�-s�n	{��N�'���p�������=(�rIA�
��wT�v��K�<ʀu��P�e��ߌ�0�����Ţ���nAgG3+�!�R>���A��g�!J��Dhz|�����S7d�|��,�)+{.���G�*�+���u��9���L�g�X-�"H30�(}at��K|d�����9�M��{˥�:k�/8��2s�T|l�?��V����]��������8+]- P�4��*bӕ�5P���Twz�]S��X����a�s���"��G�����|H�2]�b<j��$sJ�u����
rV������_�
�i��������Gި���׸ty+���7f��C�ִ d�ݩTѽ�#5�S{��o���IX?��ԖJ
5�'L���O#�,�Mܿn�S1i;�ѭ]f�!Wݖ�>����7,�gr/��y���T4{����"��B7����D�rI�#i)V^Ia����Leӽ ��թb�	!|F�1IB>)b#ǚG�6_����g;~�|B��4y7�E�~L6��R�󱉒���Ns��ň
w��c���}��N���8��Na���b����.�_\	R�O�KDߦ��,p��Ɵ�lM@�Ո*0��EDD��H�6��6����8r��zP:""�|am��V�`�׎C�{��8�f��jok�{�����W뎃�{5)���!ؕ��Ʉ��b+r2F:���R�Vzt�ܼh���R�9�{e�dEy�`�ϭ�m���t�Z�����p��a�ӧ(ss�,@l��Lw9%%;}4k�+�9�Wi8� ���XsT5y75o	#�y�Y����}F��r<y�$"�冇�����_�b�M?0����-�k%����6Z�v��c�_&�	%��P�Ge?H�68(��ݱ�9���R�l���ދ%����⛶�M�.����]n�o0d����+���S]S��V�P۰��\�Z��8���vF:0�7Bm�Z�d9�U�VY��c6�\|܇Q�a��T�O����^�L�,��.F��S��z�q
vA�����].�,^iwo�ڥ毎?/�Q$��7�R�G���9��y���P�8�����[1��^I���۸�3��LKRR�w��f��fs���x���5�~��OcgD��3�r����۷�.xe��ҽ����hr���۷�>�����-��d�{��P�ڑi���x�b��9:b�i>׸o�ԕ�/}���h�v�{�e��wiS�Έ�w��e>;s�y }��@V�C�ܮq��M�B$�����9��K㓲�'��Z5mt7�Ȱ�D��p�]�'�{��e�v���A�Сsm�;hf� 5�(X"N��U^ /����C�ꃈ� :o��=rFH��w�5��^챍��$H�$���L��u��������'1� ��A�����
�l�l7�%�~i򓄄���e�e&�����O\��i����pllR���r������亽܈�N���}m��4:z���;vިʋߒ�_etc�#
I��$!Gl6�3/ڇ�M'�|\?z$���h��[�������9R���e5+�k�`i���!���_Z���4��S��8i&�ӟ ($D
�Ç�y�EOE5���ngMh�1�0��*�H�+��40�',A���k��7/K/�CF�իW7QʊH�~�����,��4k}��ݻ�NMCc������e{D��9R� n��c̛�N�#G��]�V��/(,,����s�M,����i�X4�lиGg����B���!UA�5v���Bcjj�:t�/w��y�(�Y_;d)�|c��޽����AHH���yO+�&��ą�KBZ�х�� ����b�Y}Nl#������8A�O��!��v+�V��zU?]���]���q�QQQ�PZ.+�����;�<�}Sa$)-ݶ���- *��+��02giɓzO,�(�<�����c5d�����Tf�SoU�>��^;�JII}��L_ ������kjv��:L�Y���z�{{�SC�=oĈy7Դ(]�4��)�`��ꊐ=�+K�0f�~+�bW�߾HF���GP���5��q`�)ZC�dΝ��ՠ��U�aE����E
D���> �����i~P�a�^9n7E��qT�2F�����%�G�86�V@lKj�A�:���w;V�����Q���j&�NƷf�ut����v� ����Q�ƌ�o}Dqpp��C��MǸ��@�9!#��&@gWWR(�r.>���fkM��b�y� ]"ȿ�P��?��oɉ��n��5���I.Q��y�e���7��
E�8&f~?2n4/�=F�5.,�]�8Ti�4�kj��������H��߻wo
�"��x������������ʪ���b�̢w����qjx���w��.NT�~N���tD��+1�����c���I)*����S��xl|��c�;͠��duy�;��kUP{���i*��-��W��~H &�\��H����'N�Rsqy��� �7��Z����B��4���^�t���F��0�[����ȏ��r��t |�'m������[O�"E���E*����(!-��\�n��+r�Y�!�|�.�SVV������w���m�,j	�g�qp�hA� �*��t����ƫB�`�Ksss� K�.`0������`c�/+ڑ#�V�����)	p�����'�j\d��X�KKϲF�"a|�t���Φ�G<&�
ZJ{z��I�N&�OCC�3�!{�����$��t���\$ާ+(�/��cs����g�!	$a�Q���22n	=�NM�X�g�؋��E`�
��כq��������PkcE!��<����b}t���!,A���k�ܹ3�'����	�S,�����'���<9��b��ǧN�jjj	8����a'�Y���{��in��E] ��-�L��:���#�-��"}��m��OZ}�W��VQjLJ����ϥ;����e�r�Kum�:p]HS�\�VE,���h��(��vgΛ�w t(������k���Y@
����H��!Kx-�:4G{$P+��3�,��ߟ� E�n+�H̯
ڣ�i�0a���DD*�����DB�"��~�����@&j��}���Qd��o޼y2,�Ғ,����/e�ŕJ�};����
�!)����dv4l�Q��>x��_a
����$eV�/��\��b���jԃ�Й��Z��tj�}
|�����zIU�Ȑ�E�?^�J�<8�OFVE��
0��{�וR�������y��%�7��{���e���K��%O�%F(�?9y�ٗ)Co+�WUޕ��&�tkC���/�jb�'. 0��@8A�f9)#���S�S�("0.�k�HKN>���M���n!((�+��߂���횶vF�5�8���Y ��{Q����4w�ǚx^J�]�����?�ܤ���o.�L�����2�`)$ pB����y)i������������N��r4��x5X
Z�٣ȫ(�T)��em..��c��6�>���O;>�u-�SّR��p�o���!ix;����ֶ�~ z�I(I�O,�!>�����WcD�@q���O��"ty�����g�n������U�[�˗�1b��g��Y��Б��Mr�֊{�1/^�O�p!��؊U\_����yd��c�������3�?�"�L)�s�������ove�[˂���g���R��s����GFG�>2G�9y��,��8�u6vv���aV�������fl��o�`	������_D�N������USq��C�bb1#�^����
.�z��`mc��|}-��4
&4>��$���̢Xĝ�<�� ��8�&�}hp�W{����U[;;;��V��B�Z�K����\�.S	m؀�"m���Oq5?�uZ��u��^ּ��4�k�F��*>�VA��GC\rqqዾ�<yO+d�r?�_�JQ��1t(�s\���*�,�W*�gϞ\~�(3��,s{��LW����9I\Lw�7nF�o)�t���_�PL�E�m**ߚ�|!���̋#����3��Yh 3�|�0 Flg�5�7�wre���DZN�f�n�t�B@I�̾�%~���5�;:�~{J�;w�w��λL�;O~,ZM����c�:{h�X��ė��� ���sʆ4��	@�R����8�<	��C�U-,RVF��2��JY�\%�.:;�_��iЭX�qICc_���M=.��g��`=|��CjzzÃ�"ŧ�{Q��}�'}���Z�����������	]ho7����o�m���hvm}m5!g�j��ٸ�z_n�q��/�!L���l�;uq�y����G8�\&�Ŷ���R��U��N�ɜ��x�?u�\9��X�5�n�Ժ�sQ���Z�L���U���ڭ�"��O�KN�,j��9������?��.I�z������6<�����9Y�`R�����O���64I���vmxc^VXX8	zh��L�Wg�H-�j2�-����!5�%���G�0�������d� 4���5�k���5��~o6��퐼�{�\�a�4C���NL�Q�5`cM�gy#>��h%���B�U�a憎�ܥ��;��3u���B�r.,�`��/vNc��*:���[�1����g�e�:�B�-��W#��La�l�փ�е��*e�K��X(�YD1�Y߻x}w��6�'Q4�p c�H��/�w�o��f�?��c��)��W��Xm<ӧx��4��]���mjI�B
���ĴN1���w�@C��4r�znPZZz8��w��ho$�Ы���P�b��C�/W�~+ME����毎����j�\�����t/��Ǚ�N��}e��C�_���LJNV�I��~�,��� �������u;j�<�t|ˡ��8�-��. ����i�_��y�jj>&9ď�2T�!8,|��Dk3r�̋/�vl�N��hD�9��x�ۻ�����OmB��e�r�tu�6�E�u?���xP ���wy$�.׹eWhj���>dNs�;�c����Nq���W�z��� o�>�����]����4X�֣`J��]���T��ϖ�֝����œ����.�_��̀3��u���h^�MJW�9�������_�.�� pw��𓗑w��WI�-746�&y7�O��9�O�C'ΫU��8�����fh|��6C�4�i���8N2�j�K��J����u+�{�߲�H�guh��ДC~�����ŚC.���qMO�
hU�_ޘ�)�]�3^���'��:cù�L ��&�h�c��+ĕ�F�pJ]E\Ԓk��S*RՒ��V^n�,E�4�K�����Y|�	fY�`��+W��o�" 
���JYfa���!���G�(<?��u�~[l�N9ԟ�n�xy����!j��&�"��MO?�]�W1C��[�$���>K�f/�����AJy[hߓ�w4	�!�K�h^Gq�� #��O5�����c	�:�G��s�[����xYzv�'"��7-,���\�`�H{��� t�����e�};m��ݸ��{Q���"���v��w{�RՀ��@��gfBzz�E;�h�*^��7�}e��4��#<^y��4d����V�Ϥ��X.� �������k�3J��Ϥl}nȝ|e�E�Y|nY|�0ڍ���'��{������������N��f�.#Me�@J��-�͑��W�k�r�^ig4�
6�4�U��d�C���F����%�ѓ ����%e�ͧ����Ҝ�E�'�����P!����.A��������`��ꢺ�I� ��"	�����������cp�g�l$��+R]@~Ǩ�4�D�����m�yOd]�����L���E�a��XlJ�<h�=)�m�,��y�y�<R@�0/Y�����G��6�rR��'��>���`�7�K����E��$t�H頍f--ynl-��_�Ԍn�m��|�ʹO(ɛ�@������U���+�G���Z��Q�h��/�s/����]��JJ��~�mcG��y乶}=��?_�S/S>�{#��ٶދ+((��k?�D��q�G���sR-^�BڮX{��Y�Ssaۂ0'�[�F�_�st�};��%�9��"
�j|n�@������iv�-����$5<����x����7{� ��q�F�r�:�=�x�V���j�V��zZ�]��c���]�H��J��"C��щ���8;�1AV�,�.F���7����!4��I�����e�#"�b��sd�
~zz��J�@8������
��&s��O�yN�P��}��ۛ�}������/�N��,�^S�y�r�����}�ۑ����I3�=��e(�P���O�۬�1W�˗�'�"4/8!�~D�/_���Vde�on�zRl
�dI� f�o�v��؉�V=���G29X��ZG ?`�@�k��.�y����l������E�$�:�����e*Ѫ����_��͆o��U���L��=�������� Vz}�N�ɦWf��	N|�h��N����ݓ���6�¡f�5���ڐ�`mD㻻۫��>�#��Mrs�sp�;$���^+o:kh|܏<w���BDH+��ɫ
�2��ow�s��'���222ttu�41$2$���a�1�K�m��\WJu��>y򤐏���sήx,=U�\�S���u�E-��
Y?��`��mpx�}���������r}�D�*�?}�d�9.7Y�^�=��u)��9�����!�D�k~�������5�q���g�5���H��<�P���I硺03�__ ?Nٌ�֫����?��x[:q_l�/�>��Y���n��gF�M###s(-��bO.�dQ���~uq�W��"x]W7h��T�A>��B,{q�ܹ �>9^"�@�C.b�s���h��r����o}�o���u�s4�bS��N�ss{�����-�哴GE$S�)[&
�!�dm>�F�!0�<ҀN�͛�U�`�s�&�bii�"����*L��c\`�x����j����8�����o����"}}}�3���2_�n�S[�93B,�]�ѷ<��2�_�����H����6� ���S�V�i�p?>y�_�T^����U�"���0N�@s$�?��{�0.Tt��y��Ok�z	�4 U�Tʖ�ɴ���S�:urs�����yJzl�k��C!�̾����9�q�2��Kc^g�
��ȋ��7���s�?�C�=VX��(�� ���/{��m��~��d�'��Ĩ�8ᴴ��+Gg�24⾵Ӷ�0O�||�}��-��)]�v������h2�1`�����F���Ah�|�X��}�wڪ��|��x6�>4����H�Ƽ����@��Y��E�cm�`xz2�}m�̹�ź���S�ϳ�/˯���@����a|΄pg����|ۘ7�ɓoJK��i��K�������0����s%����oIB��=<<�@Bu�G	YA�*�,͆��4]_��h��/�_�Ư��J :5?�@& טY�k7'z��
"���-G?'�9����V��l�L�%��\�04�\XV�,0����w�DXC�XI.�
T`C] �t���ڳ;�]�.�=]��Y
e�	ĒL�I�:)��)l��yG-�����q@��]�����pf����	>v������;/iiM��Ŏ,vi 
���-��+���e�b��/��[P���o���x����B�!b�]���0�Z�p��y���WIۃO��:��	h��O���۬o�Q��(Օ�|Y�}8bW������z�8��@��]�bif�'�xL�N���e;y	R�u�8�����.S�+P�$p�
,�]��A�yIC�(r�f}]�h�,���yL��iCV����AC�ӗ���r���;���i��Ou;�z�\�t��5'��dQ�h��鋃���*Ct��`^���Ni�p\߾{��k�0m�B�ޜ�i��E�\��7o~�����X<��\(�8�xQY~�ԏZ�H�t��3�~��!��r�s�~#����?����%���s�"�.]�Lm��Y�׸�w�a%"�v֗-�(�/6Wy� [1{�����Q����FfA�5?γ�}�6�����d
�Ү���/��Ƹ�ñ�U���A|�G���ɜ>5�|*ÉE��CCC̙99�_�=�s���"g��<ʝ�`K�u3o�i��Խ���Hq4�ˊ_��5������-�黺��U�b�!�v��X�,��i��_O�5׮��^��F���^�oyS��NB	�}��1w����Wo>�.U�o�
�8Sѯ`��[��������-DHSӨ6s�B-R�(D����>H�mSƸ1�܄^XqYKK��6�B��8�?RC��][|/�!�c�d��m�2�$��p��Ȁ��װ�7�~\?_pB�X�d��?�RΪ1F��6�(�F�o(���˺Sy^[\];κhebb�2����Ī-��F�/�c\����;P˅DQ>w�ߧY����_��;#�b	�tz��t��S�ۋ]���oɭ�'Rj�V]�+p������~$9���T�����HR,�*�G�3\d�+~}5G��7���vq���P"gHMK��nd�z$iQ\;8���;+���`�˗�q�.�]h��O%ɲh��w��P	G�ܚ��b��2H�H,ʇ�=42��|O��W1������;y	��L7N/��b��Z��~�����VQ	X��<���v�{�5}�. I�L�B�$�L�#*����7�$���8@�c����)�M@:�5�������|����mʝ���������T�b��a�j��J�-)���@��_�F��7�Y&F���v
���t�)��ĸ��r�)���WL-��- ���{�jy�.�ďX@��\�/~�`�R���f�,K |�[�E� ۟�>H�ծ�����m��$�`: ����X�ȒB��|��^�gϞY��0������jJ���\}T�������(������ҍ	�"�-��e��HJ����t�tw�tw�� ����u��z.�>��޿سgF;��:+�Z�y��~p�7�|i.��~�E��ƿ��qٕo��|r��J*nJ��Iq[;"�{��s�<���*��M������(�@H���D�_�\���	�dk�dv�^G�Z�\؋���:ת�j4F��vMۿ�Yt��K$�ŕ��h���6{�Ĵh�o^��4��1����x�y��&����Ծ�M����⼛�<��δ�+��]�*��7�IF�}.s��4�R�{N̛s� ����`w�+���2%*k��^�ay\�L��:`z&&��$k��8�ͱ����-�~�����{���$N�/_V��8$z˵��,� �X��Nutθ���lw�0:O~n�������n1+?�i9�h��Q=V������B�me�BA��bdxx��p�	d�`ߋข��m�J�~��\�w�q��.jJ��� ��ms��������������<�G�;���QU9t��ݢ����Q�{��$��e���n��w�	�E�\�t�&�p�\��D�Մ����l����8R��j��zC2N�Ć;l�������IH
xV��>S�;���X��d`0j��\v���� ʗ��n�O�n7�LAU��x:k�����i��Re�ot�.�L��B��@�:Q��b��q���CKn\�=�Ac�D	+�v9���4��l
x�U�Vט�$a����t���5	
x_���ǉ6�Mf�Ӵ���3������ߺuKp�"R;g��1
;�i�8�Դ�����a:��`�Y��og_����65��eo�y&���BJJ��$�ኇc�jF|k�a�ϐ��8���3��rW;ށ"H�Ծ#�A����u�E�;w�|��3ߧN���o��	�4lڵ\�	�OL<��U�E)I:ن?������,8HKK{[���!GѡX���љ1j�\�����@���m�q�n��л�Y?Ֆ��:��o��)>YPHH���fB�CK�8���Б����ˆ%=��I�^�X�h>�t������m�lm-�7�J���yo���u&�o����M�y�������<���<.p�5�ß̢��Wf�y��`�ǐo�m`9�p.������D�@��-R���ֈ{H\��إ�Lw4�\�-��d�[ԩ���.5��J�aH!�`_�ĩ�|m�S�r�I�,!!!a���j�O�!�7��kZ�Զ���'Vu��f+�c�
��I�� �ށd�U���z���g#��=�!
Yz؜Scgc�7,l��2[�+~j�!�7JP�m�uc@�!p�z�!���\h���%{f�QT��a۠g�efզ�ׯ_z)�{6�x�,0���BB:w�+��G�����o��h�sj%:R=��M:-�VQ���v�T�-�u���t��A�����ϣ�[z�W�^L�;��w; $n�f\RT��#��',��|q*P�`dQ�r�~WTh�:Ȧ� ��`����a����ʘ�����57b�¬Q�R�t"
5��� B�y�۵�* pr�)�AH�r��s�#:�����t�VdED<E����8����u�vC�̍ݽ$і%]��q$frz�C[Ձ8��E8����ѽ��
Ix��:��O�SĽ-�"�:=�@+����>z$K����z�sT�P�=����?����7���)�W���q��l�3����iii�jeG�<yr�c�=�������د��*S�y�?]Ȼ�e�1ӛ+�Un�؍e���~�~��u�>#1 �ʆ�t��i���qٟ��������}ͳ'$$d,�q7��hD�!|9������&�+���E[�v+Mj_!"�G��G�n���p	k�jk[�0[��#_�J/h*�{t�g�6�M^^��b_n�;J�[$��*= �u,�쯞=^�*j�XH��l��{�E��lV��>K��JX�6�Iq��R���{!@j���dh�y�`�yk�l��-��9G'�q�M��J &y��*q����E9�xI]]ݗS�	���i��850���G}�Ap������Y��k�/�WCX|�=�_�}�"
���,�����y�}~]��,53ߩt}{�<3�Y Ƴ��#t��A���,)t���AG]mlX���û0��t݁y�h�^>��Jy빔��`ɯ3���馦�PYIt� J̏?*�N�s˂%�f;��A�k���Quuu�dBCty����'wsU@� 2d�=x��_g����!W
!�����"���E������X������o/RǨ>ܕ����n��AA4篋�E�@H��χ�E�-�^ۯ���m�o��[.�D������b�f}0Ͽy�w����1�	��S�o��λzno�R.@Sz��K'$$|�
��.[<+���i6^�戳�	K��� xI]`-tuE�#/���J�3r���n�X��"��kSr{��I�ݲh���S/A�.�0�8t�Z�h҂�\�ל�@ ���+�;����>�����
�}�Ǐ�+ʋ|�Wj���B'm1��f�Ny��ո�̕YT�k1Ĳ�AZ�Ha�XrN�/�ς���~��_e�Ҁ8���j$58N���53��Nh��S-�󂘴���sA�z<j�/K�¸i ��ꏇ@���D��� �4�i�����1�����

����� b	�7������5TM�.��e_�+әλ���An�577w����=|���OBs�� �Y���\ϐ5�c�&��#.ct�7�����a��=P�g�cw�:Å�������lb�����!RQ�����;��Z�O1f��F@�e���ht��ۣ��;����~�������"�Y�s����Em9A�S1r��j!2%<�H#�&@L�I<<�6����U[���5����s��F��C����;���(��9����c�>ѡ�%@f�;��k0��!!YLe�'ͫ;�ԩ�wsS$:�܏n������m,dgg��*�Hp��(�I�'y�k+�-�u�fO)���\[��w�6x���N)w�=�.1���ʿ�O��>����o',i�[
(�DWo�r���]�hw���������]$"��}���˭���k=j�t'�v߻rE��'�k�Ĝ9gǖ]щn�{Z��{�x��BŴ�M�^{���׃hG�$�_��|���f��>�����ü�h�� ��X ��=��y�����O�8�@�&�bu����с�>S#�����n�S���A,ӫ��h�E�\�&��S �k���-�a�
ہ�{�W���a�|�S�F G!n�t��.?Rt�����|�F���O�hg|��������eof�wJ��s��[�A��6-���R�Ac��T�k�~j�S00H�� ����"�,��{ ��ƅ������ix��? ���3Eװ��.s<�Ob����Ak�j7�Q4q���8]��|��5�r[/� f��P���� �U�V}B� ^�KRV�����Bz�P	�MF�3�����������>i99!mqQQ/��7��r��[���o[�4Q���d`�-�w_Yo���JУ֨	���`��M�<V>�L��
���'��r!�:~�������ԡ��&:�� 5���˪���-��������������L�x�y������pϝ������G�zċ-��w����^]]]���������Τ�����L�����/0��4��E��\�KU�"?��浪0Z�i��p��
)E[S߿�b��L��=F?n��{�G�K��Ʒ�Ӎ�z#�Ή��.�	1��Q��G���?��R7�|)�A&����h@#�9��+��ཛྷ�Lѝ�_b�*Ĩ�&^<�],���\�vG�R��"��9glL��vQ���&?I���$��AL�7���C�+���R΀�����Ni{�B�z��5�.۬���v������#�i80��m�UQt���Ǐ��N��"t���)H���&ZH�%S>�+�G�w��w�T�����\��ߴ+�y<�$D *�s�2l���^9�����"3���>0+�`C"!$��j�����K>t9��s��Bب+S��qH�B�^���c3��ݑ���2S"�#�߳������@�4�c�����?��R��O.�NK�"��jJ�u66���atAAA��*f��� ~c����yÍ�ˇ:U/�?64LQ|�&E`�0:ח�V;�I��deeU�^����)�6��:u�����^�N�PάA�����5��+� 1+]N�f29���ﮃv�����f�E�*R�������uI�@�޳�4��{IЉ��|�)����C�
���6.]��)i#
�K����R\b��J�S#R��O<-H);Kߞ��lqQ�)�4�S6.�etر��"6��_�t^�Y�m��C��ڬ�H ��9�4�R?���
�,�#�?�w�'ɺ��6�oN)���_�>�؁Z���_v�o�Y����c2]Ml�;�G�C-�Σv�m#��gd�W����O�x�����`�7)*7K�x�]|��L�l	�������,�b�LxCP)��>ˑj3����썩���NQ��O����(�S7M��B��;��~W����бj�!�R8ۥY��$�x���N9 G����ɣo���R��,N�5qX�P�����V鵙N>�B����4`˼�O!���SG5�-u�e	�[q��cЯ]���o�y������(�(��}��2������\�rV��jA�������C�����;�;�,Cn����8���ħ7�,��ׯ��?�#ɸ,*])��6M+�=��Wz��:����V2���xgP[Mm(��ε��}�����1,�g7	}!����? C����#��ͱ�$9�����U��C��E��Ԓ�����&����������Ι�����⵻�.��9�0G���&N����[��堗գ����M�������SE]�H�e*k�~ ]qz��r�]�V��gE��NO�����܇---|	))ʨ��63D��{n#$T�866f��u�r�:^���ޣ$����8YV�YVl�|
�,���ۯH$|�:�(�Zw������8<>�Tw��5���C�H��p��q�NGW������h�[�9�^h�ziwޑ/j�r�ұZ��7����=k��j �ޣ��) �kڿ��F�d�~~��J*4�М������*v��=�^|�2ǰ��I��L$p���!�g�О6@֏T�n5�$ǼH٪�ɸ2�(��wdԯ�{����8K,�NuvʎG�;W��'D+�Ͱ��l]�Ұ?�Af#NX8�O��5N�ڕ�l��8�#�������7O�S覀^3��{���O�6m�Y��N-��`F�������G�k�Zr��s`�A��rZ��O�O�tɷ�/F��W.��[[6AlFa�3���q�0|9u+���-Z(����r��6q���Va!��޳�O��m�|a7�4qħ�f����.>�TM�7��mȸW3��(�O���QI.&>^/~5��[��I���!{����I�E����5���QɃ�qog(`��U,	�W��jѻ���+��g�-f�ϓ7�>������n�h'���oO�����䪕��F�xl�*=I����й����0��>�l��6�j7�RAW�"V��
��Bvz��J3jAgBXL7qx��MJɻ%"u8�Ef������b��UI�(�Ɠ/bZ�9@T�.�<�}�����;��q:�,����/�|�!�h�����T��=R���Vٔ��.�m
�������9���O�tA|�����Y��l�2k7����˹�;���j�W��Y���Td�\o�^���t���Sj�[�X����CF��3�Fd�f�/Kș��S��&>g�tw��؝�,4�uꗑ���d:��a�D���| L����;4YE&��l���P������č�����SV�����~]2V�C�r����UaḶ��5ytS�v�3s%L�o.�u�s�HI��}��jЍ_Ihm}nj���Q�X(��Yrن��K }}}���eV��ܯ�u���w�{y�����^�ǻu��������;�m6~ݺ	)�|U�{p۽�Ұ������"�;��^9�}�ȹ�/�E5�(���0�7��M�rN�1<�2��7�t��C��]2\��D�� �4��_�-{w"���ދ�?k�!�����A--��Dk��w��0��9�抇q˩��e7��6��u�n�h�hˁ��0rX&mko[>ߒ0�/iz���/�Pqص��	�n����ffC�f�'' &R,��
����z̴e�q	\;5�F��\���'��;�������R���\���3�Qߔ0f����)�/Gv�5�b�~���1r�+��/�D��X��m�gӨ�!V4.����.�ё���Ϸ��o�t��%N4c�[5�>u鎪��̕�_n�����C3�<k�e[��� '��m���{fJ����r��ŶbjGR�d��۷�ֺ0����9�ž|uqq1�_Ev(k������d���z��gބ��T�����!�����t�|(���;���b�ݣ�����*P+��%#/��Ub�3-z��v
1�Ą��d����8�~�� I��~����fm�������[|ލ= ����w��J����M^���w��Lr_��H�TT�oN��/����5��S��ᆯ��bk����1k�_V�����֨��C����������pǢ���^*Jʕ�����\�TЃ1�5C�ܙF�@��߶m�����54b�[Z�Z�X��_����1,��T�|ߒ�w8�>�����P�5aA��[#�A��OnUV>Aߝ7Қ$��q�L��?
ZfY�S�i���w�1'���N _��<6;� �&��#�Fd J�Wc?����gϚ��K�|�����!@�s�t�v2���.�$�C$�!XJTB�{Q�F�AH\\FW7�@���t��YO��u�9ԑ�g>�bZ�&���H�|Vu{.f��Aw�f!�E�(��L�����{G��e��S^M�W�Z�x�x���6k�7ANDDD9)&��BI�A�m!i��"������YL���ѣ	t�L��7��[׮�4�B[��8?�x�[��c�`����lr�(�����ժ�*�(oR6C5]]��"� ~R!l�4�����2��4��@/��U��M��cp�q��=�K���	{��=�x��А��=3E���m�/�0&Bs��Y-�c���T�z�mv=t�b�\�&��K�d+>w����01V��Fw'#y�DP4��#�������Ы23��L
�q�B�2�F�zNv=���TW��Kȭ�M3p������{�9�/�Ys�'�+*�Eg�����^ZZ"�t)��ڜ0@���o�V��#��n��G��c7�hk��%��N�u���X� �e�>@����0LE��Z����w]ؘ9������|Q�L�18�}U�c�|�ɴ
r�6#lz���LLL�v�zBXƟWكԻm�9bw`_JD�3�I�f��z�-2˴���śuF�,Z���.1�t��7�C�ߔ�y��7"��_t~��֗��wúg�@W�ʤ��R �+�W<6::�>�aT�3�`6Pd��1�:۳����߼��)��>o�ru�O�Ag�&f
"�a��S11�0��8I;�MLL4¿�}s�΢�<Ŕme��,��\c�9��d��Vܼ�E�z�A��iih��Hz0�V�U �ꬁ8�A7+7y0i?d�ܙ���]7kmm��m�����]�Ŷ=�+41�7�ͥ�	*A�)�qv���}ċ�}`��ϟ;s����{d� ;�~�Cv�Q����t�-۰/mi�4�V.+H�U�jȹ������VJN.hƘ}���|���>'�#_{}�o��\�r�EN��^%k�g躼��d��y˙N� e�������x�Be@�Ǐ�H�J�&o����[zO�m"x�le��lD���C|?��>K6�ثvsq!����e�e���f:?�nB�		K��$�`t�kF*4�M��"�h+�#�?��4����F@�0�d|�fuc�G��.�U�(9���t#V��'�>]�ll2 �<�1G�Q�b���_�t�c��1�\v�o/R�����R`*��nT�P��t-'0�kO���� 9��|��ed��o��F�;8VVUјC�(f�����KjT �:����b�	��|cA�EB����vڗ/�YXYu+?\��BS���O�����o�J�Z�l,��L���n�v� �<߿�f�zu����X�&�#$:�0��&�C�y`�Cxh�]{�.�"�썌��Nڌ�Db�k��O�?��!����A�q=��{��3���5��!��q2���4������RQIE=d��uG����1] %M�����qX��=V�������v���5�մ92]����Acv��1Ϡ�n��ppp��*�+�����a�v��,T����Ң`
�=��M&��<~߇�ݙ:ѣ�/!�{�3��$%?��wF ���R��s�+y�L��8�Ç�-&;B=�T���|�>�5�"?�GE;S�ײ�&� �>w�\���Ͼ���ݱ��5c �8{_c�����Wۦ#7-M
m�ە,�be����Ĩ���m���ʇ*��$+:�c��S�j�M�zF�VK��Yn�����pf!Ǯ�	��}�j�l>�Х|�QR�'V�0�������{�2!�}҅������w�8/��$^��	 ��b��3���tz�cJ��������]޽�Y�h�e	�h<}�N����H��3�� ����i98���^�o.�h��Iz._�EC؋S�N(�i�~����w�����J� ��ö�?�������BN�S�)��y�A��{�| Jm�>����B���0�q��c�?F7=h�k���#�T���
V������X��F�ߞlj��;@�r��=������Q_Skk�+����~��emN��|��i�� ��"/�&-mH.�\G<��ȟ?��@[qqq9�"�)��Mg���D�nMRդK�k������H��|��vD{vz�﹖�mY�7�z F�X[��䙚�β��?P/͉��g���!!��=/�R��W%ϕS�g5�����\��W��5=���6.��yz�]�O�����p��33�,
v�t�r2���O7�����)`h��wb�SOOb�|�̳=��~�.�vc������ɛ�,�k��Z�b6>��E�Ƀ�A:��^�b�5�e������w���zv ��7��oM��z#`B�GrP���b����q������.r��Bc��������-8C��B�Py�.?|P޻w�<�Vނ���;,n��4uk�'0	0�7oݪ�n�'!#��b.%���y	w�nA���+�{z2�U�����������_��g]�p!����~��p�4!!�+n�=M�ByԘ���߿��!�S��f�"�6C�.���aQ��?��4�.f���Jy���ge��Y>��z��&�A���8�{��'ǨÛ�K�3�
#�ۇ"�C�V�i�Ȇ3|�����]�~�C��#��Ds���jH�v >�@Ȣ�NbR����ײ����#����y�S;B �o�$i��<|�0�a�K���
#o��f�9�q]�.��֯���r��(���l��y�Z�s9���鎤����nolK8v~ ��u���lq#G<��f�t��=|HJJJ�z�A_MC��� v4��#ᵳ�65]"_b���1羱�a_?Uօ�AjT_��j�Y�'�YS .��Y3���c��%ӫ�]��~h]\CC�����"e}Nl�4<��|���hrz�<i�gV+;�r�0�7�o!b��k���rN�S���˫�:@1J�>��� ��[���Z�����!�9�^ �[uz����ڜ3T�q]+����Jt�e�S,6u/Ş�L�gߔ�����{e�������	�8q��wϱ7B�#�O��J��TTԫ��\9� r���c܂��
�:-S`������:�ۋЊ�>kh�9O���G?�@��y�O���Hv&���E6/�n*O��e���T�����$$	:-qHM�a�KJ��W��&x
�����9a����-&��S����� ��Q ��j������E�����?J�hl�����],�?Ɏu�����`�BS��t!(���4~GW#�kR>��.�.��0@p+>���B��&�$������o/Q�}��\bųdd}�1Ԥ�����2�y2E;�'��u�̫��������ׇ~���߂]n����"nk±��o�����i�~������˫�ys��\�]u�����'�)[[[�a��R�f�^?�]񽲲��?���2� 8�C���_C>q%(L���t�{���{�@rq]�`0�
- j�>�`��;�L�3��G�\�o�#�ᅡr�=�^V�Kѵj��e4�kЕ���Y:��]�;1!A�h�	�4x�6`~��$�t[k��[�n=���a�5����">��@ [lL�e��r�X�-֍��FθFצ{�S!It��3"22�l�
�<���x���������8o����i/@V��5S��6BS���C��8/��������*CT���z�=/��Bۜ��tY�Iכ?��񩈆�N��� ���������ӊ�`��J�(�(�MP���q>|�t]}�ܤXBW7���o?~l��ի)���!/�Ӱ��r2�������Ѓp���v�!�0}�P�En=J��G4�Y���ν���gZ��+(�����Y���B�9�x��H��j�H~No�xI$��}ȓ��	�>��\�����"R22�SI�{>�L���� e��̷�VWW�K=}���-���D$D?�r!�W���Sc��)\R����	����aL^�N�{'�o꽍�v|��T�-&��m�ޑ��!���o-�F�E���0���"��"{[�$4��;��&��j�3����Eb����J+ڗr�@�f�z� ���qT��_�~m����M�_q�Vx�\AFF���E�ǥK��0���������0�2Yk?��q�'h��#=@�Ƥ��6�..�� �����"E�����8&#5r�Q��u`��M����L�q��-�������-S;W��P�l+���f�c�7�����5#�|��q0��@p�{k96���/����@�X/�x��<��1��/_���vA^bտ���#㳿H��=�ʞ*�&椭��+%Ĝ�����k	��/M #�ܞ�|SV^�3000�@}{�3�+�4N����77���}��ԋ�~k�Zգ���˗/3�8������Qw|N?H�����BCA0�9t5zr�ӫ�B��C�M8C��\�v�l���)�G�@����i���j���j~��~���-)��}�vE�[�>��.�Jw~8��i�wH�@o��-����x�Wܰ㔁�!�sș�s�t;�+In3qU,�$�K�8Pl�+ݎ��I�d~+� �g�8�; @�&P��E>� �����X��Zn��3����B�
J���������QQ @�II}��#��{"(�U���R��]�c78.{K>�8.���177wk���認� ����_�%��?l�i��>���\��11?��1�F���"ǵ�-�Y�J-��	�8edA�rJ�NQf?$����7���t9�81=������y�vj�W�<#�ٵ*	10ys��֮�&���;{y��aAhv�潧f�}�h'�\�`.����(�r݌�ׯ��0*�R�>��'�ĵ���n�La���d��Cs��7sB��;��e�ߥ*���y�����U�X�);�~�|���Ғ��Y���c=�:�
��>�[t�qq��`��+z��]tF+?
	g\%�l���{r�=�������u��Ew��}�0w�����]�U�)E�T��6���M�}=Z���#z{C�M�bM�����z#do_�3Z�'��Mƣe���h��]NK**~�d��9��d���Nm|>�O����Z�}�ϋsG*�[$����/�Yf�Tm�!�� $&�6��S9�縿��0�	�+E6���\���4u�,���l-�PN��#����zH ��E^f=�d�MÙ�쪜'�6�:G���ʏV�b��P�g�NA vrȕ"[��������3{���-@��ڄ�_/���Q�n��&>9�,hwq�C�X��G^^&��ꊪ��̌~�\���-F��-�E>*ݓ���ʨ�g�
`cW�?#�zYS���@o�`���{y_���?�(��{�Z[Ay<9����5o؝V��USSSUg5*�c0�k�x`�۾������k�|9v>Þ�n��N��N�ᱼ�<:���+`�� ��p��^��y�N:٬>�+�g��&=�q�~�w�s%$U���\��=F�}���܋��!Ă�V���$�W����8���rj��^��(@����K#���g�\�OmPX�1�\���S�K��F3 �	 ]iJ�
,�ҷǲ���X��a�H�i w�Gj��X��?�q�Nbjjس�ϟ��<�a2��>M��\PP�.�-M] )��x�$�ޯt:� o,?�V������n�^ݓ�1�c֨&<ik�-���6k�->��,:}/��g�br�N��f��SBv��ڭhE�/�R��;��kU�Uu��[9x�<�:�{?��i��t��%��94Ԁ�?��`��WEE�7�w��l�Ll� ���n>�Y�*z]+a��3�ߚ����c!�e��?�7�.Ow�jxP.y_�B�+%�%�ה1Tz��6�g>�o7���%�~ۂ�3������Q{w�|����=��7�6ߣo�XT?��I3�N��_>1h�d��6�~{-N�Je���fՑ��F��gIIkԹ��3���Ï�oMU�2q�E�� A����C�T9��xS�$+�$&&V�vz��%���I����B�ZgT��Xs�	���%�5ҡ:1|�Z�kyd|�M�Z'a|�i�|�d��ǎ�,�����_o���6̲|��d���W�Fo��
'ɤ�������c
&0((AIuM�'�	m�����zteh%!�ya�Pz� �T1�U�P��� 
h6g�p[�0�nפ������ʤ<71I�dw�����3-X��O��.��^�L��*�%O �7��S��Z�TT�8�8]
�&a��d���1l9(��8��c9�@�袓�v�R~��	x=��l�z ��"�c��ɜ���M�k�!W]_�τ��-&��t:a�b����W��l�9� R������i��D�e��.�]ڒ�5���JBLb�W�t8�it�����i/�O�<	O`����SZ�oOS�jɎ�vzõ�.�D1�]���)H�Ʃ�$�W|����@0e�r<6+�?LF��� ��ԝ�t%Ԙl6�c�Gh�akڑOyy��r��~5c�yߕ�OUIE����v�˙W��IC��6M5��j�W���0+<|�f��q�! :̋65�|�9Ş?�S2��C44�1zP*���}�'w�/مl���L4^E�kk_�x�@R�����c_�o4�|�^)�@BZ�
ô����*�ʀ�oIר��N/��+Y1��I���d+�?hq�nFdȚc��X��]_0�zXK*q��&���~���������� 8@`��6���G��1��\JJgw���#��zY�=Й��y�fa��pH��ˮk��~04���qT�t|�!=���>g���`���^֫iiT��u�6�1vu�Q�5����3�F��Q[%R��6~	������/O��] �^��x�+$$��МX�����G�s�"AR`2�O�av�$���]L�/ׅu�(qq\>���W�7�Z��Ł9��>4	ld���#n���ʅ�UUUy;K5`i48�-x�021I=}Z����]Ů�b��䋒��/t�;M^�Qkk�M..������3N�={qө��2J��2��߽��Z�DKv��/rb0�D�TX��/��ho�����]��oI`5������|�3�E��	i�݂��0�r�KKKϟ>�Xn�S	P� yl��Υ���]���:d�9����`�@(C��UZ��c8��u��в��ra��>j�F��U��V?�w���V˅������Қ���޽�]{�ϲ��B�@P�hjv�+`���abZ]/���)��k�Lj�z'!;[����
M6��㨟Z���eO���o0%]�h�a�� ������ˁ��߇Y���&k���01�d��Td���7<�����`jz�sP�u�vm(��|�|�G�M��ƨ9�<ev�I|���ɖ1��3���eee"''�ە.����v�^*)�H�>��y��u���ۊC��y6�{3{8��������æ׿K�z��$&��,ۿc��U߶,��7�@*��{YĄ�F,�bϟ���9��#oa&`H�
��%!��3&��"iL����q�����r-���X�P�B �e(����@�"ۮBW���Ft�m� ;�P����u����
����kq����:��B�:�=#���u9��L9C�%�¸h̽�,]�q�ӧ�n�>��8�Y ���ѯwS-�>�##��n���/��.ށ?�M���t��]@Ω��t��nwƀLF���'Y�C�Fv��c��B�qw5o�^0-x{t/�zo��������]2��0�x(AQg=z���D"'��U�ڈ7o���]�j4P�>���I�3�I��o�
8#Zq���QyO9�]���"ϝ;g���8A���r�N;�A�8l��(6ha����$���L6��(Յ��+��J�߱P`�����zcނ̧��S"�`S�i<�D�?�nF@D��Ny8���nMw�~[����T��:�"P�9:��ϟ���f��GN�݉�復����iK�a@����h(�[=_��  '�`)�32V�w�����)�.n��o��;"�a<���72c"��+���0l�?�M�)C�m�ey��M��W����s��l)R�h���컛?�o¨�r�'��˫L�luU�&�1++���AFL�LO7V���xC8�V a�?YF�h- ���J�x�B�\�jN�^G5�]է�7��1%]������h�ې������D�Ċx�?�}��1.:ҹ��mr���������~xX�Е���D�TeT�洜���se�"�����?��w�N-*RF�6����H�G��T>���0�� J��1�7aJ����j�1@����o��^��+A>
����L2��f]��u��3�"�1T�x@[���F�c�9AdL�5�7��>a���+*~{{
�_WW���f9�����k�lv���,�&J�X�@Z�k]Zq�%w���IT���CK��:# ���IO��U��xbR�����3��˧JpG���[l�8Xc�oG�&9�b��5�1}ή�����>�<�Yz2�I�U��W��'�6t���0���@ ;�2�)7d��m���qbع�Z�nB��j�-�>2����kws	�孪�%����5��������|2'RRR`��vFo�I����zp��o.��~��ll�]�X|ލ{��Qwƛ'��#�)�%@�f�GF��_�4%�%��T	`��k *���k�&��v��?�TAGq?�)\r]�݇�ld�;Ñ�^qT%��\]���r���uoN��� ��{5�����aff�2�	�,��9����=:�c��`F���7�Ο��ucêeQ�BM�se唲���
�5��q1Xz5���eq�(������X�V����;�T6�����[PI)i�ͱ �CS��o���cΐqVzw�~��) �;}��q)V��◢��1���h�X�<AEӡw��Qu\����E�h�S��>�v���{E-*ƨ��L�	�;��N^Ĝ}�`<���>0IУsh-F}�R���ETt���)N��[44�A��[9ur�8'��*	11�TVl`a9�Bњp^�>�:�#����g�0����g0vI���24�g�2D�0ᨵu���y*~�ƥ10~ �a�4��G;��8J\x�O+R�� ��@tc朧�O]��@:ԉ�M�s)Z"c��?�&�! �pqq}c���Z4�abQ5�֭j�'|&SX)�`�1@�>+�ژ�)�=�o������-�������g�+� ����jo+�c���N����$x^ggg`1�k�'j5�)c�[U�ٖ���V� �|}���������|(hT�rŧ���]X0F	o�`"��1ȋ�"S
^^^hi&-WW��X��8��St��8<��NwZ�!B��i���s��(��s[�#����,���򟺖`=�'�3���R>k�s�� .���HFu�56`2�@ZN 0��Ł.���U���L�h�� 1�� 6�����sNE6Q�ϞEA跄��J��{�⅘�#�nH@@p��#_M��i.��2����T62m�p�pG�W,�"��o�k|���!$*������+.���\\t	�κ�~�%	���M<��f26����rˬ/�UKk�$Rp�>�D�k�x
ђ�����ߤF�d8�����p�-������MV�5�bN�-�q�(�yM9������q%����K���-��J�6��*���ƶ������!��$$	nn�Q�t�g��v��l�с�ί����W �ӧO�/J������y�v��lbR�A�4:�K�j�x�A� q�
���^b��;@r��8����!R��0CΓ;N�C������P�����|!�4x������ory��9t6�޽{7��c�������0ڝ���	C�%�����?q�C����m��"�{ ����;
٥�}s-J�F��(AÁ�I[���Z�A)�  2�	{RdLՐq�y�ÕS�On����א��g�^�]��o�?���D�xX��㶂�@�VC���g��-���5t���g�ug�s��tj�|��1�*��)�
t̓�o6'İN ��3֌�r��B���_�0�wqXxKq��ݴ.3��O�]9��|dq����?���w4���Vl��؄̂���^�N��2oֲ�3�R0݅ͮ__��g�.���3Ja))�F������m]�S�q�-�Q?��G���elV&���A����l�:%C��TR� �aԨ&D�n~
Êd@Q���i7^�]�q�K�,��4��˟�� ��w�#;�~����T@>HP&��ER�a�b-*�[JZ����w�cu�顰?]Zro�A+�D#���l�@�V��&�Q�_T5����l�D����?��dE4LZ�~-U
�EL�%u�8ήv����lيs,�^�X��ฝ���1��(ir{j���?]O �o�n��*���`ǀ�p~�E�%xY�:�I������!��WHE�d�H�����+�����Ә0�=����[7�T�N�Κ-j�^M���F��b�z���V��xD��*X� `b3���у�s<������!���0r�&��2��7P^ݜ��ՠ�Ê����R�ʜ�.��N�}�� ��6E���@g�� ��5HK؋��0�X����9�N�Y��RG����i;�z�����X�'	Ө��9����Bt��3� �!!X�6�{4��9�}��t`H���ف�be�U��#oy�:m4<��z4��g��,��į7���vr�/8�`�Ss�מz}:%���B��)Z`��k����ڵGfj�����Eh�����X_�4�A��+�jos|����da>��B�b͸�����4+�Aa��M�nf����jw��kt2<j7��7V�^RC[XXc�gj�®6]�Zf�l���	�f�l�t���ק���K^���C�����՞Z@j���N� �����r���Lj����7�x~��F0�_4����'�Р�<}���G���FI���o�`k}�h[S�c4�(F0�͈��4)@�A�o����Cmq�A�4�S�a��|�.ƶ�v��ƃ�`<�����Rr�����if �[���ؘxЍz3�i���y�I�B��,S�u��wh?��f=�:��*v444�Gm����M���;j��X^M=wvqٺ���ݽy��/��ж�3'2�p }֫����)���1���܀�)���8�~��
����(�>������0�п<���+�Y��M�.T���ؗco!"≚��&��.�-��H�fGߞ��!J�u�i3 ��.�OeUe_c{&��F�wv�)��� �x�ʬ��x�zD��P��_�Iw����`o,��z��uT�E����jPoss3�I�[\3�[׮��c�%/f`kg�!d�[}��5Z���=��
ρZ���ͨ#�5���K��E�?�8�c�U�z)��/��Y�� .��kj�,��tt�U�{0��Ǎ���SiG���R�BN��***� ��w�n,cm���g�1s8m�o=>������dd��hCOp�\�Q|�O���"ݎ����f��Y̕����ޕ�5u-�[��U�Z�,`@AD��,�(hĲ��QE	�@���J�u�TR�%��U��f �[��%�@ț�������{���'ܐ9��9���f�̙�G�j�`���>u���#���˗Q��כt����|
�0B����d��� �{3:z�x����p�`w���B�aFF�m/u��Q�L2�n٩ �ş/T1|��� �!�R?r�05�Bn��F#���0Y�d��g��9��,Y�X���.�T4ڲ��rL۶��eVnIE�������1l�ʓ;}}C����a�v�.hَ�R��p�o��A��;r-�Kzp"^�Ԛ�1��UGk�:��Uj ���U,(��
�P9˩���ASOo
a�/QGk�v����h&���4j���r�.n\=9�ȫ1�u�q�+ 	��D����>0׀.A���W� �Tu?)	e���,/�F��09��
l1��>�����*�m��P��T�EaR��b���'����;����؍�(g.��'ǗO�k��	�5""�.*��	�S2Aɣ�Z � �I�S�Ĭ,ë�7P�.�z�y�X�J�;p�DRǚ�����Tj����%��m���d9�0b`���K������H	�(m{��+���a
"�6�7@�V0p�]w�J:x$�s;�����^;1L��b@���z_0&���=S\�T���`�+��~}i]ޞ`og�����w�yS��?�(��?�������O,��ٓ��\q�ZzNsN$�ơ�n��>��6��lcS@؅�ya��'WU7��;�"��XH��&!!��%h�$(tr!-��ח���b0�R���6��V*h<d�����M���q�el��R8k�����S��ibt,�I����vD[`n˹�7� ��A,�8���x{��`�?��o|d�S,�IիJ��s4i�K�MiPY���u��[���5�̞w������������e=�^A����{���,��\eu�xP�nU\�EFFF8�� �C����i�9�՗_&t�cu�I���B�Oo�XS�_�9��'���!��B��ҭ�we�"Y��U	
<*�R�R����ƺB���OiS))hЩ�F-�}���tk�g�d���~����ǌiow�A"��~LEE�����&��dQϪ��<@8�ɻ{`D����Z�5���Yb.��(�u�nғ	y�P4�Qkk���\Lv^FY�h���g�A��}����n(�i25	�c�Fj ��"�8��"o�@�k�6�ڼ���O��o���N(^��12Ŧ�}1 ��-#k*1
���3�=8Ҟ6�.B1/����L*\��&����?^�R�lHƚ���^G��#%֥�z���>;�V�o�y�ui��$����Q呾2�MA#T�ڧ��Т�k�?���_?~���g�Ș�\�����m�2�;�	��P���K��IjlJ1A�som^�9�5ľ���k����@��Mks�����y Hd�~��4���QzM��K���c�>jn�: 9�<���we%tq����Ͼ��+ 6w�G{x�oJaJU����Nk��D(��Y;��jc���[���I���\jA�X�=j���w�;�|�����t ��;	�4��1�o�U������q)��[\aEY�G7S�-^��<�0l{ɳŅX�V13�C^�<&��w��Uk`�0���~E;�"��F��><�������<~,�s �3Op=����b_V�.5v�f�vRo^[<�itHd�/���*�_�e�h�YE�6Q\�|�^I�R�ֽ��3ؠ�>]�
`.�W}1N�٨��;�4tg�"�1�;�z���e��{����P$V_?GBA;��Դ����=�z��k���*�~�m��e:5�t���O>L��upw*Ʈ�WB�����$4	pm\�լ�^#ŗ��f�)��f���S�(�M.���Ӡ�߉�[Z�r�xG�w���;���3O�i�Y�����K��]��u�w�Y�7�c�#��r�X]v�!����C�w�h� WdS�4���A�-��`T�';:J>�W������m�A%�^|@ި�n�g_����fNY��^�-�xy
ѧ�$��Rmm=�z���� ��Ͻ����T��p�d�&��B�S�W�D�B����0�Ca����0x�SG����О�E[�6P���ѩC������ S�=��`��-X��`_[(���m���
˹\{N�7����4.�[g����/�1D�z��ؙ���9�u,n���m0��������8o ��K:k�7?}�i���2��?Er�V����wT`���B�����62pR�\$;��į�����i4ư��"��A��|��ja3�ܸ�y��,��8�Lv�͍d^��RQ��T&��zL+t�Q5|����o�ս�8!��m���̉���۫������qd3^�=5��;M���o����8�3���ߙ#�x����J�ĩ
��#����]�^򧕵&��n�ΙN�a�z��Y.�rb`آm� aC=>2_�rc�G:��w�"URω��*�I�@J6|@1L��b#��Þ�O��Š��Rf<#���`6��"�ӕԷd�+�$���èQ0V����|ڤB\��V��
f?+p��v����/�8=w�n��"��]��B��!®�d#�`:�+-e��FZ&��`v��6W||����)��@��EVJ5�R����x�ӂ\{Ir�i��ɓ/�G��0�4��7���l���ޗ\���8NNN�n�v��Zo���N|�3g<�N3XWu����γB�cVff�����K�>��ǚ�%����>-�osQN('��	�rB9��PN('��	�rB9�H8X�y�|��6���go�)�����ˣ����w�p�2�љ�����>�7�M���B������?0���C3Ev�u��f���r�@o���A=�$hd���E����������f���]�t�����ak������PK   �<�X=A�'>    /   images/184639ba-f95c-4173-b99b-7b38d7e1948d.png�Y�S�>��hDi�N�;�SJ���>��V�����.�.��FB_�~y��wgvwfw���g���l���.9  ��Bd5�y�Z��gͱ�~�s�� @������ik��y��{h�X{x��[���9�`�V.�6�gb�  �'������خ�qHG|�;p,�~R�f����B��6�=<�8B���b�ŉ��������ʈTl�%=�WF.���R^����N�dppl�c�k����MU'�Lk=p����z8P�]��������
c�XE9"��߻	��1�N���9����u���onS�B��YNK����@uþ��Wl��2�&�V�5��q�T�O�����Ǭ��Ab���W>[��aQ�g;�W��ꎧK�E��cA�.A�	�~�F���o
]�\�(�w�r��7�6����J�UU��My���...'����(��e(��W�]Ե�l���Ht��`��o���{g[��H��;�Aw�w'�C���4�vs4cO�􏯏��k%��A�Ӟ���ӜN��p�z�J/���c��YN~���_<���n��$�?�DѲ��VÈ�����z:e�H�{ÏL�������'�?�(͠��@�z���)��l��j��*�m�뮀C����������l:��~�pѕ~5�����ّ��~v�I��i<fO�a��fZ�a�
���RP�ƴ[�j�����t�ʀqo_r
0�t�)�x�_��k?���f�D��횯Q7o��_���d�������U�F�d�V1g`�hB�+٧J���r�\"��ԇk���Ȧ�"��7�K�="�@�w������|%@�_���[�?�pXK�]MT2��!\3� ����,�r~��|����a4-k��\�=G%��g"°���h�O=��*B��Љ�,�y8�jw�X�c�D�=<-��D��%���jM�|1��|�H����mf���ط岍�-܈?�f�'�I-�F5m�W3yL�/'عh4����K��Q*�Ӱ�P耴�ňZq�S�h]�q�����y���Q�gMnl�H���؞i���4����[Y��6̹O��\@�NRl�VU*Dx$&d��L!WD�w3!�u�\?�*��N�ͽ�T��aѬ��R[/H�(���V!��G��w]����^#����-�F,ol�gkmՉ�0��֖�U����"J1̕Q��J^2q�j��=��z,"D�.g�4�Vx�̣���G�d�t5�T�5X�n�Z�����Vkb|+���U29�a��E�]T8���ӗ�PlO{�g����7�(��P8Iii�LW�&ZH���s�M�U8�Cp�~]o�������u# �{�L1%
a=���eT�k�9��C�Z���=¸�MC������R����
<��[�H-r+�x�",�W�l���?\�aC�X�B�B���]͝��0�pV_ܷ��j%�C�^�X��?���ȟ�̙Τ�m(��il'��0~��Z�(�� �ДKՔ:��$��:0 *R�bd�+�]	?�G���>;#M�<�Y@�{�ۺF�!�&�9.-/;U!(��B�J����9�]wFq�ma:[8F�ƛV��~��
�ר��h�y���*�Ű���ɸ}pt-�m���᪢�#/)a��H�������Ya��2s.�����	��n���)5# TZ�h��Њ�p��UnDѱ"N.���y���{��R)�	�(w�pI��eYX�"�UgYQ��|i�N�����ʫU����DI�@Z��c�Y�u�/�m��<{���g���O1e`iz�\�`��T(����,���a�h�����@��U �auS�U�}ǯo���OV!�����G�yQ<A�\�%��O<�����L��.��L�ᣲ�a�tc���WJ`zX�8~��w�E��W�X��0	��݌H�iQ@\W�@¨�zT�Ūn�2$W� %OjW�����Ls�/�И91�^���7����c���V��u��v�Uz�2Vj��Ξ���r9aP*<SI��;�P�tv�?_��|[����YGHZ$��pH��F}B	�LZ{�-#�o���qp=&yAҸ��z���R����WnA�s�2t���%F(Ja�7�b� ����F�V�R�����
̡�|�D̸ڪZ�ܰBԍ{O�Te�r<�+�h�����J��c��f5C��Y���V���w�oN��|[��8(������1L������Q�83��*�G2�Em�2����Ͻ��WS%��q��ֹ��~��{3^�3R�i��~��,�M�����o6t[�´W���:ݨ���}q� e?]NpD��)j�9;h�L9�Pa��u��d�P��=S�*.��������B:O-�R|��P>Kg���r�c��X�w�����&U�����9�3U�%�%��g���2.��P�W|������ zzs�-X"�O�6��B_��/+��c�]d���-A������q[ �ǥ����J����R۷��+�H	5M	K.yo{V�z;n�Ơt�><J����x���`H��&zz�QU3�!��$�.��g�ү�У�v �c�`�����%ZE�q�R�.;��i2fEH'`W�+�eD�P�����3k���(MDh��D�~�R�B��r5U�&����I	�؄&k#0�*��QWd�n�1Q(���-į���[%�:�`�嵔�]�J��\k���W�^ 0j ׉�%ҷ��n�� ���.�v�rC'i��������Ǻ��9e�R-FY�����r��$�l���d��SF������.̏!����Z��7X�U�����H�GePoN����)Q�O���e�1��L��I�D>�G�#c�2;-�N�5}��P Ԥ�F��뇣ۣ.�����2�4$�+5,nf��4��]p�U�=V0�O�y(�����"px��ח�y�/[�J�՟�"sY�$?������AX�)H_&�;ig*e�ڋ�%&��d%\=[�$��,p�"g�s��h�)k�$�C���r�/��!Q�~�1�$��v:V{�oZ����x�b�'�>ںZ���g(8��g�Z�\�9�m7E��>�V(��D�1`���l�`m�i��id�@�k�n,V�$������Z(+Sp����0�����È��@H Zs��n��k;�6�����Qc�����u�>�i���u�ϳ�6	%���F���}a���`����'�ܐܹ�袀A��,/�ǎ�e�������n�^k1��� ���\��S��֊����[���P}� �9�\�+�$ɨ?��ݖ��9�OvR���P�P0Nh���2��{=ld��1'^|��L?��Mj�N��.�)�&,�9x�+�# ~�б��r��eJ5��~ [�#{BYS�k�r��Hω������V��P�Pa~^݉���z�篪�L�U}����C�_t{���Auvz]~�Dª��c��c�ټ�6�7G�7,���m�A7E_��; �;=�D<p�mWm|ː�S^N�OJ�ˋD�Gr}�+}��ql�h�.W�-�`�ǖηչȖÞ.\eD����jZt�"{0�GA�w����4d���w�\�pD��n�mc(�^!������?����T���35նn�[�}���>�ՍeaL����,��|$ž�(��22T����К��&���Jc�	Ҳ�uT�b��0���� ��:��65&�	(�D�|��:�<H������!����kƝ�7i4* ֶ ��E+)�_�*����T�DJ[�k#85$�RD�|i��O����^<��&��{YgҞƘt�9��T�&j��f�7���(�0mV�6�.�GD�'���T!����
7frPZ{���d��1��Mq�lϡT�6Q9'FO���=4�"� �u�e�¾g�R>�T�2���X��n��5��"F�sf�h��?IW�ȷ)�L�>�z��Y��F霂��zC��N[�O��oG-Z0J`ak�Y:���{�Ў��f�&��q��m&.��Ǆ��e���j��#�I��$�/�!��X_�ﴆ1�� g0b��"�V�����RR�F�o�R��{��#-E*LH��5��"��S/�ŀ~�
�L�D~�lrQ�4����	�j��§#��,����-��h/Y�WZ��NB��i�O+��FB,@-�/�u5O1�7.Z�:"t7@�Kz�ONº)��F훡-`����΅�����G� Dg�.�,!fHW�&S��EqPB�֘��)��9�y嫆ͅg���Ao[��'|%���;ʰf@"Kx�HG�O-ƣ]��6����1I����HR�ETj�y-��$!����W��cuh|��Xp�}xn�_�������M}���*=��jX��L�%��s7Y�*��:?=|�6�qW�h�4��9	
��p�J��0lmC����q�0,i�lɾ?�w��Q{.��&K��&/���־�O�ӊ�z>�}�s\u�0&�㔢7g�w��`�ȸ����݌f$l�E<Lew����/�ց��M���k3�9�K�υ��,Z�����ʈ�g�c�@~�^�D��B��V_WPQ��Pe�I|�k��R� �/�RD��<s܈T���J���ʷ[�)���y�eǕP�X��Eݕ�6�V�unC4��ș���k�p@R/iq���ȣ�i'��q/��vp�H�kyڏY�][Fu�j<L�8
���eQ��c�*��CK�N��uy� ꙴ�G2��������9�liF�
��E��E���˔2�q #���"W���TX�ک�+9��n����
 ���>S5�s�j�S�K�Ff�q`U�>C'z�6�9:>��W�L�m�8�1�:����]��l�F�T�7�g^����h�KE"��U����CȊ'W�~W���l�ă��F�i2��PVpİ\�� ���]��'�FϋI�7��v�v)f�IQ F
�n�{ރ�� ���(��3��)̹�v�ľ��a߸�����?ǓŞl9��b "3=�^��}t��ۗ�����^I����5�)k��E���[���%��~"!0�������*�fP��*)s�*M���\�rr���|�(dn8|��p�mɒ�/2A�r,샢�kR�i�?7��/�4vd��%�w�yR���`��S. q�	�+��)�5�/����.�B�cC���f\���QТFɽɱ�����/���r�yzA9��h��1+|.��v��j� ��j�+��;�0S�TRQ�e��>���r�G8,��=�����0$���6���n�'�L�6@�X��Y)K�8��C�۹��ba��B���h��m:�C�H�9�q�,���K#I���(�0�wru�kA|�~��|�H�ȋ/��_�i�a�<�QG�R�'*d�r��l���s4�x���9X�;�M1������Y���F�\y���֦#�܃_��fg�p$`���,`ӧD�����(m�F5���]A)h`���X�r~�2��[ʈ_8]Ѿ��ya�TwO.91·��.��r�pf�V�Hvm�G[#[�O�x�v\�b� �pt4|z`^w¤��u���?<��G+/'�CȚ��r�hLoZ��;�(xK��e�>)��n�b�������D�Q7�
	������Kf�3O]ض�[kh-
�5ޝ.�@tC�P�m5W����M��|W)q����R�ƸU�����Z?�vg��R^;�?��P�-���I�+'700b��^�-x�MrQ�Ȋ18�%)�^�5D�c�H�S@���]:�����Z���1�8��W�dQ�R+iή��QU*��,s���0��WRN�P!dzײ[PG�i��U1mvI���9�8)Ɍ�w�j~����66���s�	q7��}
�����K�E�5��j)fC'$�c�y�TC�h�|�g�u/��}i�����.7�3��u����1���/N�ܕ
~*��ԛ����:��-<�!Z�Ab$ ]��vU{`�}��t��<v5�2�`�{�8����|]H��o��\r�➮^
��B�|�.z��3C��RY4��� ����$���+e�����Ri��wV�i@�.�x[{�@�C,�1��H�X_=[TE��6��8^���۶�8����,ˆ{���>~�R����~���0�"���VO�2
�a�??J<mm��t>f�@32��uS�+�@�t��q�2��ux�osލm��q��2|�����X�Z�����5%�"
ߧ3p����d}�b]��n�%4�1	�A����C]�㵚�b�0��Vv_����!=, �xyX��h��`��6�&O��NHj<����?���D�u����溴c�>oM�t.���x z����t��<��Sk��c��;J���O]gʛ�ڞ@��'''��E^��b� :!�4�D�L;?��M���g��-W����I:H�ׄ�����9�Y]m;T��s���s��N�Lח��o��׽����~�}��n_���t���2r���b��As��luI��M�s�������Л��_��m�w%7Ø僯DJ$"���)��.5s�]7,<ܪ_�o>,4s�_��[�
Ӱ�x���4�x�^*��\�}�1���5�tTYE�z{DjW�x�M�aa��'�  (x�a'��ĺ]�P����_�n�L��:2���4��S^���l{z�-�Wn���Mx��H���r�Ϡ����qmCɍ��fԦ���px�ud������ʣX�4+�ti�#��9��ڷ���k �|�%�3u���k���GܵG̋=L��(+	��H̪�_����rS�����q��Q4r���x~�Qz�1�W�z"{��:^� �O�r��U�f��PK   [��Xw�'<�  �  /   images/192efd05-ebbf-4f69-b47f-23f46b924e86.png�YeTг�%�nda	�E��kI��^b%��K�������.i�F:������9g�3�a��7w��U��qipQPP�d4�I�?����w�U��8.
n((H��0�o��?%5\V��l��p�F����9ٻYY�Xs9��f�Ҡ��~T�����:21�B����l�1*�(WH���bZQ#�,Q�Q���C��T��DA������I��׃q�t�}��1X���PRj$�km@���1qd�j9r��YG��]�~�Y���WX�z=[��5ҵ�� �G�2Ǧ&��PI�c ��p2���*t���7F���3�7!���X �R�Q�n���aI�2v�̩���A����99��}�w�ܦ;9�l>`�E��8�������Yz��a��O��W�q��O����:3(a�{4
�u��Wᵋ&̪���F<{�j��kr���[���mUY��KR�x�P?�%�^T�H�m�^����?�`�D���Fm��H�w�⡂s��&L��B;�Ґ��oԒc�MR\���������![����Mb�'�o^u��O0��'� LP7���9X{^�=��c��m�(SL�clv=���п�-o�I���QRּXI�)��A2�v�����?�jj��G"�Z�\.gۻ�)F}{��J��� RΥ��b�zL(�;1.��>	���Y����^��cD>�A"��f����Sz]w�m��a����8cAeE�ʽ��8�+0��Q�
A��*2�<Q�b0Rz8�$5�9ˣ�U����t��/a���F�$���>��ăU��VD��aa�}>	v��
E��幫������m%���iW�:��	o=�{m��ڜ��X�z��T(�^�xPG1�36WA�h^����aqly���RY�?�����Q�1�LFv/(]��|=��jg��X��\V#s1π��ļ�*�D�]v�o:��K�<h�^�Ә��nO�[��
�X���Ɏ4pc�8K�S�p�[���*�>�;$	j#C�0�'�,I��3gIi��F�U�E�k]wS/c]p�ܜn�:P��8�cn�0�_�ު�T�1�Sa���)ۻG8�,:�e�PQ�ƛ�Pd�:q����B����U{`u�g�`�Oq>29�h�6����%��9�4HO���7�(�_%)#U'b�GY�O�:�9�W�ܥ�7��,�]	��S
�2l��|��z���]���^��^��Xß3����f>�(M�r�|�5�K�&`�|�v���Vz�Ԫ�^m�y^�
��U;�&�����&�U�S�'jϧd��=�ڔřQEh�%�Zfp*q�TTg�`͂��K.]��ǭQ����1���䦭|��&�Y�o�HĈ2�$�ѽ�嘅*�<MJI89���9�ֿˏ�X��͗5�������Q���Pl����}Fn����Y�w����雅&�|*�V��ee\������#`K�7���di�/@�H�ᶗc����� �2f�qp vug��>�V��u$�*H����Қɕ�����n]��5��*�Lb@*~�Q�Ah� V��9`�j{��
��@N<4���p��*0�r�y�J۰�1� �Ef�pZ�4d�f�5�L��F/�V�@�z�.�SLeC1a�H�ڍ�B�������~���ݠ|A�� L�Tx'l*��GG�]�!�3}��+Ղ�[����<�s�<w��4�-F���"w�J�\\�!����Js��x�;�t��e����O^�皈����w�f�d��/8β	{ύ�IXh<Aͧ]�"��[՘��Y��n�?�c��ގ'�����$Q���k�u��J'z�5����'\�/��}M��[!����@��my�w�v,�d8��t���zrH!J��/�8�9ɯ�smdN��<وD�a+E��x�0���8f�����c_����n:c}��4�``b�z�
���b�D�P���L���@j�R��k��q-�O[:?�)��+�MD)����tG�X㾕�D�]��2ڟ�*)�Z�dxy۾���(v4==�,���o[�T���QbE`TfD1�Lfm�p��8��/{;��Ze�u�s4~���ī�������uO��cno��o�OX˙,p"�m~��496lNRU-��go�`�[�G�j��3�az�|1��6 1����t��M�+���s���Sh��5�?O�~'�v!L�n�p|�c���@��ޠԟ�g��P��7�aY��]��"�P���[f_���7H�\'�2�y������pM��d�v��NKѾ���<��$��6E��#�|o�t�7������v�?�N�򕋑)������(��̑�{�K��V������1bM~$�ل�*A+6=�͑u���6@gN�ԑ!��g�"����Nh��b�4��r�5#P�>���g�4�ӛ�q�ַ/B�z�a`o�6<J��*�mt��"6����N���ö_��|q��/g�1��M��l���5f�n�Vs14X�,,�l��F·����S��})�v������Ppy�X�:�N�E����%��&/�i�l�����؝>�~��{�=W]㉞a;2S�1x�G�y�M��|���U6�-�H���]��ơ4<+v4�ae�1e'Z8�Ύ����~ȿ�3M6&��t���$k��
K{tg�X�l��o�!Fd��Ż$	6丌iho��7�����cO�P����J %炏�{ 6��Z����dSk�W�qO|�:U�̇�	�߹N:g<�JO�g�e߁�{��Jݦ��UBD�'������T�������䆘,aI*է���^��Cn�<� Oj��;Қ���bU���/����WE�t�M[aam�����޴QY�v�ɧ��8|~�L��6kI�&�|��݄��ز
�[����4�l�۸��9/o���Q&�ox,bOK!:�ՔzX<c��IB`	����Ѧk�q�����N�|�Ƕ�]|����4�����jx�=���G�݇��_ϐHU'���j|��Sdot>n��Zg7Wl�룳@��n��`.wR�vA�gwRs�m���
�E���~��2UDMjH�2:x�Cӵ����*�9���E����dɐC�S�K,66d�!�1���Xp�qS�#��8����1!^�,�̞�)��+�0GX�`Do��[�w�k���*�Ŀ�v�����o��*��7�R�-���v��gj��e��#Q!~��?yxW����}�����&��֪����CA�U�%O��F���-�E��a���K��Ծi�q�uS�f���G�h>�*�1i���
C��L��&����zz��O�+�/�]}p��m<<�XfRX��'j)QL�3��	������:^tű�q�*�PQ�I�0^B��l"pp@P���,��-Y�죷$�7+���Î���a��SЉ�vb\7���a�#f�.N���e�G��L]��$7��Z�m���2���Y����Xf��^��2�hT���(��O�)�%ԊL��W>,
��&��dm�{�ew�>��� ��e������ǅ�m�qF����{f:���l2�$�vf"kb�C�`&;`%�����"��:��c
by��C��g�����´<�]��~2�o{ ]�/�(u��<*��~ �e5��D��6�ng��}�~�p�D� ��+Z��N�f�>b�F(qGg*շ���s�$n��5/�������Z� ����҉�ٜ¥2���1�E�����pW��,��ߠ���n���[�p�Mx>��f���xd���$P�a�q��Y��{�#���M����oi@LnU�U�b)��՘��_lm��q00tX�z��JU�6��[c8��\r�U}{�y6�awp�P�Q9���eCe�F
xD K&Q�'}!TϦg�����2��o������ٚT�u�G��ő��/"�2�5�F�e2�,Ww4b��e��k-K��7,�BM-s5�/�&d�Kͧ7�\��c���ù��v
�޺�iI�.��Z3��E-'���_����'ٔU���*�� 3�{��!�
��w�L��X��
Ņ�!8xO>]�ԛ@��_o�=<0���%������P�ph�H[��]k�9�:'X��r��l(N�J�l���AQ�Jd�qjQ���YT	�M>��>V'Ts?ܫ�\T�s�H�Ǻ��"vʛ) ibF,�1}�NR ��c�}I�L�C�Z�P��P�MR-?=�qP ʕM��*P�����}5��TG'�9�J��ᐒ��ˢq}V��6܇蓜�C�aT&5��2��Ut���-�#�8�m�؛�)
�|zMP^ݤ�;�+���ZI}�������)�u�,�3{��{uE���6^���p����d'�	n�X�e�~Y�GT�b4y���y��4�@D�e�6b��%����r[hH��7�����4J�67�D� �;���� 
�G�xBm��z�o����8�vp�s^���U�"���!}�%KL��c)d��YЄ�����6�.?G9|��0� ���f���ޜ���u)��ڤ��G,U�:n�T��@4Ck�.��b��#��D
��EA�s�s%(��B6G�s��o�x$�!�!�*eO)Y��N�٧`⛉(>��W�F ��A����M��G�f�+�J��ƥl)~~�g��J2C	vh�n�?0���Y�Z�㢾r��?�5]Ei)�0`1{����u3��O�xF;|xE3��a�w�t�7)!"�R��`x[P�^�]������"2�v��Vd�"���=����i���'<��MQ�Lh�11��Hb8fc�3D�j�,UM��1$�f #�t��1��>��P��|�oZp�����|����Z��@&����\^����j����F��a�+N��aq��%jm�Pt���p,��@���)�)�ʳ��戟6���I�s[s"�E�t=쁮7�{��X_����1������O��I#���k�W!�^���
#�j�c&�Qq�I�ʳP}��C3e~�dZ��E���}LH��	�΃��O`�j��*�MA�߿��"�r�I�CzS�~Y6M�
�7�J����n�*�Y""�3�L��K;�V�(����M{+����)Z�%�Jy�ȣ����T�M��{�ai3�Ǵ"今K�^@����V��(�����/�-@�5���5�a���CD&#�'Zkn��Ԓ�jf�z(�E���o�wH��=�RJ^��������V�9�h�7^Znt7�"/����F�6�o)WlH�*���Vx�3���%>l�W_�@Y��$8N���e�Sw21E52��g]/v�	hy����c$�9{�r-4�7���[zw��:7��7/�c��,e=9L���Eyx���{��ũY�H|h/�
��0]f�(��|�PX;�����zU���w�%�}<IZ��d��0�;�me�z� ��/��̈�2,�n�3����ǟ�ا��:}�E��a��1��*���������,*���cĦ�ȋ�ʩ3������S�T_�l�p=*�UjY�J<SI���p��yZ�5�����W{|�\	✡�o��i����>6�����a�W{��UB�H�C�i�� 0�Eg҆�rԼtf�h�V3	���P ��?����0�D�#V%��0����~@���R���ՠ��b�v����w-|���Y�l�D�@i;� �C�;W�T��c-��H�&Aެ���6[�f*��}�Tj�7/K�S��~������yI@�<�^*�y3���8ա�^�r�\s�w�z�I���&��T2�ۓ����7�����2��`�=^�X�&a'�^��𼓻S�p��/�n��v���ˠT��H�qi��#�l�ŝ��ܰ8��X.gr]i\����E�~��z|���	����l}
N�	����Ki����V���u�hV���^�wv�	����~sCM���
cb.�����"���(����n�ޢ2Ck��l0��5��Bt*n-I��CFR��9�i`���C���,f@��'�C�̲= ��į1�$���Aπ�(�y`��OJdD�q���zO�b�Ot���,��=�-��EO�޹1��qa)�򞑧�)w���ٍI1O�d�##����rcǑy�u$�6����)퍭:F�5��и�|�=��8�դ�^�~�К�!%�IZ�$ �ز�W���52��sm��fx�#.MKw<�ǓwT66����0E\�k2w�r�$%{�p�B|������b�>9��i�nI��j]�K�}0ߍU���[�yTήzM=�y='�� `�ӕI	u`�r*�[�R�I����ߟ|)@Eirx��4 �я39¡ۻ6�.((2�;Ȣ�3kO_~��i�:��e��u<��u��b1���+��V�$�hUh�gB%�B��ߙ��ǧ�6�}4$Y�9j{1*��m��c�@���&��,��u˱K(tqbV(�6��������Υ|���]r��[Wtaq��Z�d��ی� ��9�U��N��,����uy��-���ȸ�����E@5_?b��A��'��eun����}��;� M%�9��k���z�:�h+�̟�w+�-��t]vh��UN}�X�f��P����Xn��UZ�M/�F��fn���9G8Y��PЋK�]�G�oւ~�8;e,�=�>�Y-����3�l�/Q��Y��I0K�mL8�ķ��W�{��^��L�A��&���u��k�:V�k�@	s��2�-�hm�rO�Zܺ�q1�=��`�HkL������=�D￫�#nk��f�7?�ͤ�|���/��6Z ��g�y�1
�ތ���J�_����u���Υe�T�Q|x~�ՙvm���})����H������qڑ,(r��Y�Q�R�>�lrϋ`Sg�}��Z���+���o���ׯ9B��V��2;|=�|���m����0��7��V��d~��]�)��V�˥�0��/4�e�BF�� 3o���C�~��'&�����������=Oѹ�_���<�h�xh9w���A/ٿ�ޚȟ��7�)���ş��G}P(qt-���uB9#�-3i"V_c�"�S�V��%�C�)�����J�V쀵Þ�Є2�If��Qt��]Hn|0��e��r�c��#���5I�L�����Tn�)[�o��]Ჲ��f�X��)b�3q��T�#~��[�*T~�1���=n)7R������ë->�R3>5��(�*S%m�?PK   �<�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   �<�Xv��� f~ /   images/4d249bba-3190-4770-b321-fb8fc027a237.pngl�	XS��=��-��P��(We�@�U���2)a�)2�\�N�'"��@9P0̓��0V� �� B � ��oZ�����<}�޳�~ǵֻω׎�Yl�z��[1��9HH�TKHl	�,�䧙�g�|�+��f�O�f�����ly:TBB�9�練�'�*�9��F8�-A t��C=�{���f��A�ۡ����辱Â����{N���N������-Ү�7�g���װ��6���������7!AAQ�}�C�����w4����K_��������R�{�����j1���}{k�<��=1�VF^x�/8o��P�p�[L,��^Fi���0UX�����W�C�ʰ�e9�N��'�"�1����J3�����B���Y���@�ڌ6Fն|/e���YMFb���7Q��yp2&�(�0�6��j����Հ���_ڟF�Ǡ�����c�t��ZD<$����}��p=�bu�l1|�m�)L�N�Z�ش=�Qm_}* �5�)�6�dK�.�
�}s[\�g���L�
Gwj��Yb�>�T�n"X����m�Er�$	F6��fw�oV�`r�������AU��b9��X��E;Y�{��x�nް�m��C�qF��p�8ƽWW��^�tO{���1����?
�1�*b�~��wң�(VN�[���i{������ ��91��\�-~�sA8�O
���R�x��BL�ġGgº���j�� <��qx�V�{沴1��tfo��qҀ�aHW��@p��H��׳����*x�
&Έ��X2����]��;_�O6���P�Z��D_;j�g�9f�몫�fQ�̩��22s��ܾ`_�?���0H;�Y�\�ЮB� W�?G<�-
�ѫ�С'�$K�<�lɠ'�����D^��@�P>�p��9۸�妡��(�n�O^hb�^�a��:�*��GA�0~���A�̨��r/����
� ��T���R�>�z�
��2��7G�jL(�PL-y���J�#ݖ0|6\�ѝɒL
��/�=����FZT�GA�`���[�8-���P����B(���0��+:���%��<XǞ��F��ʤ֜�����t+�&<у�R��(l8r�9��~�[���@r��2�4Qs[������^J�+��s�
P�L�|�H�$t����Gl�5wZ���v�]7�௠�2����'��|n��K�NcB�������œ�=�O��7x��̹v	]�+��6�ryS���i(f�=a!Yx��b�;�퀖3Qk:�����m
c��AV��/gG�,��WQ�e��^
(��WupA,��}F�o��5�()�75�t��r�U�eo<I<�s7/��a؍;:�-�J��c&��>��:� �H�ys��q�5�oO��Q�E�1�h��h��~���p���/Lg48'�����yb��J���;�70�����Є�8�)��G"w�\���*��á�|<�1��Oq���5N�7��3N�	M�	�x��wJA�I�AS�_{�ǰX�4f"&-�nӒ��Wh7q�>�\,�z?�Ҍ���:�
���M({,\���-��\���ip������R+np�4ބ��������
��(�Tj	O�D��0���.FAÖ!X| ��(|�cA/x¸�bt(7��$v�'@���d� IܑUYZ�<E�F׬|�5~_�j��l�$��p��l L2�$��M���U�#܇�Z l;O�aV�\�e�p��8v�*.�-ʜO�%�t	��bA�3M��s7A=�	*e�&*�d��c��P�s�4��w � ZJ���2p�$v��ʵ/�'��QP�N���y�r�S�$��6�(�{��)�Ѣ|�1 ��"ju�౓؆�)��q��	��!�fd<>�B,�#5{�'��}S�;��d���B�x��~*���۲4�*��%�ݟ��0puEb-�����}����,!Ḡ���3jA�X@�{��9ǰkA��_u���C���Uv������8����^b��`���Z[{{NFN�����fR��M��A"
<p��O�̬Q���@7g�C����L*/���g�Ν;o���<�x���ӧޣ������fM�7�.w��$��x�p�G���e�\i�T��=��-��L����Km��*���'��m��t��Nc-�O���0V"���&����������Wd�nl����j/�~�����Y 02�s��]*����E?�'CY:ї�)�//'�������K*舃��mɮu3팆�t9��\R1Qy�nv󐁢�*p{�>���=J:��a�o�S�ʽ(���#0.� �-�����F��赶�֯i\L��h6���Nt*�*#3��H��ȵ���>F]PLla��a���㞞}u�#M��ȸ������ᄞ�R5^���[<���ZҴ�Uߕ{wt��dge��v;��� �ȋ�/5�LO���I���ynO@{?�.�,�A~6u0G|�a��P�=q��P9h
ix�~��|/uf�Jls����p�%���XGz�ٯ�8��Og��C�ePG�*ãQ/8��z���0�C��>��7��6Ӏ�97>��&���%�j(q�A`L��<	k��L1]`�����}=�R g}yᖸ��J�=��� i�A�탢��^#{ל�-h@��)7�2�K��W�^e�K�ڔC;�@Q��	ۤ��1����+�NJ�ݎ�yL\>Azس�Z5��k��@z�H� d�,.x=���Q^iS!�F���ȕ����4Ǌ��:xB8�Y��&�&��Zԍ�۲I-)櫋�����<6��
�6�i��W܍��yF��/�N�^TF������=�i��t��|`F�$˟Z�Sf@��t�XY>	*n(lچ�Z*,��C�k`�=�E"L��{6[����S��
B[�~e�*�w���`O�6=�8t�!Sq�����^}������fO��"�I���ΈuHޟͱ�Ep�mS:�#��d�F}|h
��V��o�/�SOF����8���$>���Q���l��N��3#f)'��rCe�9�Q-��s馧`���)&ô㜾�tHE37����wS[�&*�cJm�x�MY��}�cl��7�E�����b�A"]�.��^!��f��d�d�����Qը�2nz{e���-��w�`�s$z�%���E>�qP�w��y����d����`V^�Y�D���œ����˙i����| 7�yy�"h�H0��_
���숙����r�C. X�誀3��$�6Ͼ����R�i�ho�c��m��ZsKQj��I�4T\�$Pv�ހJ�C�r�jζ%��7p�C�<���.�㥧H���f ��AT"��`~�ސ�O�,��Pw����[��6��ͣ�
��(GnW9b�����T_���}�=�������b�� ���ct��2jؒ�����U�cDW�pC����$���c�A�[���ױh7���ⁿ���|k��4�&܄�@y�,��s�*w~�_(+�X�1x��$	~��=�u��aXL���F��;��j��&�I;�oj��ωf�D����\�3U#h��S�s7ܗ?���Eb���(5DaIf;��}opn<D~����D��F�`���s��s.�*M�ܺ�BG_�
aۺBx*nP��ǰ�4kv!z��u@,�(k� 9�/���)�#_�..m����2;w�;�L�uT�?�VL%�<O� �jv�"�J���r�kS��-��X,��a��s��%���s�Gnl�f�]�,�K	R���#� Y��bV#8������ќM�"�L�C)�YX��c��lT[�/(~0�L-�4�96�VP��-Ud�7Rf�9d`��߽@	��+z�_?:�;Mq�� f5DO��$�=b�v��ſ�P��KVA7F�����~��T���2N��~�0PE�F�O�췢6L����<�nw�Vr�S�&W�ϑ���^Pa�Ą�sR�������jf���j�<�p��(�'�4�Q��zZ�c�̿X��F��7[q�U�~@t����w����$r���=�S�=`�. �2���i;W�7N�wD]q�����Tz0
����O�0S6U�KQ��j�KjQ �LP�17�|p#��L�ɏ�@=�����?Pѹ^�� ��b�޻/8�0<uS:E�;Nw%�.�u ��椝�w��3���MI�X��h�L��t�)���i1s]m����F �C��oq�F�9�qh}J&�s`�-P�N��Yw��'��YOM��y�/F��� ?n�KŨ��=[����*-�?M3�+^Jb��$�i�����M��u;��~xJ�`'�o����������a�3���2��R?���������#6'1�"<|�:�%F�`���	�h	Z;VmxC���#rbR��O���4O�3@́֜f)�?O�vm%��Ew�#�����ϑlQ��9�J�&^n�_~����G��$�%���R�N=����H�6.M�Vt�������|������}�#�4%������XC���@���P�뢒�AMӏ�2��<݋sv�⡬�:�f���%߬�� ��*��b�r�N8���7/{��I�8W��r"�3�xܱ���ίw.wH�|��G�m:f�LH1���F�.��]�3�0:�!>ÏZ�ʽ��J*�~8�=�ο�rB�G�}�1��%��uci�v$z���|���ypq$q-t��V�O�րB�v�9���Y�:��>�VyJ�W173[�ĆG�g��YԺ��S�a�
=f�ik�M^��'�\f,�ԟd�Z��	5=ͱ/I���b��8�|:�.(���(��v�E����\��XҶ��ҝA���Q�d�j�D�:2�x�Ǉ/�ƻ���e@�L\�t'�=R��eN?��LX��͉l_f��_��]+δ\��W�Ye�Y�C�-(,4��7-�2u��5Fż��}�%w	e~���# Nt��6.�������NS��wM��:4=K�z�2C�5�Q�_�4��>hl��\\�M� |�2�����U���㙺 	��3�qC����j+Wz��W��F�B�@k�qCC��|��?zX��y�_<l��8X+X���u;���!	��|/�~�ƶmۈ��[C�����)[�ϊ�z���̹��8���KՊ�@5��Q[^8
�\baVH���XQ�a`X��PE�����t��ZrD߇W7̣�ˁ����&2� ��������sZ��.���v����TaHQӈ���,��$�J �zМ�P �ߢ�[�}o�io߾dh������y�����ϰk����N=��a�29J���*�ts l8�(���q����!0;��E�ʁ�ؙʡ����	�I����b���â�~���/E����ViY~
ls��r+�q�ن��  AT��u�"g{m�&�L�?C���H�{��6���j��:���FtB�ٙ��D�|#�fw )�Qmz��8��afp�0&�Gʫ�h�	��ʋ��)�JY��Ճ�΋����[���k���i�����֤�*Fk@�gmA��{0?
�z�� y���K׈���0Ú��68�v���61�C�c~��c*�'�n��y�FK�ݼu+�2��e(��u��3F�nTcO{(P�{��G7gh_��Ϟ�p�O�8z�Dό�	홹]�q��b+#�aڻ�(���k�_
���R*��.���G��~�〴�(��܈����^G(S�n��M%�젩i��˗/��}O���-t_�vm�SO1�>3�عx�"�?�o�4t���u�D�Ak9�KpT46���,�UY��[dj�����kY�mО���TS:s� �Z?9��oP�1r�5���;�ewLw	<l�� ��6�(�x��L�����$aإp�So^N��5Pw��7�Q�������:bL?���D���vgݻw�����o������)� �5#�/�F��|,͍��2
�~�c��d�;�/�w��0E>'Y*͡�i�d��? �k�N�
'���+dj�9�ɽ§��w��a:�@X�j�+U׵��z�
Lz|Y�B^�'4l�eS��M9�l @�@��וz���^l����>�Q��o��B�`w�b���b��2�[2zf���^�L&�\�{����[��d�����aܳ��/��>���쵈�5�S���d_�:�鄧��;:Db�^K���])C� �~_;\���k~
��X��BOZ)���ĜB�6��whWMۖs73�|�Z[�^ ��lfH�L���;��H���tJ�gV~��dV<���~��0�%>�WL���kV��FIw���FO�+�\4��M�{gMF#��cfӑ�S�2���7�^ݺ�@�����"2�Q�'��ǆ[q~�}Ip.�'!��\�<�n
�W(9]1n����&�z#��PB��y_� w����Y�^\S{��}��B��u���=	�̜�{e�cP?��z�k]��B��g3���2�5I��L�\�w
��I�m��|b�Se�Sm�~���O.lB&4ۼ3�sW��B)؂~y}�^�S&�b�΂�RW�;��|�ra]��i��r�k@�OQ`���"�;�I��&�4H���ʔ�_?�]{�L�1gϞ=S��i�����5�)�E��c&��dcgɵư���84J��N���f���Z�+A!��n�|˼#��n��O�<��}TS���YY1�g�.�V� 1� ���N}��D��5J:8�;� F�b,�-**JW}�N�OjQ�]�p#���x3���j$�A�ry��L�������ٗ%�- �f����F�c?+���M���n��:�U�L�	�B,��fJ	Uڌ\/	2����u��bX<�^<��8$�I�:��n�n<n��%֏C�:a��	�O}��%��G.{4zrL����C(��>_x�+��\�%��I���;n|�{\���~v '�Pz��{��޺�۸؊3=����8w�.'XrQ��p&<Յ%W�o/�c<G̢�_5ǂG���+�yV<��C'��[�f��{������h����*U���o�F��`���ͼ򷙼D,V�ň��d9���^�B
͝ȼ&�_�w��	�\/�F,�	�g-�0��}�di #��>�WRW�3��irdw�H��#+�H��/��N܀��R ��b��(�VG�V	I�y�z�{l��K�G�5d�ʟ�_�3��Y����Co�c�zz��o��Qڈ1$x��u#�C�>����t�4�5_�������526!�=HƯY@k�6����';��)�b�,L�il�VwZE��[O�3��g�7v=}�tkϧI
�<n����~G���΀/@[���d��1�ӈ�|�.S�9bs�`qp��O��Z?H��\/���I+ŀ��>��FI�3� ���`���1ڒ�z���`�.ؠR�UC�й��.�+�@�'����	�>��.v#ԸSV�<�q� ���S����uz��X�{��v]O��f�Z���=����%���*��Щ������������e���}��X�O���f \��+U�:WNw�������в��v7�im1��r�CAq���d�ۘ<ώ<{2Ԩ!�w�ͅe��f��ؤ��/�d�K,y��9u�=��hl��G�t�W��|��fϝ��`�k�`�0��A�l=�+v�}�6����'�JmJ��+U��I�q5	r��E΋�z4�*\[w�'}'��m�o��U;.���:i��$����{��'��w@%��q�{1�s�oL,�Q��s~#�s=�� ����}et�Z�Zw��J�?eKa�2���pGlC�}!Y��$��t!�G���a	�))�������\��~~S�7SRxv��wPj��]�V�{/��`�-�o]����H䅶�]	���DZ�f�;E�h�����:>�&����8: �I�c�%��0��0:%C�7��c��Ka�Z�0qY�/y�8b5Q���j~��Z�h'��!7�%��M,�2�簈��������S�]�ČRC"�6NHt�:�Gzr��y���rA���
�C�A�ȈD���,4u�����e��w[�Cw�م	,��}�b�����`rr2S:�����@�;Wp��#r�l��O3Ж�cF��ݔ�x �����֔V�0/cv
뉬[�=K�ӟ��rҨ)�nXM1]kt�燌Mٱ�P|/������j8p��&茺�D�w���6�(�4�9 �f�#�k5��.
���^����j͈8�f�����B��K�̓�=�v�\z�R+���I���v�7��a��-$�^S�b�*}����>�&�E׳2��%�62ed3�0�i�51��i�Ob]�c}?�<���䥘�>���}f�	�}^n�B�n��o@'H��Dq.�������`x^T��@�?���yϦ�E�vj��q/�܋W��Bb=� ��FǞ;�r/��gg
�'��.~I����k?P��LdVN�eB��`��6�R���K�mb�f.	�h_p<ΜȌ�I�p�eJbZ��$���Pkf�0P�K�"�l��n>xY����^��Vi��l���6.f|��Uf�]遗���n����/��͋���0���r���Ϋ�1,�d��{�5�����+��[H�����		)'��/��a����r+C����ġv�"�������}�0���-�)�lKfhU�� ���r�j����	�]�W#!CD��a��ń�l��D*�J�=T������=&P������U��ow��H!�)O��Q�Xm���|o��� $VQ��ޠ��b�Z����/:u�C�!���[�4��^��	��:�mE���7�H=��/���E}3�J.3���;�Y"�^�R(��7����zP����j9G�&'�r�
.5�~��
�������{ٲ1�L'��[ųQ�V0��a�(�0썝�F�ڇ8pT=�/zC�"7�N[���Q��755]���
��{�]�F�ͻbK��۱�0�
���NK%�����IO}mo$��.���R�k���|��LO�����5l�0Z*
����wPN���%n�����g�=e�tP�;�οv��mz�j>�a��bx���W��®�@h��o�&�۱k��SX0��b0Ă�L������������e�5>�7m���d�ơ���>�34Z�Ʉ�r�fҿ��f!&|�Գ�~NNNW �N���0r���<l_����'���b���!Z"�����b#@l6C�OF\�*	�#�c��P���٣��p��K�M�a����]���]�1&6�X��)�-�v�X�6��r��g�]���Q�|:v�>c�'�}5���(w[��-CB�@"�̖[� J��D��j�%�6�kn���a<�/v~�r�ޚ����U8ه� 2I�.Ҿ}�����m �9�b�D<�:/k��/�EwL�!P�|+���A�sJ`)�� �te��);t�frՔ{���xjZ���shttt8�r��xr�v\g����<^�ܰAv�> ��n���7� ��o
��H��mL�ڶ��N�30�����aml�3���u�]��(H���&ƀfkx#���.�Ef����i �Bw�@�?R& �;6�V�<�����%x�����<�M�L���1��w��;�JXn�uA���g���K��Oa;�,��~%��#V͆k	�h��}�\�c:�j`XgJ��D��_�tu����%ڋ+2��ȉ���*�Z@>��Ø��2�h-���1�g 5��_'�jFt����̣	j�<�w�չ��T[�_>����:`��w�~�u����@⯵�;B���FW�8dn����1U���R�/��En���
m*�w]�r���հOnq���?r
����x]���Sߝ���yݬ�nS}j�r\�J�͙��;�C�Y��e$��!��8�$O yݼ	L�F�;����x�ꗒ��z���~��*������+7{x��s�0�?�+���b�<ɭ���2�=T`�F���C?YB��5�¡=�V���Z3���E��׈���&��҇]�j��z���0��R�
YulX�J��!0�H�z��i�O�g������{*m�ּ�M@˟���bʟ|�W�cV`.V|1gOݒ�%�(����3�B�7�U$�C��w����5�Pi�u��
��B;�5i����M�L]ҙ���������������u�@�s���ߤ�@1f�y�����5~�:�'}�탕��F2�KS2?5�$�oO����9C1e���̎�L�����f���O�;��g>3��jD���*:$HQ�yp�;	�IK���5VJ� ��{[��r��_P��d�͘�:���'��d___�4����19(�C�Ńhʩ	�^P1�>/��P���;$y?����1��yq=QԊ�[��=;�lb]��������N��%(��LA�E��Q�J�c�}�i�\+�3��Ä�z��
G�����au�O͒Rl��q[x9�6u��ӽܡ2�Y��]��OR��-]B�5�\��X��7jrU�8<2�hz�BGqv�+Є�{�k�z�\�2��5�ĲC��Y�:g3Me��v��2�,���Ĺ����Kw����H�var�x�!_�7־�Q;^ߏ�-z=�k�L���D�**U�����VZe��<z}d���xzK������cv���MgY���d���\�J�}|N�����~��}w�cφB0co1�	�Y����2cv�Y���K�M��tp������j���I*�n�!!!�D��kmGH�%<�E5�f*���m@���:l��zs{�y����K��0�ѷ	Ԃ�('�'|�+)<����g��Oz��5��e�j嵅�k�2U��� �_Ǳ*v
����^#f��H����hN��PC�#ƍȤ�X���@��vIp�$��u��ܧy]9		�"s�ZO,&7�RM&B��<w�OM�e�L���m��-C��4,��1��&\�k��]7$�g|T5~y���N�n�8妀�����Ж8��o~�dovv�­��㴋�K;p4���n[^F��%�:�=��H���yM�8����YZ�ڊ�˗�߲P���yyO*+%��)�Js�%��]��6_o�|����MOn��L�����t�ȁ�EQ�x��{�c���E'��'IJ����-�ٍc���5T!�=I�:�5��}�"E�밼�����~���u'�I���C8Qjvy%'�M�5�}%��|�z(�?ȫ1��p�mb��$�}D�$o���]�����Ę�q,�m*�Fŉ
���cIj9��s�j��Ir*��֛$�b���0!O�Q���G"Ӄk�6�4���<Q:�3�$`&;�I�4��7�ԥ<��#������)@��?yr;QZ^�oT�1���T�CY	9�,�"4q���Q�ר��SQ��??���*'�p��;�	b���SQ�}
�V���{�n����Z�[@�^���֋�,*:��=���/\��.�f=IM�J��{�>sÆ�qP��E^�J�[8���#���O#������D�Yq�p��~��q�6I8���ar!�SǪ�'qo�x�l&a��0d�xJ]��cy�jl,9�HA⺈dyW��r�ti`R�h7����������wČi�e�t�f�&�t@ZN��k�4�Xہ�1�H݁���X.�\u�RÚ��]�ݛ�bs�&��ƀ}�*��͏)QIޫ���i�Y
��O����V����@�&�A��9���4�c]d	߈M�$8���fh´D�-�5n��hK"�d0����>\O��m��Xl툺,�2]I�/�7���IB�%B=�z �$�p��0R�NI�+Կ��bh�i�ǇIR�h	���Ƚ�L5�ɫ"��Z��|^kf(�l���	������8��.ryq�/2��?���p�&�w�9� �R��`����.��*{��Y5�/XM�_��C�*��$����$�覠���  x���#f?YiI�Tkex��;�,�b����zJ�)�>�M��I�=�^c�C�hb#�ʂm"-1"k���G��ʊȫ��q��'~u.����ƍ7����]A�զ !$>�J�l����0�t��O�����~���Y��r�@>���Rjm����G�~mmm]-	o1l��E���."W���8c�MC�p�ed�w�o&6i�$O���o8<�m�!V�m��w���Ν��/$�?	NB�Zci�.ߣ�Y�r��J)QH�8Uň�#�A�5��|�z( %=�����r��N\mxKU,�y�=���v8I���V��R�'Rq�x��|�؈kp���4N׎�m��}#"�S%%<0���߲��Q������8��\!����h�V��m�6�#ݦI!~WK�WD���Mݴ��*��ȳHOs�$ʛ�3(���d�K�?L���Y����H؏�d%kV���>Í��>���|��7�I�B��űv���B6~��|[��q`&�*��6ܼu���\�	�9���<K)!�=�gy�v�&{�3g~D�撤t�q�7 ��G���~�&��NR� �%��.�b�A�&��ִ�m��`���C�Y&��:Aʈh���n{3`a fՖ���4rn����'&�>�i�"dnǥ:�;��v�Kޝ�'O>1P������{i�S����d��[�閍9���������̝�+T_Ϩ(װ�&*=-��=4"�!�T�2�:�T��$�aN�����٢G`#����<$��L�.��G�lB��-�]�T���*	��[;��!��W
��2:�pO��HC��!��p|�K�7NVEJi�����u�W��B?��FZ�D��L/���Px&D"Eo)vq3j@,7RU&�>�ΫKsa�yi��m���2?�a�Y�۞n�/�ޡ���f�ǩS�΄=w''']�^�;h!)��h�MF���_<~xc�u��ŻFQ�?~�tɑ�4�\Z�s�j8�.i��(�]��b�j1��*�Ӗ�-�b˦�>˛�Ns(�$��˽;�?C�5�R����Pd�(�겟�͗?�������o�$Y3׍���~g""=S�*�y@]z�c���Iv'X�onnn�Zk����dz��545�%$~��h��!�t��w&�<��u�Z�C����r�����]i��8��� �|���U���O�v,	)ֵ�]Mv����W�\A����ݮ��<�U5 �!�N�c�Iᶢ2��'��	�c�y,��wi��oh�N��#H��Y�� ��V�oDF����V���Z�y�Yic�����V9��D�ѣ��
v?���;�x}^���J>��6�|	���QU"���Y��?ۡ�Q��S���\���G�m? s*=��d)�;�w"��ݢ�Dcp�Ν�tL�3����T���#v����D�0���0o�-� G�����'~�V���x�('2[�qFF��pcC8p<+YW�e�];�|z�����b�赞�

��؁99&؄�܀���/���bAK̐5���[5��e2H�R�Ϟ�)44t�ə�>��k�= kk-ށ@�aR�e�h;v��g۪�o>|�P+�;X!����	�u-H�濔L+�*QhN}� �OL�c���X�ہ�T��{'�!��
Ę�a�0�#.��sU��:����2D"q2�.#+������*]�o��/B+#�dx<��g��OU��xO=�YN͌�E����	��

A���5�F��S�Q��������,*�����ۀD�>G��L�Sw�J?'yL��|\\\ijH,�A�&���"�~���v=�
��X^��b���O�\2���*��@���8JLL9#?J-ph��՘y	m���[մ�ZS��e����L YH|��cPx�!;Ā5��`̈́����>Fm~���\F��G7�� .j� ֓S��$!��� �����}��6�_5�EOe�`�pV��,�ʖ���i֘ �i�JI�9::�/*���֭���6�DG���w�h�� g�u�	Y��x���Ԑ�B~b�XzN|ej�Jr��{[GL��cW؋$5��cv�i��zN(LnI�sL��@��hP� d�WC�|���@�)��PU�[tOxS��,//�h��օ[�� 㝀,�_�u���.�c^�^π���J, �\�����+=}}��PUU7@����{�V�W�
��lSz��|�x��U7H��Ջ#����tedd�#h��(���Pl(���b ������R.�Ҩ �gQ:J@~�
�q���5+��R�zzּ��`T�?��Qw6�(�?=Kw�LN�`@�(۫I����Y�D�l�����BUj�/B@b#����u��s���UTz�.���S���T��>��}ܭ�����R�n`���Χ;�{�]|_J��8P��NV��������s�� ?��th7[�֜}��*P��?S����'�o�����ۋ����Q̪%�Z�J���d��'���0��֣��¨�{�|�pVN��= 3���p%p�,��?�G�c��~���y����������{  ��������Hi����b��X�@E�p�r�wՁ4O����������A����>y�ys|ǡ�WQX����� �Z�bd JK��B����kV��o�w�n�\���u-{��˸k%Ф::bڲ����_=G�����B3w_��+@�;#nݺ�`������y~��[���C�r�a��$�`���~mo5����C�� rZoo�9K����c��z�:r?77�Nk,�6X������W�Ԕ��G����$om��+A��y	�q�8�E ��a[.c��}�!�>H����D0�u��볏�vQ�0��ͯ���h�g�B�Ɠ�0�����v� ��SK�L�Y�G#�w���#diJ_��2��� P�`=V���Z7��E�oL�*!5A�s��X�/\k�G,i�K�R������	D�i4��Pz^eô,UI�U����@(E��a��)�[)���O� a�`-�B�>�-�T�B~R4��"y9	�f�)���i�	�O-9��W_9A��k-MM��8�Є���%�P�2 �ҽ�u�z��o3��VA9��1U [O]��f��E��ٛ�@��F4G;� U�yz����DϐG=�p��s�As�u�Z��*y@�21q�4�,���~>[:,A�jڥ����7/Zo�읉�73c�����k����E {r�$�h�VCړ��I�U�V�vj�kf`U�F�	�x��ъT�c�lA�1�n�3�o߾�I\Ɲ|?	`rz�8绮X�,��h"V�Ov�Ծ�-� �a���e�agg��Pe�֫t���u��9?�$���}�NG���Y@7
8��~��d���u=O�w������Oh��)v��I�?@�;W={13VG/q�*E����W('M>ɡ=@������g���u�"��;�5ѝ=P�����70f�����Ѫ���)�j�Wfǭ��/��I��-j-2Lu�L0��]�* ���	ľ�Ӄ�݀%ש�m�%(hh�*+��H7��k�ĭ�1�4/[V�!纈 ���6vv���X�?�a�Q��n�$�l@�t�իW)�5�;���n�-�!cO�� ����%	M�NB��z��m)��R��C�.���!��D��{)A�g£J� k?�������])�)���Ǖl�g��
���ů�aD�
2U��i���6�b��߮��҈�H�]�R��8Vڡ̬,���.0���7T�t���N҉��Df�H�����r����B�'�����';>������ۈ���xfcqq4�I���,P陃Ue�P`��%�cJP۵�%!R�O�4��H��ȀsF�t�Ò$k����K��~?��\�w���\%;:�C��}����2T�3��*v񈼭h9?�v8�k���sp}���~�uua;6zz�$h����M�%�{$N�DO��R�Lq��Z�v���i6S?B�lY{~��ǜ�ˏ]�x���WS��!�?��c ���G�0�1G�S_���p]�)�8V��O@�lml�� �\/�u(�~۰��o���
M���͸�Z���ΚY��YY
�������7ե����}����?���g�����|�F~*Oc�Z￀�.�,P�����EYr)VB��moVI;fm4�j��g���@��q����s_��'�˷�⦥�.0+.Z��}q ���F�(��2m�S�	���̈\ǃ���2��P�4/�;J]��A�#N5��fv��yg��?�Y+�(5��v�o>���@��m��x��-,�R�'�������{�� �DjZ۹ҫ-Ye2�dߏ�gdK����="d�x��I�u�,϶@����߲f9�_�ˡݽR��e��T��Kx"`��T��g>]����{�A�O�UkhxO�g�KOj��[f*&4M���4����NX!�QPX�<��PL)5�S�OjJ�y ��HNIq�f�#�EE� ����J�����6��r��y�왯o	U6�V�4,�z/�t@O!�P�0�PP�� ��=��F50�,�ݨm�\�%����B�	jCnQ��S;7nQ�>���|��������Pf�o����I�]��ѕi�(z��'f��i|���	�A�w�Ø��&����%b��^ ���j�ZBh��!��,��

@υ#��-�E��^�(�(CrRg��"�&�A�~���Ю���O�g�qu��m
 1l�E#o~D#)�Z&�{?�h��af�� c���r\�"� �7IVA�$+-�Ut �xy�^G���C�`�o�k���eW"�1?uP����w�T����ű�� ����|�f���*CD��]�a�/7��;�h��T@]*�;o|�o��s������#������k(}dI��`��052���c�%F�I(�ۓ�Q�k�$`�ÿdkV�6��m&$~�*dl�+wD�W�+�k�4U�������/. l><}�7�����Dy�#������)�й~��\�vє���"��h���pav���"�� ��k��^G @�`���~([3�<6����9�뮃��S9����Y��O�7B��t1U��N@��5�k�B�<(�`'  ���X�W'�]m=*��R�^�X)�f��5"��  �4��G1��ф���z��oP4��QZ��By'�Ҭr�l50�X�׀Ð����ue=q�"c�Ƃ����/�o���-WT����Iȟ?UiD�j�9�2�
J�r�@���4��������"��P�'ĮO���~��a��Q�
�1!����0���zP8h��(�a~�ڠ���=��D�O���\m���h+��.$��|��b�.v���В�SG6q���D��+��j�Y�����G���e� J�n�?�̆k^�z��)�j"�	�{�\��#U�5vQ��K�_ׯ��)��0O�Mg�Me�0�`�)7��d��{n�D�3�'aK@o�q�=*���̊Љ�0�b�!0��vG���w8D�����k�������&�^c�o:G����ˣy�90��Y���x�-�����	��=���̭��2�Z���*��[�5�/A�T�_o�=����^ ���O�G�W<sZ��o$����ǯ5U3!k�_4[��:9�(>�?ȍ攫^
��O����p�F ���fh�+��������W���^����k~��Ly$�n�\s` �@�=0��s��,�GGyG�)��mC�* �V�"�qB�Z��m���w��a1q0A�:�˨�uؖ��3�4 �/hU������ �r����8-��l�J!22^�4(Y�d+�M�^�SVHB�5*+��{UV��[F�����_�����r]]�㹟�����>���s�l⋞;\c,�ӛ}d���9��B�г�+f˃�r$�X���lV�~�����Q?YQ,�cҰ;ТQ*���R�Bv��/�yyy�'Q��0�m��O��.� �ߠ�j[�����~����1��T�*B�ё���Rav+	27���O���0�z�Y5S�}�1�L;^�3ˆ�)�B� w;���QU\�[Ā�\7��_��2����ō�T�O%� ��#��o3��ބ��ɾ���_� ��y�8�����a����DTV$E�Ë������О�I���nc������9]���F��%���9y����&��f�+�av{��������c̫�vW��t	9�E��'�~<�u�vt��x�<0D�����?�N���9�Q{)^�~��P|S���]>`$�I�ɹ�B��VQo���	���{1�/�k��3:::�/���}�����I l����j^-��`�4128�˟���`�k���@��bڹt]�O�����ׯ_�S�V5���	�CCC�	u;4QUIde��������d���zy
���p8�d�Y8El��
t��leuu3�}	���&obb"%%U\T$6]|�/**j��ډ2J����]W���~�)m�{K����p�J���Vښ��W�J�2w5���Z��Bwإ.Mܖ�i��O
��������VW�l���v�I�17][�n@F�2++��H<���N~d�]��K���c�q&>������:�iu����}��FI���eJ(��&U�k	wn�dV���x�1��n�U9%��T���c�(p/%Gd�(���	;�����wmy��e�L탛�h5��Tt^�re�⩍Ӗ7Y-��˖�l:�^���jְ�`ee%��2	�U]�y"��5{��u��J��ˑ�\���
循�*�P@J�ǥJ$b7!�?���?u>N���2<���L��sG�:�`ĺ�����E����p��)t�,e�X�H�2Z�R�T��|Te��TG����ġ��n���O��4�@a��C��P�Q�!��3�C1m�JDSS�H��*a�FZЫ��g�K�[s��4�F�RŴ勺��7�z���/�G��kH222z�4������kLyQ��(]�گ?-��KY��(���yTq���P��4o}���
�W���KPWv{�wKB9��3<�֩��|W
!q������@��}SS��
���!�f���69g�w�MHꡃ�����-,D������>ׄj6�����.�rN�y�Ǥm�>�:αa���go:a^T��A2����}�D�c
�q�����1q����C��)�Й��r%w�x�>��&�
� ykuyzE7m�@��=T��@�op����Ẩ��������9Q�}q
����l8g�t��o��$��l�����Ə�\3�&r'���ofȝ[Ӂ����𗖕���g%��,�ro�����T����'��JK�tʶ��b/�TPP`������P�p�x��d��hB��V��-;�*��uĸ���F>[�ƍ�s��z����J�?���r��>f�������7�A�nB��]����3P�������m~�
�K�ӗެ��`g�����oE�-�]���>o�\�7@Q���޹��41z���YT�Pq[|�+���w�Q˳1=Q����D���X����J\JN���W�ޮ|��,gD�?��(�ɲ��Nc�zո*dqn��X�N�h����ڧ!�Q��w����CօG??=@��S��%��>���-C�%Y��9Q�+|}L�Vm�x�8&��(la��D���q>�}��5��FȖ	��GM��}%�5����b���;����i=@��M\��Tmc#��t��ř4�^^����"U� pa���k{컬fq�&Ϋ�+=��8RL7+,�IF�{466R10�LLL4�%��(�L~���rW�4��0�+�nß��c�]��g�
��sW;,B��E�iM�}�:M��
h��}0����^�:��Ǐ�UVS{θ�T��)��w�������?J]��̉����e�D���l��ᆠ����iJJ�m�~��b�U͔��x��տ �N1^
�̲���`y�*ȡ*<���I�pZ؈���r/�����j;8���mA�ϕ���o����*���A�-�����qw��(Agno���x��VE���O����(��R1�u�gƣ���!�F�X�t���V� "�g*8ʼi�vNL'v� 5V˱����x��x7hG�x������@�eϠϹjjo_�/v���|�tj�:�����C�E1�`�^���(\7�}BJ�p�XS�������������o�/��0�2���������s555|���&f��V6pbҘ�w�v� ��@�vo	������?{�l+����E����ܐ;�'E0�y�/���{��#C�����7x�;���+�
(�H(�lg�%Х�S��u2
�d�����a�1.L)�w��j�%�U��M+q맷���WVVD�#�ܻ��|8(����A� ��N/���+R ��w�ې�n�&^��ݦϛoa~a���Ԇґtt�=<<�&&P�|����[ $ 2�^V��Q�at>�Q��N<H,�G��sssrr����/�;{�w��|��5vwo8O�h"���gA��~ӈ��^@e�`Q �/S/��UN�s��%�39 �nBn��J���;��:��)���3ww3C����8�9T͸��K��M�:�Z�ߚ��`t�]i�Hd`F-��]�cQWW7]k������x�J�����&Hy\$�=C�4����@��;T���ۑm�\P��`�kbW���7�7�4�x�.2��"	ג�=���S�����H鞞�����n��L��5�U`�a���d��m�S��o3�5��S��-#?�~�
�500��� (;�D�UM�/utv��O�� �FA��s뼽�t�ҡ�C�ng`` �Ծv�����M����Ɔ/���$)���O��]��k��nr��3��Ҋ��֒�Q��bW�p��5Y�^Y$��T�p�
y�n���;w�ܷ� �%�e��xҞl���:���E2F�w��qt����{�yB+	�ʊw[��/�?��,�0f�|E�3%�#� P�gϞ����E��1�3���|�ŉ�աx5������@�>���Z�#����u���wܤp�*ou"7�{�M��4���M�AJ��������Oʄ�л��#$��\y
-�z�����������W���վ����	��,���_
��I��ʁۥB���셬�^R��ɐ������Qo��8���1�nX�؍щ��͛�?�K�����:��W�Ǆ���nN����b6y%�5889����[�w�Đ�>zmbd4^}��Y
T�/_8ED� (N�%$$�#=}�4�r4pt,�ﴶ$�I29��n3�V%a[�E\��&���V��>Q�X�ӽ��`ue4a�;T�g���C� �_`�`�(j�Ns�Z��v$��&rbk���ٌ����' ,,-K��"'M�~+����{'����jd��ݏj�Y6�?�l���[��x"oh-���Aac��I  3��[0���C(�}�����|轠�`�S�Ay����2e�<~�]��{��FGW�RV!'�A�����!;�=�%�jW:k��8\ы�Y�񣚔@�@t�c���+�"�&b#�v9��pjh��f�o��^�w�$��������|cWX�5�Hl��9.�&���v����E�8߬+W���e��D�B�t�����!��3����}�gΏ�#��O�s��j$ߖ��o�D�-�\�	���ZX_OJM=|���w<Ӹ���o�=((�7XK��0��Jo��@�U8��P�;�#��ZD�u\�?��>�{l��Ī*^��6hN,���GM�+immMX�����7H(�HK�O������2������ �c/o����v{��������.M�Ak��5�xM����,���[�i��ɫ�iQhPVn�E�$Pr�M]�(p��p\�h��QPQ�L�6�iRS{��T�+))�a���8Y$�k,�\�ZK�g������;�*�Ht�qT��W7G���U�G��0�3E��^+P�����ؽ.d�YYT���(��w�MQ�F���*���������{���A9G�jNh(����zH���q��@�'�$�6�+��/v�" P�Zѕ��
�}�ɯ��<4�}����*��E�,ⴚv@�JJ� 
G��T�B���'�AA}3���G�s�E?i�uˊ,?pX��E:]�t8_t
�n�3�*��@Џ�͋&)l�V(���
12�"{�H]8��)�76�J��"!l��U4Bw8�y�t�#;�|PfGZ��-�z���E��"�DD6b(����A�8&�re4nn�)cV�@�Iw��H\L�pL���*�qd	H$��sS��6>�d�e"�	�)�e���!���P����8�@��
ٽh��~���P����%I����*��RQ�����E��Ӽ�Ꮤ&O���J�� �!:�Ō�t���%%�A0���l�G����ܔ��`�#,�et[����Kɓ��D������n��I$" Q��Ĩ蚛s;M{i��Y(�76��҂�C;�nP���Z��J9[�g�ys��$�&x�ʑ��E�C��gݗ�A=Z���7�)��co����8���84}���aI[�,��/�W-<V��^��n�y�51��΢���qT�/*�q�p�>e��ԕi�)4]|��&�^d}��b'V�f�-_VVW�PNM�fCk����n�)))�E�>����{���D��<y>�{J�o��8L��������Z�a��d������Y��#�[a�{�w�WƖ��^�D=��dٽ���g�pa}cjj�_]}�&֘746��Lc7N�sv����$����5�܅���W[O��R�T�KS?�+���&;on�;,=�^Yi�U��o��		��/��-�.W$�IQi��*�Rhu,U=J~�:�q�[CY�*]BSSs�c����ӭsK.�����V���7@�A=��rC2�"�C�j�А.�����c���Uv���*�!]�Ųq�iѫke�?A��[&����������θ�*�)��E�$����@���*�����Բ�΀c��u��$�i�D�Бz�jΊof���C�8��ބ&ˤ�x�Y�gXXX� �A2_���`��`�k�~����겎5dP�ۺX����w� w �Q}z3͕�&��z��2(\ˁ����o�$A�K8;;��a���N>�Q<?ڌ�F�ҿ81! `i�7���q#`+o�����.���'�Ք|�Z/ҸT���z˨H�_TTT �_�:YȈ� Y�񶎎�qqqw55}��;��:<�?��F��xd��c���a�N�-���5:hk3���}��sQkmm��\D�{�=�Up6�[������Q*0O��Yr-���KI �����g.����|�!�vzF::̀��p����Dc`�&7��z�L��@~�ZKq�� �������Z&� ������o@�K%��zO��v�D5v�(����g����ϓ��"�jI&V�k>XEM��>
��ؘ!T3-���B����o���`A��=D~-� ٙ`� ��s�� ����^�`QI���h៬�A�B2@\z}q#���At�8'��v[��I���w��J�f��,Lv3:::��0v6���x������E���6���$b��(р��ST�̈́�I����;�P]966Vܙk����P�.B+�u�Q�y�)�\���ML116.���s�x�8��6K��l%__%_�s��,iDԷ3)YY�H9w��]_?�Yo���W�Lj���)4�Q��%hC3��6.�H��b�� �M=�� �z�9As��+�m��jl��@nף�H���r38��6w,��G+��>��&5$��t���=n�_:Θ	P��F��>
�x�΋?��4解�a�"��螁ktt�[�:��X7T[>􂔨��v�JH�e�{�ZP2��V��*C�c��i�хJf�E8 J�M&����ʥ�/�} Pk�����ZZZ'��V�Gwm.h��%ݔ�i��@����P�������u��Q(�4o�#���Crj�?�4!����R�[����N�"�� �v�B�Eڊ�L��l�9(��Pȣ���\\����&0h<,!�r�l
�MT��8�7���ɀ��ז��W�ve\`W��4�{z}�z///�)��Ɖ!��h�A�"�9�epx�/�`�ʊ��Qa=@՟��}�~[�\�E�� !턷�W]N�`"tyk\h
ncf٘u��2����ũCp2��`�C$c�R�jp��8�%:��t��o	�a�]#�����.��������h���{hӾ�����xS10TU�?�Zp��Y�c��Y�r�X(f�[oq&(����x/AL+q���}��࡙��J��?,���M� LH	`r"	
R�č��5vo�v�ҙ34��08E������i�pь��_4.y���W�����1E>�*�Ϗ��OG0UVU�zqPm=MĶ����:	#4]__�мB.ٗ�l����0RH�Dq}kK� �! ��e�Ƽ-�����7tn2Q㍨�H�t!+��S(�FH��K�� a�U˷ۡ��{�dS�������a�� �����C�K({|ᆝZ�Я�$�ddd$�Ő���@�+q24>0�����|Ң�vU�����1-e*�F�{���A���&��B�8C�{Od��y�6�A�$k�ՕN� �w�����<6qS�=;�5�p�����������#�T
�ךlik�w�������#��d3���e������0b̾��@ƠG	=t�٧O���ǥq�S�	������� ��*��:r�9��kME�<8�
��	 p'(�!(nh�gv8u��~����V^��&B��^�s�NG��~�kJB���]�r����G��i�j&��;���w����L�����_r�(䏉���j�!�P텄j�¸qqK�O��6��g�F=��������넥]A0�`4��]:�t�x��IgǺA���z�����o�{�#�/pp�!$F��Y:%���V��dcamSu�� � Ը3��C"N3ҥ�����J�7G_A��U,�W�p�Ҁ�� h�t�G��j�M 2(!4V�{�=U�z%8Eꌻ����6�
k*�i���̸��ͣH�C�HZ�&g��K_b���l�TUU5]]'<����ߗg�
�����g�3e��=|SX�t.o:��32(�f��nQ=7T����		%��f�E�6���iP�}NK��yP�W���3�m��r�"h(���Ω�O������?A�CT�,?1\7@�q�	c1(W0x���cʢ���b���áw� "��٥Y��\��V�C(m� ����\�=zb��q��Q�/��ǃ�Dϳ���r�|qC�A��<�5�,�	x����?~t�E~l�GJ{�1���2��lmQ�r{��q�K
f&���@#֓];�最R<]Ũ2�oCn`H��yl�N<���E>V�V���ٞi#C�u�z��j/abbf�=Q-�0������lcG���6P0T����l]II�Ɔ��iW�	?����c��W�[A�11
:��=h~A@ݗഠ���]�yn���_���6����'̡b"x72�G8I�y��iq48]�����4:z�o���;�Z::�v��/,�]:��T�����ι��a���&m�3���J����9��.Bq�t@���|e�W�J���}"��<#>!6�;�AGb�1 *�ˑPgF��@y�:xSD�
��-yQ��`8��/#��h��lg�/o�Q`K��"�r����֮.(R�x:1�Ah 9Z���q>Q�B�m��> ]q��t�v<�������t���ߒ��M?Y����� V�����Bd�\Aq�GNJZ:�
q�!e�	Cؗ� �)(���^dm��z�s9}�yb�|��볝�vTN�w8�|�����'�R��d?�v��yL��(;�h0������
�1�r;Q�VG��V5���e�����`�F�2@6�����#uޔ��#P�28l �L&�\�v�]6GX7���:+?	�9�!>��I������QU`u�Hcvv6��{���Qȃ�Wv�3U�;��%���颭%������+�����UWG��	�6�o�����)�d/Zлv�?C�=��;bw����������X?uxS���+�|�SC�"�R��^\II	hN���{@�Q|a�؅A�I�����j�F������L=�S����}���L���1)���jW�.O�Hc|rZ�+lTz���ϲ�s���L)��V��b��:�m���2[dX=�%?�I�M���^j(�����kK7�5�9����][�1�G@��M�j��I���d�����.���Z�ۂ��:�U�:+++���$+�����7��B�=D��� j��\_T��qW�c��V��O����p��`1�b �a�I��^0�=��ȢP��[Ղ�&L�I0�5%^ǵ��7�~��%�!1An3R���`��vA	h'4�@�L��A�|PSOrC8�^��h��07���iu��`�`ܑ�LxAgҗѷ��J�`���ҁ��oϚe��"��E��%Z<z;�Su��<�0߷����9
&�m�=�S{Uh04(xW{W�-�k�U���v�CGS���E��~zn=˰w� Q�w}*��Q�������
��eTO"](X��@�`N���?��bN؞Y<��.3���٢w~t�q��7]����)�Y�h��l8_t�A��N�?[L����ڂɦ����K\�a �-���g�@�CR�[/|�1TC�3��bAae����ˊP;::�y �T��,�qu�&Y/���n�uyC�7V'c ���-^X ���ń�`�f��`3���3S�E$�X��j�c�z����e�j�۷"�T)�i���L�aN+�H���$���E��z�4�ʦ��9����mF���G��`!S�f�����Q܎��_���=di�}V"�P|��B����o1���	����`9W>�ss��1�]J
�c��dBL��x�O���t~���Ѝ�3���c�8lQ1cj~�Qzd$nL/�$DBJ����'�@oQgΞ@z����:�&��_hh[@$:�s#�v��?��/���n�-҄a���E�(y`�kQ��L\`T���6�/�:R�ܘr�����F�8n�QH�'bޭwn�A�6���7�����	��y����)�蛚r>��!<Su��uZ��@����B�JCK��ލ�����)���1aD���7�`��"�G f����Y�}�̊i��VV����`?�8^q�hw4 �Gc��}bh+=�����Ӿg��7�@9ޖ���-,("�8��-��
*?7����`s��MF��Aa�u�bkӑ�8�r3�Ss��(~ m{{A@�ʔ0�+�FX��sp��J�s]����q[b6���*�p
ӣ�%oB�N�#�>e�u�����Mq
1hԱH����3vqG�������j>���~GE֦�4���+'�	SfNNzr;������B��ނUP�����
�|!	� %������c�� Z�P�����C+Js�����"���-��in�'�m ��뾈�^�i,�7�&�B�6�މ�|��b����n�l7$f�O�	L�
4lpp0A�����^�8��	y���G�4�LD�3�)��Dm�#������C£84)ݍO�:�����_�gKF�Vzy���Z�ݽ2L���Dg�ـ$$�����S�����L9@}^,�>�}D�A
� {#��P��ܝe�%���z�IP�;%�uza.I#����,FA����[��$koF���1�K5(
4%'�����(�֢pp?�.i�o|�V$�UE�	HjR�_�p2��r`���]@�-�346��)�wuuE���䡥������XѴ_�5�ݼ~G�9x��|�|Ԓ�N��%s��|A(B��ZQP�&�]�+*
p��x��H�x�E#a ��(񥗠�A��̘A�.� ����h_ƴ=�SOwC���#Z�0��B�!��V�-��ZC"*��^�03`^x���޻��{_�sy��sg��6���PЮ�**��=F�����<$1�@x����&g�R�����D��A�:땶�w�G��X���p�&�̰�8R^3҈3�AAڶ���&=��������Tl�md ��9��NdOLL�n��7�Uc/Csä?]�x�B�-�\2?�G/ds�r���Ɣ����]��&$�/ɛ赌���������j�?4�>c�!�R
 ���b����:��ZrӁ��-�~J���U`ܝx�Yh���=_�T&�]�mA�>������$ㄟ*�UȰ���dn�"��Lp@��i��--KC�7o�D/>�&�������;�������S��cbb�^�����(��			K=O�E8�ߞ�V�*#����;�V^��GS:�K�-��-YU�]���]7�N��|{}���QVzU�#�~8~��D�2f���#�q���<Ӯ�/:���VKb�]�wN��J#O^��9�R��(u�)���8�f�j���d��1k�������&IO\��+HxC1X���|�lZ^�×U� O����YJ�V��~%!f����!s����u�?>nxv9R�wJ��<5$4�a�B�HFr�q"�㈗_��'͹�����<�#,l�ů_F��󧂌���J�_^�����mV�^�����)l7��Y��	�:%����2��#��;�Q,-��AC}}�9E���R���s�D���(:�����F����������. �X�y;;�.��E�(��� &�����9����� 8E���0+����[�>���hh4��}Tk���C�!,��9sm���T&1���<��I�}����+`��>'\�!���9���w�X��X$�e�������2oE0 &��e+(;���8G�=��P�F�al�ii�
���Y�ZM˙�9��Q�G�����Ճ�SZ?�C����w+++���#|]YYId����Pv>��R:��\"�� cmGG���̔��_500�Vp!nnn�� ����o�d6�p���b@�<���>��k-	b'"���*Vy�s����&�r�h���ݻZ��-�RS͕�냥ġ�E��K���e=-�$<����J:ndd}��r.!_\�ܐ�f$<��(uV[����<�r���b����~N�mX�	�?������/±��ۥ�����t�w�@U� V>�~R{���{��ͳy��0�R�`Y�7����[>��Z�E����r��
'�ko����,������Þ�4�,**��"L���3_��냙�<�4f��`�e萷8:�þ|�^�L{���p���p{�T�պf?�����c0��g�.������f�ıCE�o�n���T���fA�<�^��$K,�'���|^[�3�� j�`�[gfR��
D�WF����w��
���=�,y�����]���(aSuk��A�0����B��������8���5��H�����}2��q�Q�⁁���X(�R�F3�����H��066V`�J�ipSc�>�H�mu,B�������l�Ν;<�����onEɃ��x����ZJ��T����zz�.(f�j�-_e|���(�$o��ڍ(?Q�jik���K۪[I�����h&$�����`b�0��>�ty�|g��٥���7��N�WC�A���::�~85�iMi1�)�3=���X��r��X�����Ăg�I�=�{�;V<��c"���xx��3Z���Y��\�P}##�}�ϒ�k�8���LcŬPeUKh%Ði{[ٜM���X�n�3G`Q
�����_�lJ'Q�����|��.W����Y��b\F���b,��=eF&&�S��7i����V|,GXQ<�g���jJ'��gS���/�cYH���l��'���se8��
�	M��Lz"�;t*͆h�1M,.�rHH�~l'���{�?��!���ĳdگ�����x���KJ����#ƬY;f9B�4�/�7�hVh�"��?6�R���5�[���v�r�dJPv��]-��{����n�Y���Fo�f�O��E�[����
��χv�L��Q��v���6�y�7�j�R�9gBt���H����y�`��U�Mglk�>��턺Ї�7�� n]r>_��rHܢ�����j�E�;�}p��풀@\U�L���c�(7��;q��-3RlON"t�+�(2Kz+(3��sT?�߳9�B�q?��ˋ8W��i���tK❺�f�S6G��o�'�&Jy|����~RZ��1oIW��t\�}��ʧ���$�^���,$<[�l��*I(���+�1q��GM� �1�������
�Xa��={��+> @��̛��֋�x��xE�������QKX�f�5����8"3]9�)�7�5|�'���K�^����w�ry�����27�K�=ε�Z�h,3�z�K��#��ŧ�Y.5EMA�Cu�v��b�0�ЍL�ɯ]*�r#B�DU���$4��4v�x��rE]HO���Y��Ve��U˝����T�Occ�������P����d�Q�q�A�h醸Q�gƆ���#����2`-�B�����uu/�sV�a\�+�z^=%����~�\PŌ��n��%��O�J(3!������M�~`���m0���*-}v�ϝ�l�q<#�w~nn���xbe�p�imq�O��I3aAA�fK�������QQ%͗232(���C�1�HK{��ff����R��Y!�+�UB�B� �Z:b�j������}}}�P�f1�~3i@����y[;_&%-M�������sO����{���n#���
<?�A�C���&Y��h�14�F��$c�,~~���g�d�x�ӉB���^�G��ѽ���<�~�E'?�dd<����_�6�w�����3B�wI1</��-�o�$}����'�aY�����a� ��.�3"�j������!!\"�V�-3+r����dv� d�N����E:�cUmKƅ h\j����)]���А��DOu���XM>2M{�\qqq)�s���?_#gR0Q-�me�t�y>~������%�j�Qo���7�5M���O��0d��� �ߖW{-��Op�N�0��HMMͱWic?�I7��Lח}�ʘ�(wn,���7l'�	}!Ng:�q5-9�� +o��e��_~����~��Pu}[[��I3�y�t�X�(� ��|E+��e#��-H��2�q��!!3a:��`_�J������ᣚ�������ZFj211Es˝;
E�wY��ExJHT�R�Z�H|�Qgć$]=��k����3t��O��J�s/CU�c�>|+[����d�b���0R))o����y]���̓` 𡤤��I~�y�{QЛ=�b<��l7�`�끽�j��8�sxCo���;���W�����*��c?�0|?lÚ��-�ܪ�lho��;� Kl�c6��V��o��_�43��:��
���ǧ�'��K��	���{/ji��T���MN�n�z\}О�A����v���%z���=���1�%?ٝl$.����%�-�$%�ؒ�\Z�tc��=�ٌWIJK+^ĺ<�iɰ������^ ����=)�C��SU��!�#�~' "�Bt�14wt�U�=��{��=܊����E��b,_mQz���x[=�,*���'�5��5�헬S��gz�k��\��Z�O�o*��L����(�1>Cup�	�Z��su�2��*jj�Y�.��l���c^?��~�.VGS���I�s��]S:$D���1�P��{��q��o�C��c9�E�"TTU�u����$j� Ny��O�R*���c���bUkfr2���LHUQ���Y�-������X�� �ђ�6�h�,ls[9�X
uuu���.�v5]Y-p[�<ǋ#Ɛ����PQV�[��a��ߗ��i��6WW:p� !�&p��򰔙J�D��7�A`s�92�XA���ܯ� Ì�bqw��>����FNN>Z�:��s-�eb�y���WC�z�y�n&�
!ޖ��2��G|�5��F���R�&� ۗ�B��AvQ�6�h5�<z�訷8�a�A��1av���v����(��N���u��0�[�W�[��:��G\������=T��X����3g`b/@w BS�a	�G�={�bgɑ���N\�^4����qk��F9j�2vG��lI/�:�ى���3� Rd��樨�7�;�����-����n �PU����Y�9��D�7�
S���g?��1��wR�  ���|�I�,��]?G�'�{̾�O�����W�%*���s�/~�˦w�м�̃3��Z��kM��~|$l0�k�n͐����	���j�1�.]�,3S	�`=::����Kz;6!A:|��y.�ı��+�a62k��H�],&-�+�����D�6���q���>����w|��ʲM��SO��W%4f;��S&$�d�L8�����d}�`|�yv~�n��E�z���5�|+^ �g}6�:�G�
���=�sUG�4�V����qT�dFr��y`� �qxlZ��y\��RA��u�1S�6G�Ջr�����i�ή�WՂ��9��'��7_L�B֗\	����m\��􌌐�i�仯*�02*�����#W'59
�R Rï��%�pB�/��Ƹ}�0s�on�6\5�>d&R!F&��Hl�]�/鞃Zos�x�u!ܸ�o�?��x�Z��̥���ӳ�C�p�L��m�5�+�SDY�F�%�V�nt�^\�&�7��*�S����It�� ��3l����0�7�yp0u�ǏPF+�uD�R�S���6�ӻ��_�g9�](E"�� N���K�(�QW����J���<oE������
Ik���CGSf
V����P�ƶ���w������q�y�����*~���J��kkyH���\�f�f�<X���p2|ߵr�V��×��4t|����6@O��B.�`�=�'�؆A#��BTM�	vԱ�{h�|�^t���Y!#C�!@HPٷ؛���>��>���Y�Uy`ֶ����R�p�\8W �dӊ�/.�}O����1�w��u��A��ǽ(�Ӻ�~ԡLZ���`w�~�|�7�G�$P��pݙ.\��v�Ú���� z�6@���?;��-��(�� ��*?���Y��l�8]p[H���P^^~�مG�� R�����'����Qt:==J���@�wɨ�؊��賎?hʁ�>�wH��7��ihQ��`��U b���7N��I.��
�
��x���z1����1冚BIӱ�b�L9>>Pﶬ�/		IC}�;�Z�C.��]P;���'�[|����?�Pt���6w�^h�7Y��4��J��@aP?iE�42���f������94�����"C$s̫����5�P�=��õ�T^e�c�6�s�IBd���:멃H�(��ݶ��\m�#,Ec[��f��|;">�f��haUO��<e:ؤ�A��n�٭��D�����jV��<ƹ�p~Tj�oI>���d#�xЇA[`/T� �vTS ͜>\=un��=�{e�L��n�}�ؿ��fd,�?���^�% �t���t����R��>�@��Zu��a�=�>�||��~�~ݹ%�Q=�������kk �ޞq����G��\� ]4Jq���>~�f� m����1�e>q���4.���$�%A�/;���-�(9�+Y"�F���Wv��ǿ����T��T�v���'��!��Q����ʨ=��EU��a:��aYg�)l�� |A��~�晓�c��SUEE*��P�hn�#%m�_��+�H�`"��ӬPĽjW�)��݃q����iA�x�%JF�g�
?16.�z�
�W*��_`AD�97�f�fte�5��nq+��4��>��{־8Ϊ�cs��;x� �(a�*+��LC�����(��L�Mx(CCG�05�Ǯkl�w�p^+s�� b��ydhbb �|iee%j798D4u���<N�\���ڔ�Z�^N	g	"y��2��V�$�8:2���/G�;\?�r������䍐���J]�\��JKPDS�=H���ttb�����+����A���H��V�RQ��V��32x�ϷD)��i�X\��������	���t��:���q����4�,33�7#9��F�j��>B�e�g�&��[lj�3?77��xϾ�扣,�_��4X���

D�+4�j�IH�h�#Ӳk�;Ah�!���e}PD4��
'�����y�"�GD$��K�^�bOG��J�����%���9p|�8Ey�4|]�j�c����b���[3,��K���z�������ߔ��M�{�����3����~�)��gc��隙��C��n����-� ;��:�;_��t�{�'���X����Yɶ��|�Mgg�ys�8EH=kh%N&��>��]��Z�$OG��ȧo߾��6-p�)����哖�� F����~Ձ���F��x����,������}u�6����ҫL�r���@`��0񸆍���K@�����v�2�r
`��ǈKHX�-���uu!������Y��<�@Nb���I�.y�ß4���1I��¡q8�ؔ���@ZP#f�t��d�ț����T*F�W��~ffƈ�ɪ�����R��"�'��E�I0KKY�C`�94��3�OA#
�ң
<T_z����F󬭭G���FFF�4������ai�gb] [?����ly���8���|���D��b�n����\�ڐ,�a�����{6��WU�&>F6�QlƧ�A��Z�S����J�rq�IF`i��h���������}�ͩ �vA��A3 h419`YX���Ң�x�%i�ezJ�Y{ُ�Gv��u�u��q���4�}�MMM��u״C?}'jp�E���68m�LzON�OH���F VUU���N����r�΅WO�d\h����$.���\12<&�L2�|�x��9�ү��ik�
iȻ�R��������~��O�������8��k���ݸ:l�fAf�V��@w<M#�ZF���$$ܰ���MM�Zu��6F��Wd�Ӓ�z��LmN�������l�hs�Y�ǫ�LO����ұ����]��c�+W��ɷ��%�=����E�:,�,V���?1��n�UoH���y�з8����O�������R0k%!!qe�����A�ḻl`@���
b$rҡ�IG��bvu\TT��~�/uuu����ڻ'��h0!�~��aJ/`r�Xz?u�fJi��F�it�̇���`��z��z�����z���Y+�q'�f����$]@�(J��V����@{�������S��[}Ǵ�֦˲9M�ą������h���M�:##C��Q�8D�g�v!c4�b��(��S��������'�Y�W�G�L4kj:禧�)s���p�l?��gI�'c /����Bh��lR�D�� >���*jjBI}>�Ze��,r�[3@f��A^�L	����]hf.q�{����걖#�6L6��LY}�|�PW��.rB�k�-	r�\Xe�~�嘀S�)�0E� k����-ӳ�����1ܸ��22ζg���t0���"V�㰇����'O� �&�Wy���nl8�L�>=p���ňµ�BE4� ~�H�ݭ������Ϛ�v&��m��}���N� �AE����3�>}cy��.��W n���r�/G�p��s������i�N���7^o��E0Q��M--w��+��$��}U1��Ū<�姃��7(�(nj�W�����h_���-	�~�*��lh��,����� Ɂh\��x���3QM�CKg@�31.��lL�v��Ӥk��NG�>1&%����>_i(�R0��D����c�l��E�S�%me&�㝌�{Xb��u
� '���ƙ/�7iL,�&�ھ���˅�m�s��M�)���9Ki�ugc�˛��I��v���O�#<����MXA�B���8�c`v��Z�2Ѓ�͏������ݛ�ݩ��Ȟښ��q�r��呋���]	_���X��?�/k���)3��(��:������K��(�W�]޴Z�=�š����/*��%~���4:ON�}5�:G��{�W=x��-��t���Js��R1E�bb�kIN��Ϊ��p��{��R��+���xn����t7+��)��:�9B��C�iA�ZN��Iթ��̙��#C�R�y�������ЩE`�ȍ�±�b���u��/|��e���o�W�Z�C)�;X0�J_�  5�� �Y`�~�3$4Tz������h��&K �x�of�UV�L;s�% 5r]�}hd��B=�]�n�"b��ě����^�2{\>XO�/�p�/?������U����m���LV�] MEG�7XfZ]$\i{h�'|~qq1��V�H\2k:;��*�R�E*��C����ݬ�L����$	�x���_I��$VT����Sʠ.�}��E׾�6�����=ˤ�b�D�`�=�5|/�+���1�L�I�[y��/��~��(9qqq�>��aVIN����q��gϞͭn��t-�8/9~��)�[X�_{?�;)��`�A���­@&R��7G���]D~�P1��d��c���j��xᝐ�d*4�3DQ�FCJ�y�H�Y�n��K���hB�'�Y�iB��V��Y�J��.=��ο�:�9���^��Z�Y���=��ֳ�=��{�+�ӢEV����v���5h�::o";���^->&�d N���(���i`9L��?$"�W1�궏a����e�p�2����cv���N�����A�d����eG sl۶m<�yB�m$%�RF�1~~���N��iݘ��^�N���6�6�����Qm�~� 3"U+KK}��Cɜ^�|�wl�2-���
��n�_sm5�+R}~?ȭ]a;M���խjo���fXW��D[A!�� L^����✚o��C��1�Twg�h)��F���x�cn�ea3��V�ͫ�@�VS�=W�1[�6�(%Zn"V_V/�K�򼛛>T�ϕO��+v��!������י�������Q]�n�|�6H�Fz������|R2�x���2�v�{&����ì��/[��˫ԥ�ye�W�F����Tl����/_�/fa9�A��ݗu��X�=���@�� /�`|L䤕+Vt�F�}�m2[t����П�����!Oӷ�^��T��[�04���-U d'�t��C]�Yx���tR��f�J�)YPc5��@rr �̲]k��������R�ng��{�3г���H���]g%+���S�{�u�j���˭k��]]���
�9h���Z��~�E����P��~����$~���w^$RW[��������Bo�Ϗ��Mǖ�^2[��D�����?��u(�ſ��233���}��-fƓg��O�ך��>�����k�j�|�{��}zTz� �s5�U��?,����W��N���ލo���{{V-	R�q,Z1��P�DD1��B�T�#��܍Lc��:���+<�r~Oˏ������'O8�
p�y�n�֛fK����Ր>ׂ饾}T~�< h�@���C�� }3O�)z&�q��А���t�2H��7c�x���~��x%~�b����YR2��G�o՗I�F�˺�B��S^��`W��y��y���䏐�t�SP55�L�v�.�1~�-2 ����5�e9�YR��J�*�|G��l�6�Ns@MX����Ǫ�Ĭ�J����t������t�LR}�uѳ[�����,���l�	��@1ǽ����J�>FEw%V>���GZz:��C�E��8 ~�-�4褗����ֶR�_��nT��h���UE w���]��C?�!v>�n�d�C�k����z��s[��1Qo�<�5��_�	(*.����1V�t���k��FD�����O%j�/�@�K4f|||T
A���6��/�Q�XQud�\������
���n����@��-�IH$�%8�!*�9�uq�?A�u��	4��ޅ�S�$C�.�_YI]��g��gQ�@�r��
�PV��{M5�Q0�1��!I7�NI�RɃ�6�<�x��Zvvv�/���}�C�����QTTԣӑ������^/�7V���T��*J�ض�O|f#b�Zy�X���Ǡ��l�-�uu�ϕ� U��1����lr|�%ϽG��*9�����p/��}x�T�����>���Xy�&�h���l]Pv�\��#/^SZ�@Y�~�+d���t��0ק�Ŭ�[�8B��f͚5�����1�9�w~������Į��a`�i�*�3>%*3��~��Ԃ��4��*�"�MM�C��#TK�S�k�轭n�����\��U��J�.�jP,�����h�։V�ǿW�k����sr������f�̋-^[�>8%���f���D�V���!��_�O+**Z�b1����>�Q��_����g���v�C�~CƊN�_!Xn�����Y��uTħ�R��6�{��,�11뇃< Ӈ�QBq�q�{������X�<=#A��錭��!��#6�t����]>Y�4���W8Q�^	Y�E7���}���h��4L�P5�O�$�Ƞ:�9G��h唋�%nnn0�D"q�3�a��q�l��~�ePYW�L�ʚZ��ѥ?'��Ǎ�	(��z�<���q��b��:!��W���s�b��~�&7-��OnߌMi,פ����p��aze�U�.��¡L�	M#��F����c\��3��4X̽�Ƶ�.����V��K_��ж��w��&��{Oʏ�ܸq�WH�`ҟBϏ��|�����/���R�Fs�)�����r�	k��N�x�.�ĖKL "�F..��6q:,��z8��v:�Q��j$u��W^VG���t�D�}}^���܉k "��j7�?���ac�n~kz$�Y a\��Ũ�N��M8���%}�"�<�Sh��{�)m=@�κ��)��ҥ�k<�C�^�*fG���jV�����-�9@�E����Hス���ǏAm����Pz���Jn���#A�۸iSJ��j�i�Mר�h�d��|���e333Ә)����l�t1wN�w"�a�b~�g�t��|����ml,���~�4�KxB�m�-�ߵ��$~���c?��������=��|T����J���b�}�>�C�9� YR�k�*H��
���g'#����աq�.$���W�x,�VRR2�i���]5���u�t"�ENm�V��4�����g��p�Ѧ�"���8�)Z�B��ӛ�>��?�.��f��:���:�O���)�Sh/���=�����|����1�
�A(Gs�����zgQ���^ul�,9�n�~�0�������B��Ç����l���4����*n1{��C w���g�
÷��]�v�*���*�~|�

"�km�N�u��=Ŝ��,t$*�������,s��kEa	��O�v�:+�$m��o�}���ѱ�{����;��]�Gw<W���C��mrIގ66��Y��=i��:�H0�P<:s��`��dS&��N��ڨ�?1q���;��4�B=[���˗c�8�0I�"���nڅdY��q����Έ'O6@�������]vko�e�R@�I���*(�7�Q\^o}&���.�����H�S�5��Y(�])�}5L�iP���]��#;�w�ccբ7�~�Dgg��M�D_�h����RHTsg@�|Z�WE	 �!�"P"��\�vM0*H����6�F�_�<�o$���E�P�qM,���
*��+����&)�+�W�Y��U�F.�l��P|���T�[�FG�!oٰ���*���XdMŁce�WXL�
��``FT�f����Z�%��X\Q�_�8�Y@�Dhҿ�;i�5�	����Í�w��RE}�$K�0���Ϸ��ٛ�::��>�YI%B|�=��ܶ��0��&�7S�C��Ϫ��D~Z��8�,~�,����ɡ��R�hNʽ�:Ff�s
E#1)��]NZ�fJ���f0-������Z�xr�ӧ
L^�C��qt\�s.$w���� s����,�p�m�{g>Pu��صV��eܒ����4%�q<�t���^��EU�gve�������l��-����q�YN||�5#��O�[[/�5��
����m�\3n��_Մ:
27�|�����H�6.V� ���Q��e��F�u���0`�6&����಍1I������j$R�=nq���nxt��Kv*�kjjR/t�6bvoF/}��B�x9""���/j���|���R�:@G|L�]T���V 4X���<�t��#E�OZ��}� [__��[�wS 1������Ȏ
H8�3�65���:uwPYt�����t�BtC��kb��3{$���b��W�f�s\�,���&'#�M?����h=��[r_gō��2=lܾ����ﴒΓyw�.7��x߳zs����<��O����ٹ��'�f���_k�2�z�ȓ���q_>�:}�כKm��ٍ�ο/�l+5K��� &M�A/�v�e��Z�}�B�!�~o��5�ͬ�=;���E�t	ޮ��6T�O6Bexb��8���WUt�W]�b�ϟ?��탿C3�&�!.�{r/�K7H�H6̻g�H��XTL��\�0�1�hYhX�lt՝���b0/��ab����mTӼNO$�6��;�o<lڴI�wɛ���֢>?��R�&�������g�����5݃#���~ű�zw��*憫Q�<�����U  ���M����7�GR��7䲠��5��+ ٸ���o�+V���%C~<���DhI۸b�`��4��ArG,���f?����e��A'.�uX�;�=S=�������~d�P81��60 �$��<^�a5W�<V�5wV�%���g�n����b�Թ�"��^���G%�:��vH�A��W�o�� �.4���͛��Մ"��+۶�7�jI�����s�>� ���녚�����$W�U0=��F������{��N7\�1KEo����Rv0�� 0�\��Ӫ*M%�Ƣ\Qā��y�~��'�7����B,����v.Xk����j���F+�$��4y���BM��C������hD}oT����Xxcd؜2������孅�����������d��u�'�0������w�SbEm6�#5Q�r��g$�\�$ �_��X(27��'�Ӷ�l��1)f�ak"�{� �[9Ւ(0	��&��-4���M�����8��$\�i!/�9��:8:��? -zخ����yy�����������{5�_�*Iz�4<5ԭi'�fҤ�zC� ̈́B� �s5�e��C�o�C&����?�oMp�/J��-�2�Yfә��y���u+�����ՎX4�E���k����u����q5�AېQ�ɬ���<��e�MB�x��5ˍ�L����QuJ+�����%�o�OV�r7�n�4_@hX{"+;��g.^^���{�J�宵����6��U�����o�h�;�p�%i�� |`��r���Lw�<!.Vko�ת|�l��7%���N\\�4S2����@ݠ�X�|��6 �<f�k��3�%=%l�NzOH�e̴���HMZ�M�7�d���o�k�:�y�ff��=�e[��M�M:%iL���'m����$3C!��j���ߔ�G��4/����LP*&��#[�L[�|�� �u�U�;��{	B�0U?�iQ!��o�%�v�!�I#���C��=��O1������z999d ��V#�:�>I4�s^�о#a��Gž�<�Q�jo�#�B�D���ߎC\�m�x-tE�����"�����F��l��5ݑa��9�sG�V!e���헃�
[!����'HȅN���H����&���ڮ�v���P��TI=W��ۜ����$0���2���O��O��	���Aw��Z��m��Wq��s�F����*�!
���OW)	9gut�NR)�N4�ƊŞ�DpHXX�]��B��,�Ѵ��g̢�R'�$z�]d�z��qZ7��ll��1�������6��_� �p;v������t�fټf���>� I�9� ��Zvc��NـK��m�cŤ���=B�V,��-�'����߿���F߿Q��p3z�����|�351�hDI���ېEYXXl�]�J>�
>H௩L޽Y,e�����o�����ϛ�jo� �>�^��F�m���ݖ���h1X�䇢��4���2.��yr�ѴHک�|!�V�K�EFFV��<�tjj����WΏ��UyB�m�v//��h�������{'�"?��^�fS&靘��h�u���8�X�����ޓ����P��b�E�	;�~��� ����t��
to}	B���ӏW������_e>��G���A|m?�;��al�R��OK^��#1�~A��e����4_�$�='AX`�K3�$x�b�\��#q��3��=t ��
�������$�
�&ל��;t6�x��$t�%��ˣ{�Sp�h���>���% �?(s-�ԽbJ�L��q6\
�[/���*���H���*�hs<w�T�2�ߦ���e�"�����h�֢
��Z߹������/�t#;�˙��9��!���4�c=���if��}���c=}}E!�Z� ZH��mn��!Q��[��OQU�3w>$.���2s��XrTV� ���zo$��p%Y w�@��� �:�����f��=1118�g���i�/�il�T����D�n-m �>�N9��X�B2��ja[��"L�����%�J���O��\�����D䱁'`��Ā���/�{�b��v(?A�N#=:��h�ק-����қ���~��A���r�g��2%o��ܹ}e���tw	@��$H��s):���X��N��HKKS�Xв"�Z���*��I΁YP){����c7�y�c��D�����pby�ZrM!��=��� ߈Y���+�����F��Yc������2����@��������6/^���[����0�����9]\\^ggo�k�4�	&PUU��B��\7>���H�e�O!?<`�z��P��@h8=�.�lQ_�eCI:   �>��3�?p�^��v���雒r�7�O����`}���#@��\~~�S;#��橲���=(�!��8��
�%�w���{���S���$�w���;��;� @��O �u���ޮ��E���%� ������w]�zn���$'��#�h�]�Ҕڜ~�w�~�.@R<9���#P�Ԡj 4�yidd�U����Ք��j`��>A��[��AF�#j�!��C8L���*p%栍�a����w]�	� $F7�E����<�����Z(�`�U�fA��I�cp	���g;`�ɗ9r�|D�_/]�͜���H��RQGJDM:p/7�E�L���ӎ�v���Q�Ǖ(#��_�^F��|4V���C��y~�GHL���������;��]�=:���� �ֲ`�J�t�و�q��iH�M͏0f��"�7��E@�i�����aB(ף[��F�ggg�NIiSw�H~D�@��#w���'~3KE�p���X��#*@TK!%�5���!�T^F_f@��@&������,�ѯś�?�#D
�Ի
�84n6�#�IW���yHYzTy�+��
�Κ 2ˀg�JJ����D��u���@���r��\cJ��=߅�|SLR6�K�::���k�M�2�3��m��Ex��,u>H��@����@ ����T+��E�(f��t�������@�0׀oxX]�[-�V}���
K�6 ��+Qso�����E�Y���������fS�����U
i D�p��I~l.P�>�:V��\����t�[G�#��lZ�.̈́8�>����F�H7�8�$%M� ^������q�v�q��֓t�*I��*�<#@֐������n�K���Hˍ^�O�k ��W�R�fl�X&:��'������ad�]Uѯ32��_P�L6�ŷ�VVň����V�֜P,�eKǥQ��P�
ڛ��kH�sD I)\ʗ�L� ���n���S��߹[��n ��y|p22Ǘ�ߺit�u�7%K&:��\E�[vVn��R� ^ �|��ƿ���C��==�WzE�W!넄�>��1�V:���p��U:e
��O�i$ҿ���Ħ�êw��}�l-T���1�5f�K
�N1��zR�u��$==-]��d@=2�XI�!<<�f�./C��!���q�\�&�i�l6�������5��7�t��������_U�������\� $�E�<�]���"�<������t�廬d!�B��Uϡ��=(_Ƀ��^�'B�)��ucTkƯ�zݿ�.Giv0�Y	�--��`��F<�u`@Ŏ��p�F��^��BAY/L�y5J�|��-�x@���۵(�itH�c��Y+DPd�`F��Q�����q$�ҽ�%�c�h�&77���l$�)3�@��<���mX�=�	��sXpɐ�(��q�&����ۣbmpl��Dt�LdY�4Ru������:��)H���B���$���S 3��_(��Ӄ@/���$�ƅ�}�������MdQ2uuu�zrss��W>UA��V��'��s��ZL��_�ta�#�𽍖"����� ӏ���;{���Т_Z�z����L�i��������z�p�D{�ʻ�A��*Fx�/i[:i@��PՋX@�ԺLaj�f�A���ڌM��5� y����kz��~1vv�҈�f�R9����Li���+}j{�zbں5d�U��U~� P*d��VB���<$S��sj�|���r?@3���^����Ѹ��*:�����oL�h4��Ż�v����s\[O�U�"�u/��mP����/?�[(�$Z�����mT}�&�`%�T��e%��k0��Ç/XX����./�<$��$�M�':�P�zMl.m�M�F�В]˦PP*�
!�|/6cK����9Y��Z���'�6�'
�H�Kx6�~�ƿ>B5V�
�,�S��N\��zz��b��S�NA��������m��R,dK��h݉�D����3�\'�*�̱�q�y�[�Ys1�Q�A�(��8�C�jM۶��`oOK�t�re���c�]=��/�ӈ��6����c���9[jB����������Q��Zooo��,� ���'���(�Y�N�\1�Q�>�}�a�aE����C�Pa`1����X�r@5����Pg����m�C�9|Q4
���NCCw��!p��O�|뺶��MuU����V��]s�E�B�օPf�����WiƝ*�p�9�P�c����Pۻw/���Θ�������:G'*�iR��' �_�H ��L=�y��ә~
���z�ȏG�c�˰���2Ʉ�X�����󮀇 Ę��y��5��=$$� �����d-5QT�t;d���64����/��W@EĬ�e�M�6�'��9D�� �4Z�ԛ>�Ґ��ⶒW� �9��}����T@O�}R�����҅[����PG�S�w5��:��
��@��yANW�(��sp2����_��Z�	���4��
Ҏ�԰���;��37o��տ|�r�$��iG�n>0�}/@��$q�3	����Y�b~��Ŵ@��.���s���(��z��2��(��םṞ즡O�t/;�z���ʌ��}��95ONN����%�g�i��xH���$��t�4�����F_w����+��ď�y���OG&u����{�v��#[lA�`��QH�NÝ*��a�vV%Kq�Y��i�S��Y0�����pat *�rDq�66*l!�?�so�
�E&*x��;��èbho33=�?M��VA��ϠSȼy�" N��::��$5�Ԏ�L��hAC!aax��������
-�))�z��������VQ' 2���3�)�.���n��}Tcע/�@U���)��"�>h��0��w�m��l��}l��'�X��U����DQ@׀�燺��~f�� ͷA|E��u^�Իz�\�A9�@{ie!���^�9g!�F��-���N��V���m�����Pe�/נ?�EݧŪ $�
�h��o��Ѧ	�}[[�6-GA1e�Ж�7`����%�y�oDA4�J�܏J~��֡r�w��`�eAw�n�U��c�aO7��<H3Rh+
���$:�y�R? &HۈŹ�[���%��o��������C��h�җ��1��#	&z��h=L$-=�D���h&���Uu���9�!��բ
| |BϢ����������	�DM$C��qdn �3�M������+ShfP9i(J�l)������:����V�� ����𑲵��E2��xI���"�%�=��=��
��h��F��NII� ?��R~d�ٷ��[�r�Κ-��o[A���wݻ6l|���F�'1 �C5Z�S�6���NJ(Ix���px��+�6 %��_�~@�D��\"*���p�P�#�DA�~��̙3q����� �$�����Bݺ��V���`K ��� v� 7!�@?��}��IE���9#}�w��&d��Dx���@�/�w�}Z}�s�4l��!g�d���
=�C����γ�o�:m=�w>��}���`] \Q�z�"�� �@��
)�x�PA��-.ix�[�e�7�vȂ��s�� �����f���W���D����^DU[2-Oח��P�N�u���ٰ53�Dr���9h��6�_oq�ҽ
�/��;��Яs!G0x���iՒ�o������8��Z`��|XG`�[��+���Y�*v�*Fw�
,���m+����vvB����y�o~��l���$Rds!���
zO[-��W���&%GC" �!W���0Lu�F@��UY@��G��s����RT݃� �A� `A+ kNHN����`5��C`F[:���蘪	���`zE}�2y�������ޤ�K��������ab�A�Z�]ꍾ:ea��;-+k�4
|�m]�ȥ/R\�jq�2d����U�o�
�,T�� �DD�w��Ǡ0)�l�i�s��R	aL��i �/GNf��Y���hi���M~ŕ�U]�#��s�=����^[����P})PG|||���е�%���4A���谿���A/L��ҧ{n��� [��V���V2�oiu`c�@�[�%L�DFtA��\ 3h��H����}�>���~������6�mk�~�<�=�P��}���y���>�6���V�E��[�[9^ۥ|�l��X�~��haa!:������`���v5�b���`�ԃ� �4_-4�2���YX��W�Ջ����b@�M��!��T0`h*�c����㗟�[O��� ��7\���y;1O���X��TU}CCïz��e7?"ɒ�6(	`A��]�/}�xA���p����t5�p�r�>{l2�EŅ���̒t��/��M�h5��m���[����
w��/<��%,��7ȩ��&���=�F�y��������!ˬ½rBd_؇{Va�u܅&�5���fw��3kW"+�|L�:Eu$�Θ�>�3?�Q�Og))Qѱ�~��������͔���O�d����*������M{W�reZX �Μ�9τ����#�y3��M�,�#ˬɜlҦա%����S�h5,�:K���%�����深s�2�3|�h�V����c�(X}����%[Q zG4|M:sz(�;#7���A�8�h�8�]��K���,)�%CP;�1_��F\�8�^�uN�i`U�����!�Jg�:�Ƒ,C$��c$��^Dr5F�
H�. �Ia ��Eǥu0L\g�5��L��%xg���Z�L�4\����wFNM7�z6����K �
��;ܕ w
8��Owb�]
������0�>l���3�[��F���̓r=p�r��I�Ϛe��^��;�L���⦻���`��܋{R=	5p�r?� �I`�6��|�@=xX�ql�z�l��5�����Hr�Sn��-f��'�?�`�Ӡ�r�jue��?���A�Mw����,YƦ������VC�m0�P��П��p���:xă��<�'��I-�V�E��`����$�Q5B̳��k�����5)\P@�z�Y(���@�M'(�{�a̐��&�P#;��@O5��5�.V�F��Ƚ;-Y2��!l�<o�� ���&``���P��}Lj�,6�G7��;��)�}����ܛ�]?�3� ~�0�S��A��NO2�f� ^�d	�Q��1��la܂��:5�Ђ�p�B�Q����Hg;X�#(�I�,�U^"�ryբE_ާ�~yY~������	a�ˍ�'D��ě���n�7���^��bG�����%�7�~1�f�}�x����{��4/�bhc�'�lw�x�����<6݉��>�0�U��Ln#�}м [�aඃ�+>b�k6�d�~�m��}��,X����]�E���Q�o�Q���|�:v�(�K=�gZS��x��Jg.���0�\.���a��;��<Rs�9�`s�	�+�0F�B�� ږ>��C�%����дݡ����]�G��ׁ���8���@��9�3q���v)�tȶ���������J		=0OP�X+ a��9}�h����A�L��=A���ى�<�Q챫e�d�Ŏ8�_Q�I�Q.VL���jN_�7�=��+0�1�1��0#r �y`%6;s���6�[���+�n(ja%�b���0� ��-Xo?PhK��3��XC��8���P."�c*��jw �|�qr0=g��<��D���9Z^�q�8�1�uI�  ɂ� M{� .��b\�(�ԖJl6���<L{=�E�� �3B̯8����A[ڠ���V�A�F�Pg���A�0�!Ѝ��y��`�o�F����EY@:�X<�A*���C��zй�GN�1ȡ��=��������64��M�]n�`����uє7�O���d0�1x<z�P�I!xyV��z��<+-���j��G���!~@n+�ۍ�J��7���6z� <&�=�=���[�<�#��t.m*hT\[�=�6Nw���2kAL(�H�2��[��f�"��K�{Xg��,��)�A+`�3�rK.�� 3L���<��1���$�G�5�&*����a�%
3ʑ0иBἇ�\�t�� ���'���=��@�w�F1�-��߽��y9D���}�fl�ϐ���V��F&�̂�l�R.�}������Л#O�4�ڽ��]柈��-ւ��h�y��	���롣7p��!x,�ėNK;���z���Ή�)����߀��7���o����d�|��,������o�����?Tyß�m�$��q�M7�����W�v�(���(��%�mp���Zv%����.����)��<����1�R�25.����w���x�,�[������w$�R��@X%�����~�O^��v�����*���_ծ�1���#��9���F���,�o��l,Y�x���nof�Ϳ��:���������՛y����d!p�la��"�LK�:�I��v�\SS3���o:{��#:�rqq�`�s��U��\����w�ȴ�`k��+&ѻd��;��`N���І���C��&�ᶌE�mĕ�\W^�m̑'z�Z,�;z����&����f�u�3�8^��4�V�naU7����Q�*e@�1�
/PAGq)�-�w;,Y΁D�p��Jg�]���HB�}��gqcK�NgN��2|;<��eǵi��8g���4���ma�mÿ�o����2$.'����G�a
�Іی?z�ؠ���NÌq��|u��_7 ����m�9���^���#�����q���pM�ΞH����t��vVc�@�hÝ"��m��w:��NK�Nk����V#MK�[�vǷ�:��9������fh�yP~��ݲ�8ۑ%|]�Sja�q��Ƴ������#}a�7�3��mE�V�ZZ$U⒣��n罠��Pb���P �X/���FÃ!G�}�AA�����xP�]�{0�A��G�8	�S�Ծݚ%w< ����H<��=��u�ʊ����ߒ%ȟ�ݲ7�r9��P9T��n��Oa�5�!�ȴ�
.��~\Hp+L�6�nq�G��6�U�� �5@�G#XA&��0"����x���&���cp,���~���ha��Ex� �p���J�����v`j>�
��aj��=(^D�8FG5A��q<m7�m� ���Q$��ë��r���fl�0ƅ ����	�@n�	�����6�{���XW��~8�͒e	Lc�6�9���K���/��w��1�P"���k`���Jc�KnN��cx:� � ��Q__o����]ϴ`��v���?Y�$���q`�3fc-���i`w <�a
{ (�<�Jm���A��_ ,���n�%�e�EϘ��Ā�� �g츶�І�ۂk�!.߇��6D����6"zH�*�6D�w��:=����:��6f�m��D�������w������^_?�Ӕ��ǂ�ҟ0+7箯��y��E��������(�F�1�^� 2; 2��d���5�hǨ��D,�n��q�ȭ���]n����[,YZ$G4a�J"��Vk�� 1�� (�bFM�F�:�?`Ѓ��..lv���`dn�Hel����Գs0�	J=y�/=��a=n�`(�l#N���"�K�vূ�ԭ��у�@����"賥����v=�6(�C����{9@�W��a<A�@�ژ>3�e��(k�G��|sB�������2�B��`S� (9C1�W��NDp5Fp��>�wb���gG]]]C`>�!�%���b�3�][oς�bzр��J�`��w�L����T�
q��U^�D���Qah+��]�U��GU��]L2@O���6;�:���M~�; ��,Y�f����<"��Wɵ�}455���ߴn�q�EG��)�X6fa������bbډ(?��e��چ��xR���� z)y�$P`���*������	j�A��Sy9 ��0����R�|����� �P����c��)*6"h`��I��bn5����*�
� #ڸŚ�q��gv���-���P�ȳX�j|�k[�� s=;���$�`y&�z:,f+���0��5g��C뮑n�����c����%����|J��Rn�W��S�qmm�Xk]��̞fB�ۉ�����؟����F���c8}���|�Q��׌'�e�u���E�r���i�K<�$�Ý"�l���g:��%䌗|��Sd���c���D7C"����_$t�2��z�J�?}dE>�������Є�O2�����2���_���+�ꔈu���?+<
V���4�㿎��u��(ϑ�2��&�F��n5ޚ(�}}�ʢ��ݷ���V���\�S�^�����	��U]e՛(&f�O�}~v�Nv�Ԕ�?v�:^`m��v;d�jSM��#K���G'&���KM�.}�Y�<6�wf=�;@��j3o��?�N2��W�B��蠣�YV����c���7�A������p72�ѡΧU�5P5�ᨤ�&Y�ώ�d�mQg'5��Cՠ�i$��rO��믧����u�	h�E�'��1t�4�fK�R�k�{�>��A{���n�߄PR��$���I�T�W_=/�g�q`�{w�E>�LmB�"Rܙ�?��dN��q�ĭ#S[&������yǑ���\{��ә�C1��_�Y��/̮��aN=���d���=,&�!�a��"$�
�VX�ߜ"ߟҠ�����0q��lE�������h���T
��B�"�������B��_83h�DPVN�?�<�I�[��ş���*9C��Tiq�*T�|�����R�
U�lg`x�ƈX���t�r����x���wP�T�7v��A�aC�c#"����j�_�:TX&��hμs�g�Sf��w@�X#Z�/��ԟ��Z�P�i�y*E�"��k���4L5B���Kz�%�uӷw�7��v�t�,s9��WLE�7)ͺyvq����J�.?=���oi�xs���_?prk��k|��G}��a�
/+�C�ŚV��IDC��wޢk�2��ag�{��?Q1ȑ�����ԩ���mV�Hځ����>:S���'JL���3p�}P�O�?��zvh��l��=��V�Q-([G�a�\�^-ꬦ���u\i�@���-q*�z�2�T�Z����n@S�M�ۂg3��-)uFa�I؍Q��#���@3�pJ՞ZjW�����d�ԭ,���(��4�"�.�(ƻG�Ѷ%��c���,�!�!�9u&k�d�S�'�*�2�R��s/���zn"����Zo�|�d�5;4f���"���db�fMigف��$ܧ���k�f��>�x�?-)����I�y)b�N^���ՠb�㿨��ء��rxF��}*P\�雓�*�^v
��k9CU�.ػ�.�k���1pC�\x��v�eӡ�R��88#$)G(,q�Z$�����z�V�7L(��.���6���&n4�n]3���'�숓9�5rr�oRs(v������X��@���8ůT�%��o&>�S�0��R;�z�!�1�t���ܤ�
U\�a�m'��IԎ8Ǘ�����bQ��L&:��L�RT��_��F^�"n��ݺ��{a����xn�Ȝ�_���V%�N���U(�Dq�հJ������B�k��$��fe$��3x�����cмǌD��m4��Rg��UrS洄s��W�x���]V�$�H��տ�,Խ��&;�j�L¤���J������I�(���g�m�#F�|*�)�)��"��t���T��x�֦u�J�12��<�A�]��<�ϣ`�ie�'��W!�Lt~X���r���[TZ�ckB�ǉ��q�8#��Ó��s��?Qct䘼���JgS4F�8��w��eD��ΉC?�[iB�[tU�M�&>��^�넦Nn�w�7ڀ�o.�k��{{L��I���Pqd*ى�E�HjV��	�7����K,���E�k	�yo�L�mr/�-���Z_�jo�1Ev4�}�3fI���o����s�د��l�zpb7HW��E���eP�+r��z�)Vገ,�/6W�-)�������ɚ��Yo�?��4����(d@o��|�J@,{uo�h)�9�2@Q����ws�M�L�f�(�i3Pg�ӵ?ko��8�5bQȋ���Ϧҕ�Yv�r��HRS���ki�(���g�a  }��Ώ'Y�ޟ�|�ڞ?Ш{��M��X�$����K�����JN,O0P�yK<fok���lG�w���IW7��LH2[�Br�>���0Է?���SY�9�Q�r�VO�,����Z����씬����Ĕ���觢��r�r<�<.>:��T?��\Ú��H�g��2�zL\�yp}_1s�����Dt�K��3 	!5Z<��x���ZO���&��;���ニ:�}+u����1�T�<���/)+f�!"ݯrЎ�>�^��!2+͓�w&N:~DQ��T��)C��k��ҝr��UU�	��`B�wF�C�7yh�H�;�F�+�)�(�q�u�^�Xj��=�휾�L�0�����=����j���I>�xd4�,�)�lL|1����e�^��ߓ(u�����t��?��o�u���4��` ��3�&��b':x���'n
)^J쬾�('+#�]#�iYߦ�\��2:�� B�iTc���Zs��
/E���lg10��})u�a`D�Z�L!�E�J�O�� ���P����J��r�0���%ny�a8]�r���������0L�.+}\��?�c`�a%f��C�F.u�^� G����1Rg��r0v5ҍ	8�D|J��.�� �e`@:S��O�_�`@���������J�q��h�d�.�t�F߁=��=#:���Ga�?Ƶ�s���e��M�bYL����0!�<�R����d ��5�����\�\]�0��)�i��:ԟ�V�Iz���x�*��j���l��	�b`#=:V����g=��j�b��Q���<�~|��{��7�mUթv~ף�2�Ա�r������dz����NM�d@u�����b�Pg���ݓ\nka̾R8ձ(C��<���{��fٷK��� %����bf����K]�t�����qR�S�t2�g ��n�?��w�T�&yA��'m���F�~.��?�Ni�I���K��u�{oˀ��5iyq3:S?fy*f Q�3��U�u��������P�;��ș��Q�nC�72�zs������ݮ�e7��? ��>`W�-i\��:����6���!�7�m�����M��%���5�����c���Z�z��Aׯ��0&W��{���mP�7��]Kŗ�r2 ��rq�q���ͺn6O�̿i���#���l"#�?�g]x�e?���j!���z�VMjV���}#ī�|�^���K*��dEi���_�>8��4��:��`|w���	�K;V怳����(�W1��Qj���´��L�x���G��1"U�7��:�WԽ���ok��NPn&Z&5k4�;&��F�,܆����ɖ�3����rnvS5"Z�A�{�S^�m8�"Gef���.֐NsW2�f���?O\��;�_�`����
��4���F�)�,j�T��ԯ�}�3��a���Ru]���:N}�,�J�0\R�O��8w����1VZZZ.lN5gS��9���Z�=5<�;����;�đ�߇����E����Fø�/������d������s�����[�7���
�%zm��9�F�nJJ���I��T�ʹ�H��{`v��ѽ�\�NB�%�)�rr>2\}(�ִj�&��r5z�յ*��n��E`�O�Z��5N����@���~��ި���D)�)��oY7�j��rF������]��l�xy~�&Y�u�۝�3[�.A�ya��z��B����;[��X5�,�LS5����%5v�j�j�7�[�S�Sv�~ qb���늶�0�=������-w?�}N�p�	��M���2#�w�{��Ӝ݇�� �vt��Q��u��6jd���.��5i��R�6=�
���WIA��K9�YVBd�[�G)�#�(�{9W�UdI��fxh����'�U@b'C(u�R�r��S��,»7x��ʐ'~9:�fg��;����y$����:�oW(�(���yv9���Җ�Gmn/����6jZfZ�����	`�^r�F���̰#�U��v>v����L��Tg��a�MJ��+����I�f!⪄������i�I��bW�7k�c`I�E�C+�<�8�N���c�0^�p$��Ҭ:Ĭa:K��+�O�*3��u�Tza�d�3���)���AS�ī���?�t;Įo��e ;����k���mrl7����AkS���9�_��=71�$�Zu��ඳxBgH�a�)�u��R5�v���U=��[�f�FzY�s39��D|�:�\������X�º�:����q3J��x
�c0WY[{{Zyf���@�.^�¾Q/�O~�JcnW�Y��V�}O火K-�g)���,פ|Y�m�h�s�.�I?��Ԟa����"�2���s��F��w/.)�I��[��C�����B����Yi�m�@0W4�جW�A&�jC���Z�4�v��Û�1�<�D�ב_܆�Lx��*���5q���q���W#8���>_��ܾ�f,�]��G�c<Xte�i���:���5��%o2�X3�%��i*N\�-�%	Qk��;��z%o⽞ +QwD��OΏ'���#��Cuݜ�,�ň��*�JM��iۤ2;nQ��ab'�����x��db��#�������0/I�y��j�X%��q ��˰����K=8����`ͱ�׶�Ę��O����)��P��R��{�N�4�� ۵�ô���i��
�FŞ���"+�<��ˠ�o�o�T;s�N��63L�����J�먓����������"ý ��#o��j2���|L�C��`oo_�' zb�|·���
eѠ(f��n*ԡL�g��e�~2�U|b粰ӗ�9�2���/۫���8'yʱ1��\�꥕��v-ɻC���3_�EY)f�e����=����=����/h���+�Z��b��V�S7���K�gE@�!�"R@A�a	�X�֕Z[AP�%3!��HXԊ�7������|g��=��˽7s��O:j@!WN ��rDb�c�����Ȧ�0G��FI�ٮ��뮁\XBWxu.�L��,ۄm�߅�X�y3��W����_i�׻��ٸ��Y��v+�i;k��gd$O}T%�Ti;�7���]0Wft�O��w�J�5�����ѿUv���S&�nI"ҽӼx;�\����?ȱ�5k�d���C69��cUz���)l��&�f˜���ܥ^غ�*�N[����F�3��v�O�a�V9n�y��y����)����'�ކ�o���](C���m��{Yk{�禗w=ݕ8��n.����-{y����լ�Q��Ӕ����9G�\ࡴR)��G:�t|����e�&D�|�ѝ�;�Q�����.��
�5�YmVP��#�aa��d�֩Y��OSo�5d;�;V)5�cteI�n%���K���낌��C6��{AD;��$#c�_�ƒ~54��m��D���F��Z{��`�*��ȥjiGlXM�*�U����b{�"��	��fs��%������������k�g�+f���K���/���^�j�ϩE����K��s!>�/�/�j݉���k��8^��z�,���]WIxs�:B�q���dt�ő��Oޥ����'�����uȚ7��"��7|�KA�B2Ȗ78Gܲq{�$1C�Į~��8���v�B�u$=�I�<Ų�Q�w�,���gB�6��d�w#��_���re��<H����Ir(Rv+�Nw]}�x
9K�8�N��kJ��e�X}�F�r���*��D�֥x�؇Dڞ*A��s[[��9b�ӹax�б]�B�6-�ZR(3�a%��Ʃ���*{���j���6<��sE�A#���Un7_�k�6�U،����M��y?���|7�WP/�%��j��YD�9�=e�*�ڛ��;�mT�R��&y��F!��\���=O�(��>��q� G1A����Lk�������ӻ�kB���GtVd�_ݖj�B<��IcӇ�<yED�|º���TU���: {0�+�Я*OJ=x�DS��q����,x�m1:���K�<��@�3�x��6m�
9�.M�:7%y��[��-|�z��F���wW�e���%��C�k�ۻ�a���Gy��5�?8�hp)�3W��	��˜�k$��y{�|l9?��=�5�E�!��-ݎ��̎j}��@?���6ͪ]�����y�b2��!x��+/�$E�O�2�z2|Gz���r����{`���<��_1z�nq�/�ڎ�zU��}��������$[�/���������ks��Y�l���L������Ym���ԛĎ��o/�\hd�in��l9������G!b�#����&oN+(�إ#� ���\G���S������)���&�X��6S�LO!�X]�\I�����Ǥ�fo����eP���Й׏��рt>K����r6��t�ذYr?v���NӘ�@�<!�
5�'��+���p�N��^/��C���䌽<��R4� ���/ׁ��Q_�fɪ;y�分V��'�0,�����cǸi�Z�e�q�R]-2m�:�V �7O^ƍ�������<�\��=�K'��6[�_����������L�`t����f0�C��R�j�d��&E��c�o�D./��"=�hl�J��}U��(}��q�X8�xOc���!ٞ�>!M�J�h�N�(0G(�,$�񡬐�J�Z׍C�z|�Lѓ1�� �AY(�I�H�u�,q֥���B�X���m�bR/6�a��hm�k?��C��k�e��������^�7<t[?��uHorU��G�2�(s3D �3�rnpb�q:8ٖ��~wl}����5�c�
�����@�"KQ��P%�/O~��$Q/�w��<�y��tvǂ�=P�1��7Rk����z��Ɍ�"���C�ߙ����c�L5����=��O�*��̸oxH)/�
E���q��<�;���A^wQ^V0g��R&��@s(:{20G�xj��o�����=��yn��"��jO�a-X}12Y��L�K�����	1���c�j0#<Ʀ�LD�Į&�_*Ě;�zll������=%��iMf�a����w�s�6q�.�\��ԟ'���efG�H_�H�㖢x;�ĵlJ����J녲QG���i�4o�y���5Vg���O!_�Q�3V��T{fx� ?�ß���5�P��o�E��U)����-w W1��J�ŲQs˗9�uTU&u��<�(��z�`���7l��O���d��Z�xb*۴�{�{�)\��)�'[;���:�aB�Ui>�t��;�m��T�Ho�@g����)��$�x��ґ�e�u�=�&�����s�';r��y�AD'`�<d���EJB�;f=�H(��b�����K�$�"��D����vN/��XY����׋��8��C�f�˽%�#'�5lҨ'�m<���l�o2.�`e)SX/��R|͏���x�;�"Tẋ���0�N���֭���:��zFq ��]G���������w�Z�Ok|��W���an71������o�{Ug��
�}9"���!%��c��y��MᎵ���}�<�̍��(�sk�/�iAyv�Z�u��G*I�d�	��r�8W�.Pg�6`s�'�����:E�k�-"�r�[ ���s�����X9�S�����8�=��@:]�'�ZI(.�Pj����~����GDѮ��䑢A�h��4������z���F_�~��g�dsE�0G0x^�s)\�4����E��ѝ�����Uy�<Kv���y�D̋x;�!7[�^P�#���	k�4�d}��[݋�0�W޴��v��l}�\y�!�zA��x2�6��ƺ��%v�Q:[�=~� ���j�����T��y��5��~S�X�#t�����Vm�����K�&����������j7hp�+n��g�<�@�&���C�o	"�a���9Q�*�&+��,��8)��~`_k_m�Ȱ�΢�S��+�J���3� 2��J�m���h�}K�b]�Se`#�����Y˵��[�y�����?I
�`x�d��SQ3N�F�A��|S����ى����m�Zz�'<���BT��9ۿ�kc��;�*K�F�H,6!���/���9("��21������
o��E�~�f[1i�En�����aCD�!A��B�P�(�QTooRD��lT�^�}�
�|y{t�)�^E��8ޗ�f�#3LsĎD�Q�ݎl=u�1�l�ma��0MvY�$2�h]�O��a���Ǻ;�W�#��/�P�%{�����f��D�o��t_ $E�ě��"�$�o�W����Z#wҬ� i[ɞ�[�C�F�bu!C�/� "/FV_�)���P�9���y�l#�6�B��]g�p)����C�Z�\I[*�Eb=��}�6G��D�#ߚe���w5>��"2]��;��8��n$mɍ�ȩ]��Y���`���Yj�k� �ʔ�m�-E��Z�E0�ғ"�=[�?t��NA������a��U鈺�l�t_��k%�X@4A������Q �B����y�֓�Eg�U��go�e�}��-�����`��t��(s6ID�PF�ې�<�E�Q% %oDJ�C�_��j��Wp_��@��4y!�I<�/�<�k�-8�ҟH�m��Qfs�^�lYD��7L��@��]���rY%p����M$���1�m�P���T�^FX/�2�E��K�*ԗ����G|��v���Ԋu΢6�R��D��v(���G��R��FR0�9�%f]��5�.���靹���e��C���O��
z�㤠l�x��Z�Q�Ke�AE
W᎑��+.#-r}�Ґs�{n��g�~��ђ���%㇯����ﹿ�\}h�w"�J��Պw�SG��������Ӹv/��j�<\��k�!1�='t�����2ǻx�<<���?��p�O�E���t�(��M��?�&��Y�MG��&ǎڎ�!&	������G��È�-+-�o��.�o��ָ�YYI�]�Y7R��MN�:�_�1�tD���I��<��l���7��z�U���r�i�#j�l�buQ��*a� lo�5r�iQ���:�`��*��2�ʾ{�f�_�M	�݉}�LZ9-�m_���F��W����#��r��~{�N?�5�>8H7�7W}N�u�ٲ����N��ŁX�j��E�����+���c�:���� ��w����<_X%�����/��X�������= �v����z�,�� ���-��EB�����b;�D<R�Q"����]���x�҆�MT8&dT����&w���J�����D� �pn����%
��1@GR޼\����hG.���V`o�8n7� 
��7@NK&�ũ�3C�;����A�]��\ތ��k#�6��p�C��)=�)���
;ĳ��@�b�b�J��]��x��w�t��O�#�b���h�*܃��0�a��M9���,��?���Oq��zѦh��zn6،W��G�D;u�'�X�v���唂zD>��?!��m<��ؾ�m�~�Gj�[��W�R_�<���$b��s �NdJm�s�����e�"�ђ�D�U����[�Y� 6d+��a?� 
9O)=���&�U˚�lݎ�uHhd�?���"��Ȓ��9~*�=�8�͑�&�����H	�ž�B�V�]��S���s�Q�[����2^�٣]�k�19}r�����:r(e�^�W3@��Yӌ�L��Gz���T7P���5x���[,�`U%��*�As�u.[�v�z�˗-��:�Z}*�$cq�i��o{����SK���T}�I�ۦ��C�T޸1�� D�l�U���n��*&�������S�ۢ*����7������h��W�����)���HJ��i�5
}pT-���e3ƶ��I6���kp��
�[���؍���JuTY�O���	�[�>^�n�@sZ�����?O9�$�]/cZ;b�<]h�l��!d4@��{�����2~چy��8�����nha��YI_�c���Rh)�|r��ܐ����#���R���$�G���`W�v�y��eH,��ڲe�u遃H���6�'�0���5�J��!�8C�.��
��lC�9�0�	�}-��d#�Eٚ
:�x��(�~���S�ҌH�^q��Ą���p��c�����@��*֢�_GM�6���K���W"M�B	_I�İ��
u����*4��
v���PPXg�H�L�j/#g�s�Z���wD��|}1�AK,F+�#�JjĢq�m��
�������m�OG �\��,��RЃ^
NƟfD�Wz��^x�z!�U��;���r~�=����t�qҎ\�������U���+m��v)RZ��f��@��_��L�.�[G�aǅ��8�E��xV�"�V��U�$�"ϼv���p��!�_�q��x'#��E����\f'�_y�Opp�v!Z�GF����\T��[��v��O�v,�M]��zq��7��]�S���x�o2��i5���~�]�v�,�q��=�\@���x��<_���N�A�����R����p߶Szj��U��]�\ND߻�O��˟�W$45�.\��]���~�Tg��$6��,'�G�I�r��L�c�ωA�9�:G�C� ���3M,�0ݩ5H�ޤ��U�w��uE��|��vz��P�<�o�c���Tl)�Q~�l���ކ{�K�P�A������̃G�v��U���Ux�i#�el�Y��RQ$�%n��x�3�<����Uu�Y���+\\��R�/�Q���@�K�{��zZA�o�ޮ��f��2 7�`T��U��0\;��
-$���TH���]0���4#��B���?� &Ըq��]Y� b�Ĉ=X@����{�
3�u��4<�5�d���U5��`O�F�,<,�kTCS2*�Yf��b{0&��M�^'��.�@dg�WŽ����I��u��3V���۪j���N%F6���iʟW&Y��#��ۛ���ɼ�G�%�$Fv/@��lG"����K�#�B�ݗX��&�n�\DT���|�^(���yQ�3��V3���PQu!x�?���f3�A�z�w�&Uڒf�aѣ�.�V����ƕ��r�{I�qj,��~(B���0�Ryܦ4!Ʃy=G"YUH�[uƉAo���*ũ�I<�T�_�rـ�[���]=�V��V�����#�Wo���ǽz,�+=y�]uI���4Y��ǹ��o�'�-�kqA�$S�s�u7���D��O�X�c�B���ϭs�ղ)M��~���QBl�OꟌE�fC���,�VzcF�^� T"��v 9G]�6�}@�gVD5��U�.�9}Ű�F�
Ծh.�;��r���u�8m(����z��Ge�|���\d�D��r�	gۣ6��Q�b���H�����"+k~_"�l��Ȗ�әTH�(�c]�������0���[�g�x`�k��)8\5��C�t��*����ߍZ���\T�N�#L��I�o"w 5��>�D��|mr�K�S�������-h"���(�>�i>�d1�!���]6r�+�
���c��l�J���t�B���OX%�!$k��s�?���=]v^��a�ݔ36���.tw� �DH�Q ��U����C uM1x&��
r�M�\K�yj��u�N�ٺ�*�HU�L����r�8Q���\���b�3�?�v]���2�^���Ħ֮�ф���I����ee��벳K�dP��B/�!?]��&o򅎒i1��!�":��-QfH�b�֘Dċ5��f�����ش���^�����k�"��3��T�d�����~��(�Niag��� ��V6F쪮<
o��ȡyaO��XD؀?�FfDv��SB}��nL��#���D�q>����Bn�l5e�¡�D�c�҈�0�Er� %�������+}���fL�[*ۦ�};�:1�EB{�#j�&��ʑv�w���g���x�׋rĭ6��]� ��uNG.Æ*}7A�����s��}�LX���$�£ŋ���}B+y�.-d��T~��F��:�e`;�mV-�a©�F�J$�[����uK����m'D�ݧ{�a̭ƥQ՛s�N;B�3��j����2>���1 �Ͻtq�|�X|w�㟛�xr�TY�������|%��P lC��.3)$����^��Nb~�<�=*id�i�nd��UeKx>ԹI�t�"ד�rh���M�Z�]U�����U0�p�/[U�a��~�*S�G��.A��.���K$�X�|gD����k�R�)�&O[|q�w�kb1�in�r<L&���8E��G4�VkJ�&�^c�����m#�2M�Ew
C�*��+ݕ\����D��]K榋$^-5M�1�=��#���a1Dҍo^�cX�-�Co�!j�s���规��Gx���lI����)k/S��� W��{�E�*��h��~Dlo:��(�"M��h�������
m�`�I��RE�b�UuP�o����0�i(6��#'��5d�I݀�s?��W{U� ,�VU�|@�*����+�]����S�,����r��\ :GŐ�x\�^C�$c��j����W*�6i4\��{�����|M~v�*�G6"�K��cYˤ�ċI~��k���rrE��)��i��|�ZB֘:#�"�H�zMӐd�=7]`�P��K���D3��SV���7�&��S6s�Z�KG��h+���|�w�����f)_�s������I�����&����<2����׺z����؁H�qC80;����rF��L(�݌�6��r�e��^�z>���w�J��9���
:��p���dFBt,d�1��1#��,��i�g��md=��n�.G�7�{*��_~n��ly��c�A�&��z�/z�q�ŉ���9C#��g8\�5m?^�Iq0JC:P�@�mg=�Ƞz�Y/�3(C���A���+S"Y(�%d,XT� ��@���m���@y�E�F@iTz-f��`P�l*�r,( ]`=���
f���[Y���_�px���۾��Ȗ���t�	�Y7�%p���_t|>ޡ�!q@b[ k6�E�i��}��X@�5yhdBgȊ��:�tt�����]��`lN���/�
$�@M��d���=���KGZ�[�tX*���~�ʑ2S멜��O"bA?1F��N0H�������L(�H`�,�L'�Y>�H�r��:z)��� ��9R�eS �2Ћ�P�N`�^�7�Z �Ӟ�`��Џ28��~�o����xM IsA�
���z@e�ס�^�@���FA�^���6J��X�!%���]����r[��7�!!$ƜaL6~n����4۱4�����.�jP�{u�w+L\���E�Xyy��Ɵ���WCUg�{%��Zx-�J+��ZBs�O8��.�i�����?�eLǧ%'�^��bT���1�y��mF�4���]pu���FX,�~d`[X��`�F�f�ʂ1�,�Øq��.�>�X�V�_�Lj��}irh��!��>9Q�S{D��1=&%)�,S:5�q�ʑ�	{�>��n�6 �,f�- +e�΂l��lBg���j�ME��/�ě� �8���H�T ��R0#)���p�Mt�Ft�7��m�IFtp�2�����8�-�����T|A��4ͽg|�e�:�B-�4����t<0��H��?���':V|kdv�?���J�t�q��`7c�:;듟���� �ۓF�s��a�ǣ�FR)���-�n��h22�ĸ��P�s�m;M������ �m|�E0'_u���;��\T<Lw�������`�DEL(��f^�c\m���+� ��Oǀ�Mz�Vu,C@�;O�p��M ���`r���
~+�$�-��Z:�Rn�k0��3:eB8P8w�NS�gƅs�н���J�]�LHt4I6.���ӝ�|���h(:��h-��e�J�ke�o�ŧ+��
ş��`�Q�vC��@rAрQ��5 ���v��g2�0�p�s�av*H���OK-���`�!��Kx�w_�孍��k8��-�5h�`�c����44�g$������-&3
�f ��e�{���k�����i3_f��з"�C�|8�����į4`+A��v,�8��3�b�q ��'�0Gf���eƁ�ǟ6�x�8��	ֶ`��_��-��>n_7j3t$ �m5F���r.���΂?~�5�j��O�r��q�QT�����Qmw��	& ����/��5�3!���#��	G�m��杦�F�ݗ@z��{��Go�K�L�H��K���ß�- I�	R�$cC^V�$Y���?rC������޽�d޸����po��?2�[����r����PK   �<�X��НR5 �� /   images/52cc771c-8bcb-4758-820d-da79c3626c72.png�uT���>:��GApD�tH�CiP�D��;���i$����;��A�;�c��3|������οg���zY����{?���u_�u=C�e�����@��r�з AĨ���/�eo��[ί���|y�c \�u��v��~�~n4[�S�H�"��fo�7r2��pN+;��������E�(�$}��=ic�#$�؇��o?�W,i��O���I2�j��(2���qS�a2-�"ؘ�*���AS�I�ԋ�TV����/�����J�ߦ����� .�����������N����ÿ�/�׋�9��>�mP�t� b�������׏�4���+�$n��x��p�?w�ƃ��T����T����?S�oSY����&KV�M���"E�����b�����	������KJ�y0�p�_��3E�~�@Ҿ���@�g8,��?����������ۖ/SZ���+]be-�sQ��d"��AǑ�����f���\X�Mq����U� f ����h��h<�G���U�,l違��۫2\f(.'FK�npo�ד��!����z�@mU{,)����&�/IK��#`�z���Z��A�?.���c�KN�*��}������������_O���.n�sOX^Zm*s�uzc�N.��:)�5J���<Z�`�\���wR08�,�9��J=ux
�}�T��	�j��s�:$�!��u �Jl��)����u/����_ f�m�3�!�K����@����އf��S�ͪ��/�T��R�]�_yb��[��u�(Ij�CJ˭���]?]}�4��G�zE(���]Ә���4Q�,� �ި���'5T�iy����L2���jbeg�VC.�2z*C�����8�\��$q����o��T���a9����O&���
�jVk��4�����z��q�P�㽵�8�u�Uo?�*-�M5Lz=n�s��҄ bW:k~�D��Z\}L��nxm���Y>����g�h�:i��5��w/t��s�*����3V��ʖ(0&�����U�_�W�5T��TSv���w��ް:�xyS�ˡ��Gc[��6�&8:�`����ӧ�ri�����u/�Mz�+o~zj�vTM��9<����x�PG�!�A^!T�R�>&7��p�i0.A����i�����ш-J� !�9v\����� A���J�j���c�T���ݭ_-* qNXhI�r���R4�z �.&09��AA��m$o���ȅ(��d@Э9#O+�y�`	�%r��.���l���ӖǪ�|����R��lߑrա�T��ʁ��,�k(���$�٭���UOˑ���W.�ɻ��@���|���w�U)Rpt��}E9�d?aqi#�G�唻��^[��(�L�^J�/!A�G\!�:��v�FaR�ա���A�������7��1�؄�q���z���x�3P6�?A���]�|5WD����k4�0))�$%�- ��t�cI{��R|��h��/(��t{V���?1V���0�܌!�RȓyeK��yV�n�O��*��5M"<u?��2����i���b���X���#y܌+���b�5�1�&9��N�>���F6~=��,��"���sn9��$b�&�f�&��H����45�4Z#��2������/�w�{�/P�8<�Lz��4z��)�\.��={�˷ O�ӊY�M.aČ�x��n7᠍����)�^'��՗I�5o�x�5Gm�GYr���:�_�n���Mi-�q���V3i/`3��Vlڗj9=K���S�;h{p���L��k��&���D����;s�?F��~�+L�t�X���<�6b-�l��Q'���s�$���c�k�0L�x����x;�����yı����2d���2J�/�=/�=��0��773x���O���I�e �{�ol�L��9-��	�K�+���1��Q*)}��F�蚍M�5Ml�|����=k��������%�^>6^IU+�F7X��?�cޤ>4�Eb��(xT�@�tf����&VC��Ӝm|��sn���/��j�p���B.<�����ȥ��	��C��0d���]�{Ι2��ȳ#H�%�:B�E|��|����{>�ф�(�_na#������^��oܹ%�*.��oH�U�O̙B
l#H"�wb4)�4��b���a�����0�\��:��Ւ���W]�����3�L��P!Lr-�|�}gL��+�����h��V��PM�@3���=�tcCV�V�{�F��A_�Q@F�p���a-���Q��n�z�O���7ۂ:>R��K�8�O2S�lD���׺�ǻ��Kf1���k��Ή��݋��2�#��^����`�S�E16�����	���T	�h�#|� I^��:Q�zGG�IWV[�'а>�0d�fK<������3��,�݉3)raĹ~�>Nv޼��ո/7.3�ں�N��0�{�C�D>��E���or�DV3��1�'(ԾV�!�N5D���}rjƵN*r$��w|�3�>��P'�=p\Xb ���TR�<���~I�|�<�S5�&���oK |��̬��"�jk\�d7O"�Q�4����G�w+��7M� �$&�?��x-�FǺ���F=h	��lRN�����r�3�y_��Pƿ�������ܱzG�:��)Y�Ǔ[g��^#m:0t��Q��Eiح%E��T�������M�D� ��E��#A�U6��U�h�vP"%|�ߵUԎ�P�r��4P�O�������^*G��⎩9-�-�P䳛�~Uu����1t�A��y{���|�C+�[��(����7衳�Nr������"�wۏD��\��p���G�ʂT�,#\�[Q�$��h�
�����%P��f�_�P�J�������T>Ր86ϟ*� $�aR�Gr��mR�n��� �\���i��p��Lj�9US���i�4:�,?��6�����a������MWq�x`1�fJ�|�6����}Hd���s\_Gq�-6�	����L��3���4��ب1���(K�)�&_X��^��;Y��wI��6��ji��%Ƭa�∿�G0���"��R����g�ｅJ�E�	�y]��(-�I���h�`u�{���~x���F�������2�D`�D��^WߢJ}�Q�H���M����*�nN��[Q�0�c/���}��ߩ�p�-t-��jj�TԎ��2����n:# �?�%�6�_�|�h�~>�F���m�'&V�-3��N�Vư;a�n%\!"�H��7��Q);������S��S�����|��;>���Kt�	`3쎎N�Gx!@�Ky�&�m�d����������*�*���B��vh�h����o4%(�,/zRPжY'��=k����9*�3g���"��׻"��'�Q��0�? Kb�b�
8ZX�ƌ��(���G�2Ι<#�W��b*>g(p��z�c���A��O".�!F�)�@���5JJz^!Z� P��]\�;�!�f��NW ^�`=�X�Jg���K�U�ll���#l���\�x�URh�}�+ٸ�����֦���?���0�o�4[�qT����cM�!��7����|�,:��$���*�����(bt��R�w���+у�G����tn�.朏�mxۏ7k9���`t�Ph
@�go���Z���*��� \��N�,G���������g���]�0��+�������	okϳ�0<�op��Re[��d��~r�B�j��Y]ip)�r��-R�!�X��K�	:����m��Bj�,Y��r��=��������Oe�S���-�����Xs��U�w�^V��oRe����V)��)�O�vfa����¶��~�ʖ���2F4kEa2�ULD�)H�Gs�.#m��	�'|oQ�@O{�A����*�V�t=�+9��Q[�LM��n� ��K�n�۲6����. �<����y�w��l-j���Q0�^g{3Z|��A��E�*�3�< U�� ��R\�?����[�� �"�g>k����&�M z[��vp�䂤H:�nw�lOq[���\�g�������G����H�.
Y�C|��	�ު}�,�¶j��?jk��z��
����O)>�>�� <n;$H�,|��j5��z����k����0 ���l����CA��U�I�n�pw�Е���6�E\���s��[W����<?��=�7?���8V��u��zW���5�r���c&�q@���}����^�@z��ځ��)�m��V�S4|��ʲ¿�]�ud�E3��k;�R�;���j@�p��Wa�G@�\�1��aT4��hK'�zX_��-�a�#p�#�T���(�qWa�²i��uo^W\�Y�>�[��0����#��kp���~۷8��� p�H� ��}�SN��6_d(�����]���͐�Ҝ�}��y��
�]���5V�oܒ��Gn�_ɍa�!@��/F࿐Q�TQ5�H&�]�n�D�H Nj1bv�t�(�#�}���ΘIp���v<N8L2�\���Wd�-<?����yk&;����W�_S�;0}d�&�0���+|�N���޲���Gղ�
�ݣu�v�㵜���:��!@`�Ϡ�,x܌O���Eϖ��aKD)C PZt`+�w�2��y!m�g�g��C�ne��)?�A��H�>z-?������+����K�n�e���&��ȍ�-u�.a��kd�P8h��JC��;��J�n��l%ƶ%S���r�Z·�7���>����
����J�����gQpƘ��nK���i�^�;ޖ��̭&5B�Ϻ�7Aa0d��J�%a7����}�@��03Qw��ׇ���m��]��,`�8�7��/�Vns�	*.[�W�K������-ӏ���[�&5́*)�6Iq��k1G?�����Q?*5��'M��-�_�>�c�h	C��M��Q=�5?�*���1��I��}S^>�6�/�*�3��C��3����i�qFO8*��>_�p8��o0�����ƻ��R�/x�N+ɕ��ǚk�va���#�s$���6�?���x�p{��}��� 2���}2W��]z��q,`���x�����L͖���x`�L@�ğt
�"ị;H������kP:��C��b�x�8�h�lf��L��{��ǚ��=�?���O)1���bk��%��� ��> ��VZ��nO�h��ZT�2���s�]�\l��y��a��^R���7K�����F�;:��,���\�,��gyl ������ �&��#�E�{b�/q5�@I�e�"-���!iriJQao�T����[�Q���G���V�.R�G�r�����X+���
�(F����[�w!V�Ph$����e�+U��	�{�`+��r&	Y�P�/N�s
ν�����\��D5g��AM�"�$�����f�g5_��e��Cr��Y��&�Q�L��+y_���V�+a��'��BN����թ�<���_=#���2BWe!��.��r�k	d��߈2��frQ1��DB�O��+���3=��
��;�U�ȟ�k��f�s��IdF�U(��ڒ,��`�	��s��T;�
&d9B�"+���Y�O��9դ�-�:���y%���c�)��D�/!��z�^0��2��1Ƒ��<L�|��f��&�z��NF��Rzc�c��%����
��xջ����H`�6�x��CJ��Y>�aN�V �d��ҋ���2L��-2ڣ��Yk�o[r^G&��.������Ọ�����;�$�͋]�(J9*%�'��qҼl����hi����F ���Ҟ��D�k���V-󀓖��)`璈�Jqm돡��e��t����`w]�Ƚ����$K&ݒ�C�2: ď�[K��CDZ?��U�6�w4���m����֚�-���|D*�������G�0H`�|II'0�l~���2�+�2!�8A�14+�aY��<�;k@�R��L����_ :o_IB�������+|����~!)�,ٌ����a��y�����W�>�� �(���;��`g.�?'�3�GZ�k�O��9�P,Jw���v�fSO�cs9�O;e�V����?� �q��j<�a����U���Ռ�c�_vޖɳ9V��h�!P�dsE�"=r�z���l�a�ҳ؉BJj����R��f/��RtU�����zV��6�
K`&���>Z���sC8�H��ƒ� ���%F0�3��I?��{2�IC3��$>�t�������ߎB%�
�s��V���¨�U���n)	�Y�z����6/h�
����YC[�����������u6���Nb��Ĺ}��fPN����Ģ����K�֮��u�����Y2}ip�A��S�.cv5���a��������d�"~yo��^������N����Vr��D�F'���������t�5�c�%��rz��[��)�㚓Q�:�臼��I)��盄XO_H���۪���$�o�v��=�>����D3V�e���@�*{ai;��� @��H��f�zA����)����)��-�nQ��hH��tDKbDF.�>2Q�C��rU$�q��G����u�!M�_?Tt\Q�zFԞV���|���w9�n���;�A�J�nN{�0�"(@ b���K�9���o���������g���

"�ZI=Q�ɔ+y�#+@�D���gCJf�+��O^6�Zg��}w%�o*������(
��͎_X�_͙4���֢%��è����V�?93E��ӳj��Y�+o������w�Κ�K�"�Z�k!		%a�rk�z<ص��0�,���l��)�!Ҋ���+�8 ���� oO��m�!�#�9r��E���%�Er<�����Kw]�]����!['���b̏p�"�$W,��$����Y��=A������gg֟�'|��B+��%�({��׫%���`���犀���HdyN�]�xTJ\�J�8�Sav��v�@�K EM'���Z ������*���BƁ�ȷ����K�)�.�zVjj�o��KX�
dM���r=j�	����oڹŵ� 1p1d�t����v�����K�!�C���6�e����,3ӭ�;�o���6�����0!R����x�pX����KZ~-:��+���N��*��j�w��E�>q�,%�jw�T�(����9��J���6�1;u��٫:��:��@a ��֎0�&#Z�#�ֹ-�%�k{��ә���t����p��v4��g���_�e�+ ]�xXc�-t��rs_�i@�;��h�:_k*�۠[Z�uԱ��gl��d����R������k7��2�ohTf-�xD���ki�����l]���PY�`Uз�3����Z��~�ZG����V����ٗ���V5�ƶP#[O�q��o S�KP�f��L��A �~�k.:���y"]���2

X zuD�8��g��R��$�JZ�BfF�T�;����l-��`m�΂�9��&��F��	O}����|���Жm���^�F���C��B,��BY��u��s|wGL.��(E�m�
��XE���㩓�ψnR�m����)�:;޾jn�r�2@�lcG��߳�G�:�F�J-�:6x�/�p����m|��pXf��x�hb�đ�q##�uY�h�H�ӋګAbe3��h����1xw��bӞ����n ��Ӟ�؝\6�K|w���8�EEqq+���
l/C��lx �nߖ����ɨ9o��R����+��6�Q�-�H�o�
VMQ�&�:���k�p/JK���@m؊r=y�~�a��Ү�)1��QKC���h��?�F ���ϔ��	�LXA�8
 �K�)� J(��֠�/���H�\-�c�}.f�,�
�8���#]ӰV¾�[�E*2���?��4�j�)��&H�S$�6@=�X��0��-Z���}��rgE������d�����"��h����y��xQ%t��`�Q�v�(���m���+�Q __�N,}��ta=P6��$"���pC���}���-����F_&�(`0�g��.fE�����J|��Ք]�.�N;YW��O{��1��mL�_�Zwڔ ��׽.k�������/�����+q�mPC(+���^rHK���} �%)���Y�у~Z��l2tm|/!�B4�zA^9Y�LlP��<[���8�,7N�)+�a&�b��t���\�8�L���﬇����b7[g��N.�<��m��ϧ������υ�N-u��6��{���X3Z徤�����n���Bj����qt��E�l�]Q�.{.OjW����bC��Fp����VC���&��XX�ǩ�q�����%��~b��:��p@W�d�6�I�cR��Cb��W���Z	J��BHi�~l�v��Ka�}�JA��@Q�?p&`���͓��eR�>�D��1�0�V����PoH���F�r�@�B�l�x��`�^����"��٦2X������7c��$'�jA��g�i�#L٬ˉ΀3�MQ��!�՜@
�׏�$I}}G�H6e0����B	��s0x7���c��v?ĸw��D���{5K��hO��u,�nL���l����| ǧZ�Y���j�����ȸoݖ�hc�y-�e%��i��ޫ�˽픐��}�e&m��Y1!����4Tx��i�2�12Jut<���z�l5�6���,䆠���h�����;�T�*��xU\lw^)^_U_�P˲����/tc���އ}]�E�mm	�_(~��3�{�g�\��B��Ӓ;��j���Լ<&{	�"�0 �!�A?�7�x/>s�&Ch
��Rq���ZFA�H�7{'��X�E��h�Z�
��H�zZ0v�װ!7A����S�/����`��U^$��la�$Q�1y���g�Щ�M�1�>�������)�)-��$i��hBբ}%�n�~X.]���o����U!g�w5�$1\:ɳ����d��y�Ss
	�{���秬���w�L"a��˩����N��ƭq�����iO��w?C��Ro��9w����G�Bd�}`���O��ｍ&�� �f~��Q���O�=���K|����W�ܢ���+�+���n�/bCw*�:��_�FP�ǲ�����H:#�1����j�st����Nd�_�$�$�a�,@�ݽ�њ){�>OҽR5��mw��Q����Z2��2�B.����S�X�#y�r?>f��wj����|>��a���&P��@c$�Ux��`�|��{pM�`�i�eeA�Ƌ���*�	�15h9�0�&���w,��$�Qo4'�yYV/%`���N�d�2�u�f`�Ŷ��ö����I�s4yl'�CD�T�Q���1T�l�;�h ��?���E5IQ�6f�c"�n�w�i)�<�QKEm�xrE���2a�ecP�2��jX�ƽ1��=�9k�THJ��l�*�-�bX�Ҳ6 ��gA�����Y�m%�n�����0|��e��� �	2)�$jh��+��ɠ�l������Ѐ6���zV��
:��{&�;D7�AM)�E�:~A��>�z4�-�-ǸY�VTn<��ZrA�.��#r#ƴ!n� ~V�Л#_�_ޘ�r�!w�q���5|�\[�^�^؈�L�u�=��k�'�`��pe��
�[�X&����+��O{�я�}t��!1�=�}c�"�v�bln���3��j�a����`�˖/�?lt�'��'�a�N���a����~��:�)!�b�o{ϸ��`[5��<XQ}J��׈7��<�H�R,b�|x�R���p7ϴ���\z3�b�kʄh�3}�C��8�>J>4�#��������c�mO�UK�S��g��}�	�@���mȱ�QU��"w'�f9!�:AS�2:�qΡ�l+����Ǝ�f S��N'ZoЋ��·f��v�5^�Σ���L��R[�њTi��[R�v�b~�EW�K�g�����Y���ղȾE�׀��'�r�Vy���������"K���`I^w���'񄋦�5����S���B��n�T��B�m��.��虚��m=��:�E3�}���{���{m)u?�7A�.�p��o�n>i��OJ��M�L)�l��#;�2+(=-#{R�>҈t)�,��Co�A�֡SV{�"J��FP���*�jK)��hz���sH���2)��T�CX���W���k�ݻ����VR�;��N��m�����Z/s�A����*�#��w�İl�^pq�w>�!b���3�������6b3,q�2[}T�Z����nP4�?\A�����7{�h�Z��B�x�%���w*�K{�ߺL�t�Y h��d��u�7�q���fV��@�yG�\^o���=��3<��'�MQ�d&�C��໒˼sEy��d�j]('��_����Hc8b��ԥrzхפ^�ѣ��A��֊��c_��&eDR���A�N�.���ͥ �ZZS>	�)w��~��o�͐��c��ӵA�G��>���{���m|�c�`h����@�A�����!־��e�y!αH[��)q�����I7���D��;>	Mp������o#��LZ�j"&]v+��ѳ%��
S�&�
�`+h�(����/[����7��g�/d������uPt��V��Wb����W��;��jA?�>���a���&S�7�vaͣo33!}�B�˾���L>���2ϰC�'|@ �+N�(�Fy�V'�{�ٚ�I8�>Dk�.���JM�E'�����9�#~�ƶĦA�J�Ge-Й�.��ޯ���=����}�����]�E�N��`�X���U1��¤��Ԛ����F/nSe���i<����x���u�yDx͞��ή�wOJ���+
�c��ӓR����#h��\��uT�l�4�q�|l���~-���eh%%~�[փ��8Q��TUx���:�<�-��:c]v�����b&U�z������4�L�s�t�ߧ{�;9��x\�`H�̖�n��� 9�mYo�h-�=�~MfV���K�
���I�5��9ƦC�ώwhƿ��[-����h��b��o}���cؾ�+ezb:u����ϟi`��$�.�Eh�����PX㚌��q���x�����ՠ�9��PT��D5Dwլ���heJ1��$�%UR�ZK~�`����IG���U�[	��I��f	>V�?����Ͷ;l6�E��KpI�Y�o���5�p����ﲹ�30�1ש9s���*��n�׏��$U��gY����c��xc���5��e[�**i���[��k����-L��Bu�\T�:��Z�Q�xi9��Xd^@�s���N�,��5�I ��7O�̻_k1�н'4A	5q���q�8�vc]~�LT�@�p{��������I������/���L�kA��i9����l�V��t� $:�-��C���Υ��p}7A3��_=-=T<N�!���K�����]��y6�
׶u]�������F�)��z2���YZ�@�~f�L������P��B10�H��`w�K���v����	�)W͙�,R��>����Q�Eܩß�Od�o����E�����!=��X6�7P���&+W懗��%���n9z��V@~���:j�C��\j��Aְ��Xx�{���)�� ]��ȱX҄]$���Ɲ�(�(��5������M.�d�_C��� ���[e#�TDW�~�C�{��y&�(ө��Mr��#/��8u�g&9�8�?Xv����FIun����~�|�ψ~E���S��7��-��6K������ޅnwv4�I���ª{i%ֳL=��)%j���^z����Y�t�͞A U3���k�p�?p/�����٠7��j�)|[	>]�DD�tx�;��/L� u��W��oݞ����(*(xKBx�-PF�}d�uC����@^s��1]��EH�5��_���mQ��,���z��X�Y��M����?��_��Jߒm�C}{�=O�e򾥽@qL�-6�6.QO0-[�,[i�7���Il�TM9=��3:`�.I��6,���nҞf�F_p>�̆��Ӈ��[Uf�=�cEڞ]��m�/q�=�R�Q�]��`[���׆�*���.~xK�2�ga�x�U0F�a��r��h����a�<:[l�Q��c&?��)�>��0�cj�h|Q�FM8���y��OPFu�O�4l.�Y
mU�ۏm�N�)�I��I��>�|ϫ �wR�D���P��<]G�	O9�OΚVEi̞-���9?��&��X�R��b�D���g�ު\�/aX�7�X)�.��'�?�Zk-�\+(I�|����\f&��w`$�~%/���R���%����c����(�ĳ�r�1s�	�΍~�!Vӌ�q��S��9Ǆ���:0yq��M���
�`"j;m�O���_.�<�pX�ѳW	�:�h�����-rd��N9%�'hD��b����:��n}A��(e"�N>>z&k���ϊ�"&o9�9�\����%k� �S��^T&��P�����X=U[��Ng�@�OFs�=�Kt3�i�B�e2NH��[*�׏w�sD?��Z:z_�5�-�n��%�{jZaC���Vybt"]|�����*ذ�"���9���q~�^!A��NcX�żW���!�e��4v�Y�/�K�H�א���¸w�����m�l7����į�/z�*!��J�8N�35��ŧ;�\�S#n�V@/��$���!N"|^T&G�|R�u����q�$����A�V��Dǈ��V�c`7n�[��P�΀�xe2�;}��(�ֿ�����h��W� �=_��ӄ��xF��"_ګ^�%Bx��M�0=a���Q�lNE&����H�᭦ᕑ��_��Dn��~�����[s9��K�l�����Z^��q�D%f���%�e�[��>�I�_��\yǿ/���=1��cb�Xm�,�_5����3uP���7�83�uTK*}d�W��/p|�6��/y�˳'�Ю����gO�m�q�����~VA�Z�ݦ�񑑍��2b��@_����a�r+CZm�s�U�Ã�є���6����������zk}!���2>���ӀUN�^�͙ݼ6uk������B��Qr�SK��Z�l5���l8kV;�p3۠�ؚY���.��@��;_��x������ET�+_�F��&^�.E�6SEK����3�#�i<���o�&�	L|��2W3�1�_D{˰/�{C�s�B��[����p���<�=I̛��e|̭a�[ڽ�!��ȷ�b���;�a���[��?��,@���;�kI�,%)��W�9~��i�_�
Y�L�885K��ي#|a�0�
���%Co[ �j;�L�:J�$��mX���Q8���ʟ����[��P���u��1�Y �rc��d�}mP2G�7���3)���CM�~J6uc#]���	d��@�5��8
@A-e��z9�s���?�)O�X��zut�)3<�i�Ŝ��Ηa�3���٘V'=�o~�SL���y��[U����{fc|�jMxmD���~�I"1�$_�S{Nd�R��ۮ7��8؟��2:Ͻ���@g���Չ�G-6!&F�J��y�@nA�:�)�<V>o��*u�Ҝ��B�]c�nA��˞.~���	�jDH1F*h�����jv�]�YZ<ғⴷ�\��u�;v��ļ�&���Rm�V̯gdĠP/��[L�sW{�Z/�*3g�W��`����V"ƞ^�K旲������F��l�IMPJ�w��̈́���W|g~����N�(�cB�me�| ��vpDqn+��=���C���$S���r�}��ֆ�c�J� !Ը"����ک������$$!>��@�SJ�c��ң�d<��ĥpL��m�Sk`�Z�:��J�k���n�]P��������*����lั5Vn\�q�^�Z~d����8A;�Ŷ��ix��{biGk�Ab���,x>&f��4�Y*RՅ����x������J�Ŷ��9��Q��=� Џ���tM�����wA~7�1�����o/�1Y����I=��:��v�O�$F�\xˋ���͘zn����Ъ�d���{�|���5�⧹^�R�x$��p��m��K>�\y�x&IW�	JV�������6�u}�VpÅ��"W�����!s�_�1�C�0�!R��k�r
cU�ϒU,q��Sѱ����~����|�����dR��^�۵�K�oUaK=Ht����}�$��w6�@q��Ux'>ƽ��q¬�ӽ�"oBdG��F[��c��������0)(�K,D��{�ǰ�^�u������b��s��(�M�G�d�\����M֝�<&�F9����wd����^�ϸ`$S�8�ҦU�I�N���^�H�`�O�R���;2g}1���}��|�w�m���*e�(���A�/ \2��_cD��$+|�o�d	�Э���@ ���t\{ ��-`	 ��;8bMQ�[ۀ�z���)�w��V���|��}|u����8^�eJ�y��ܟw��u����v��yY���*
�8%n�s�|_{���U��`TD�pZUQU��VD����wZ�k�9*����ހ8i���K+s^��"�A�� 0�
,9�5�����`c���a��/�<i3^!{(�v��6�G�}��c��n,��R��B��;�Ѭl8DQo}�YAjC@��m�6t,e�f����5��V��eM�D��^�^���E?z�g	�@z��6*_���\)s�^K�*�z��?�6�+a��
8�>��;]�������(�4�i�@b��]�䷖x�-?ޡ���<}<���2jab�Q������� �J&@x�lGz�`S�Z?��I�3^2��:���U��F�?jE�lz�^j����ѭ��Ќ� ��2��,k~5>^�,7��� �Z��aG��"AV�Ӊ��|�pE���,�u�]�
? �k��?: �36^1ɽ?�)w�g3$-����]hHR����#;�_> �xx Jg�+.�zn�s�ӎa7��0D�|�� �`��.�a (�  9=Z<Ā�l!�H�S�WwF����a�t|�Ы�z;5��+��-oqCo3EϹ�Bo�6��T�vD�(Tzųɖvx*�<E-�^�S�tor�\�[h%�!m�"���u��y�� �l�-ڭ��ҵ�M�W�g�#@��ֺG|NY |N�N����9t�.\֝�Rt8!�A����7x��#���Y�R�~!_�C�1U]�	P����Z%�!D�[Cɶ~�|t���&�b����X�j��&��	���V��eVS��6}ha��۱@�D0�ݑi 4ʟE1[���Jԙ\�|���$zۯ��筣u`^�ya4���Ʈ��c��h}���p���m���̘�L�nh�_��"|$5z���������������󵹕�1�@�u�L���@`D +7iՖ=����T7|f��`��ęj/��t-7��<�/��m<�3�y���@b���DO~{���g�M��ͮ�L���Qk�J^=�U&�}:2�k�dp���`��8��-�KJ?djc�����m3G7����@.�_�X9d�č�q�l��j��23�"���zc8���y�(��o�� j~�!�ɧ&�j	����5�7�/j{G)�׹�\/wZ���g񯬶
�V,�z�F
�*u�͒�m��/�ت\ y��0�M���j�b~9�2@b���F���� n�04K�u�#�Uo" �F*����UMe��� q.B�C�m�:Cx3��@��[/��,Z��ٟ� ��F�I�� � YyJ$�"`�
Ck2^�(#]]_R��O�p5̛V%D:S�����X�-�c93>W�-,3�;FZ�1��{5YLI:�!� �r����
:MѱÕ�.?D6v��13<�ù HgPFk�}
4�o�	1PW����ǹ��8�'�vd�]&5�4�=~�c�W�"$���&h�����+��+[�Cv���l�t��нXW�ֽϖ�}�j��`3��+�/E��=������P�B��~:�>�Ѽ�{��-���N]���x�0��	�� ?>A&��m��Vk7�(���S��
����j����>v��0��X�$����qU�w�^��?#l��Wn�� Pm@�ۺ��H�%$}���z�tȂ 1ڱY�}l���s��22T�����5�� hô�V�K?n��k9���\����b{9�=��L�X1`����>pe�&��@_O�),e�qw�k�ҸO�Ⓖ�v�57�����]#�Z���9<>9yz��#�O!����j�+�K7�����o��hz����6Igz���Ԕ%�mp�g��Sj t���� �o���5�m;�:}�V)��j�����n0W��t�!�Ȫ���l�z-��y��U��$��`� ��{Pm���[=����*�RF��Z��$��b�Tb����q
�4��Ry�^��&J>�q�7z���/@48B��8����O �(�@0�����Ҳs^KG/ 2�q9��2k\����Ŕ�[~�ó�%	*�s�r�{�u��ά�hMb�a�҉h١�k�-���J��ȟV�ٟ� ,k��&�G�����&�6}C�}fo�0��5�#s�i/�G�����2�f��դ�w�^�O�#xmx�ƛ-|]S�ұ��@�C+��uq��p��PJ3f3�ڎq=V$�Pimf����g7�
�Hm�$)ۗ�T�j#yߒ�����$�/�{U]������M��6�����x@,��ߟ䑨��c�	ڿ����"�[����ﮕ�l~�����:p�G���R�
��E������.�#�b��ꯨkС��@U���b���L҅`p.l���;�<�Q��"�nx3#�kKq���#�C'��7�[�z�s���?�W��Srh��a�GAf�����j����QD% ���Hu	)�%��ӤA�CE������a萘�c`��ټ���g�zV��׳eb�'�#��C�V���%ti�c"8l�w�Us�\)T�W�Lj�e@��8l5�z�>:�O�IP�e5@6֙�ww���$�U������L�C�|x�Đ����q;�E� �B{�O�~-,�g�s����|/e"�S��1B����*eLvD�a���9�4i6�Cʤ�/�j�@vpz>RIa�ޖ���0���.��/���O2|Y�c���B^�w�7{����A_L�"���L��&m������ZMa���	�J�Pb�!���um?R��o�.�����o��9�&��;���Zk�3��g��C֜j��"��@w���b��p�"�*�ST�O��],#��җ��ZI<Ix5��١���7��8w���O�ki�x�!�1K����`G��!	���S�#7>����妢�w��d� pl�����q�HzS�����qdk��=<E/��עBg��S�k��:�dk	����'Q|�Ou:�{���ݑ��˳1:�#Mx�0�����󹤭��s]$ޯ��-����bI�ϗ*Bax��IKBP�P��w��7!�2�s���ե��ѷ��_&��T�v��ՍC����7��"$�g�QW N�ON#|)۠x^���9L@����ό�9��>=�~���"�&2j�E��͗c��=;G� }䫩��:H�u�M��������w�:����9�G�DŴ�zS��M��8 �
d�
�W�� ���L�u��p2��8k�V�Ua���� E��o��������]-/(_ �;*f�:�x���$1����>E��J���D*�C�4��� *�_(�a.ں	�_��<2=/�4Ȕнt7'���q+���R��T�L��+��>�f���K@WS}+&�,���r'�Ջ.�ڭ-j���対]�x \�M��om��/�?tD��Ҵ�a�T2������G��F�����aC��������9�������<�����|��C������~�WW�*���63���W��jFR���T�[!�}��0�`� ����p���=�W:�M�j��V�J))>�x�s�������ѕ����8)/H�� Kc�����ξH������bR���#.Gui����x��"�/��)�����q����U��6���]XFo���CP���f"��~��=���щ��e�so�"J= )�Yq��n�'&��C��������/U�8�������ѷM����]��b;y��K{���D�4�l1��z�5U@â?>�t�$�!�Z"��毖��u�s�o�Ju!� `\.��X3@��e'y�姀�6�C�@���\��kL���ր̃V��].&���d��{��kꘗ��1<11Jk@3��|�ƌXK�%̊ڪ�.ꈺV��>'�eFn��=���$A���T��c�:㰜���=�֭Qp��i'C����l�]BRcQ6
��v�J&��k�YΛ�������!	|�@�9��X��4Kį���@�����s�����- �d��d(�0\ȕ}bc3�+��z{/��#���.�o_�:_a6H�WY1���"V�����$��gD�g�pݥ��O��`��6?��$hթ���w��Ϫ'$ߡë��q.=���Y�k��l�g.RG^�EN��n;䀍W�K$�(�IUg)}"�'@5Aq"ȍi�ٴ4�bU�X��������E,�F��j��,���J�}q��gM:�Q���U�_��;�h��pՂ�r��~��;�t�I��J��z����x@,�Xsn�I�0G�7�1!�H�]�%z#��
2e�!Y�W�Y,$Iy����7.��Pb�R��Fmjq�UۺmVmH��t��k4����6�� [�0~��][�758x+^���U�9_H,�;5'E]w��㙘�p��ԇ���ۍs�� ��n����5��N�J���ԟ���7M�u����z���~\@�+��')�^��^�/��P�6��J$a/��ҺGآ�c`�a�6���#�m�E���k�_g���u��=;��~7�#�
�b ��JR{;nNf6
L"&u��@H�E��`���
/qHLQ�
3iZ�C��P9�\J��d�vK�GE�oes�k�Ĝ��NGωB�D�נl.d�=�����?�e�����= �^���O�V�d�7�:�I���oU�|eo�̮4�\��|�U�w��'���_4u��ؓO��E�;=��~M	q RA���?�'=�!���`�S��wR��bM���\F�G%���X�yxYp��Ӓ�I�xU�Z
�\^����Z��Q�5���'8��hh�����J��0�^oڲ��$�y����hrK����^���e��ྮ���M	t��.�PA�RjY�[/�־�̜.���;H4-g)�`v�b��YP���L0�����ĳ�[���&,��1s_��]��Uo�s�@ۦ�f
�ߩ�g� jQ,����j����Jsԕr�7��< �1�����4�(�.�Z������lj	=���\X�[]�)��T^�H�L'c�?�|6Il+c�`(��x`ò�����	�����F|J跐��p�j��x��A%<_�e���CE����;)`Pv���#4PZ��������c5��y�V4R"����Iq��饎���#������;V� �0��!u�^`E�r|*M�moc}�ը5�?@���g����'V��� �ʽ�mm�E6fe�r�S ��2-�d�oަD�.�6�~�R0�,�F�
��eq�0IK�b���V�������y��:�p���3��|�Q
`���c��6]�t�k�W�\�W%��A����B�3�+{r�E傧�������P���o\ QD^��3ɭ��ݘe��9 �(VOH�vބ�l�J'�6��������Q�Qs}�R �c|��6ю���N#�U�>�V���P���k�G�r�◻���K�M��`����ڳ#� ����mx=��sQ�j���?΄�7��hu�.�A&Z�=�K�j;73&N�T*�:�4{�̖�~;�_Bq������ò��a*��審X�DA��N��Ԃp�G��8���@���fX	�f)���!�3��p:��9��[,��!�JW��xpq����ǉ2�ne��an����1�>Y�ܓ~k_�ɹ�C�D�@o����*��.�5ww�q��
CZS�i݋������l��'�PP�1�i]l�C/T��.0�4a��"��>E�Җvs�ƺ�|���_}S�3���X�݁7���Z���x����֩�dU;n(����%�<�p�T!>y��f*<�gO�О��3ßkMz�;:A���{�ۓ��{^NuF3��gluN�%_�e��F���߆�W<������v��1�M�1�>��k�ts1�3U�M����ZP)X���,�:`y��i�����U�q�U�M��a�����4��G��J���ӌW��]��y� �.o���m6�D�G��"�n�^mX|�_�Z�5�x�ރ)���w �[��5��~�rs<K� �����}ÏzZ�΋�Ğ���kkd4���*~��?�[��9%��j��������5�٪RK F3g�B;�p������.WRj١�JNƨwŗ<6Y�IS�{�D��J	{�A�����/ډoW�hbc�O���Ԫ���ݦ�;jRJ�� �Ei����5�]��!�{�s�ݚ��
a��W�,~��6��ԇ_�l�?��_2-��pou� ͼ�.����W�R?�v�gw�~&�&�}<���:��#�p(��\*�!`ۊ��c;�c�\�6"�-^��`���}e/��`��s+�-���O���ձ��`�~����;ѕ�/�5�@�s�Z��q�8y����<`�G���b!��'n�MB�w�ٺ�q��^!�ZS*ɋ�����f�J���Y:��w�&Y�Ք���>�p:�|���Iמ�5����m{����H�t���a59�.(,���|p��7	�F��$�%L*�xw?�x�0��V�B,qݺ��BIJ��#�:I<�xi���M�pR�v�������Z��3�Pn��m�rlt���6�'�|����TAv�܇J3�W]f&?<���틧������y�Mhz�O�P�궡��gW�����5��3���@±��A���o6�6��)�H^�t��m�v�Mk�4�W	��U�qDJ��TE��k^�m����d@��*�RMS�t�|�C��!
,5���� �"����uPt�/?�"�;�G*'^&�X?���Uv���n��J�9 �W�dui��Ο����o�7$M��Y�ʤ���j����{9 ��*�܍�uYA��}��f�e>��g{�A���,�L�AR��z4)6p��W��_@g���u&�]p8$�|K�c1~�#���&"�؀p���J�,��nQa�Z,��~�:gZR���|�~5Y�c֥�[�"L ����fpRyW�l1�a�0�,ITB�]`��1�|���e�y>��d���qw\{�F�?��]u�s2t+�����AQ������j�C����O�����M�7f_�Cfa��d��M��E�%l�-����(���{���Д�~($R� �|/޹ы7d�	<�:�~p�~��e�>{4�ָ]=	���0�`�p/�k``i��w�Vd{w�쎨5!�7�q�4�W����$�]��p��Iv�&��0,#f��0���\�!W�q�O�_ϳ�%��>� �xP�����,e3x�Y���~�JQ��5?]u�B�c9�5�������W��))�J�qڹ�?X4�gX��F�Mk;K�U���?[�+D�o�R�jZ��Y���+�����������BJ#�'\SS.+��ύ�4i,��b�\�B�$'	f���5^�p�H�[6��#q��i@�h�݉`���;�N�U�h��%����'��S��k�'I�ѹ#�����9E��zT�E�u��1U�L���v哅k�
�$޲���қ�)<�b������ScR��q�W<�
��|���$�������vGJ��/�lU`�<o��
 �l��ζ���']���hh+.�'��Fm��&Ɣ
���ʟ��L!hZub������v�K���f�'QAb����5��7Ԝ@�?b��+��?�_~����F�AZa���b|������:I�9e������曏��0q�ߤLy�P����YT��a�Y>qeZ*�=�I��Ƞ9������Q�@�.�2�Q4}Dt*�����zc��j��X�@j?m.ȏ�)���E��"c ݦ����'�P
 �J)nD��a�'��L&;����j��m��p����T��<JtI�}_QU���l�0�}D� ��!��>�� zܴ���hX&��i����v)�rן�V@��t�|n5��vk6�M���]���אں\"����˚�"Lݍ�L0m���������=/E�\�ܖ?�3�?w�:���%}�5�R�L�oR!�3��<X�����a8�5�=���q�����Xm���(<h9ͤm���d��''u�
?Zw�
D����n��j����-�� ��}i� �u*ӵ�����<���;�a+ҋ���昴�	 �D@仓ؙ?�F�#��7Mq<N��Н*����y�+��R��X�Qv��c��R���k9�`/�G
�G6�D�2"�NZ��D�D�5T%�6��қ��A��x��x��vv��p���"7�
��{I���g��vo�q+�6/���T���Fs{�;VG� ���v��ݿ(��,`U[�a¿j!��X�y��$aݼqCej������������������eq�᧸����R�>�$.�&$Sw!�W���v���]�g:W9��]�;6{�Y5��������c����Cfk���Q���ɜ4�VKX h���F���3LT�d+̼���u��O:�~<�[�\d*ڹlRؘ'N�$��j�xv��r<��.�x��W�W�+o�2~6�U�"�Q���@��V�-:��-P
�ծ�����w!�{�=��ߢ +���	a�y���.�u� Nn���`�CQ2�@�����PR�=��h�u��oq���=�·��}�ڌ*����.�8�3'�Us ?1}]%ַ�UD���&	�������Z�7����0�Y��p���.�� ��$�v�zZ�3K�	�4�q�vF͘�R)���6����t���A����D �����m�^Q9x��Zr��<$���.�m�{�hbw�f|Fi'8k��l�7�����T��HZD2�v�y���K���a�D'�O�}+�d-e��N55πO^�T�9�.�u��C��Ȓ(6{��ߖr��y����X*(���o�ʣ&��`���hK�A�a8�����9ňC%�Y�#�%~��,^����H�K���󂖕���=U�2�����f�&;o\O)�
\��V�����l�Rm�D��i*����_�dn�O/M�NHDy�ރ�g�ʪ_1��~�{ŗ���D�,<���ހp7�~������b�ѥ&ƿ:�^K�;��;I���GL�)���;��l2 �>h	��^<�_�Ǌ?��<�nv?8�h�	 ��)�ܳ;I���t�Ip8��n2��l��K5��c�M��l��r:��$�����/<:lͩ��:��3?���	�+�1I#�q�+OZyh,���|�2*f��B4&S����U+A3�������#&��K��!I;-2��Xk/Y�?��,,c<~��P��N�����g�Jߋ�W�� _�۪����0�^���������s{2ԉ�6��Yx�B���u�3������U�>��")^����߻P6v�w�(�gq�����;٢閖�+U�g��0�6�`%n�b��� �BS�pIд/T��	0��q�Eq,O�6�P�����2��Ŷ�4�ڸ���F��o
?�xgąT���jT�l7���M�8|hZ��cw�
nw�$ou6�w����>΋ �g!���?uU�&k�f�6Z��n-�s_�MOƃ��_Q}���Ԇ_q�2���M���c0KT/t���9�J����ܨ� n�� Wqt�$C�Ѻ��@�ä�T��ەRf	�����R�����Ei=����䡥�Kx[Q면Y`�쨬"��*L|k۔��N��۹p�}̬^�$5�1��}`��>��5u���K�`�j�+���;���S��} ��N�V5�]���7F%jNX&��Ǟx�����.�v���lX�c���:=���J�ܧ����4A7��S�*"��YHd� /�j@9��Ϧ~g�M��2�j���Ϯ�Z�\��ܚ�\�Aq��bP*A��n�e���$�mQ���߱^N����JR}\Ld	"�-�yr���,�+5c����ch�~�@ �n�'����o!s���v�����ȯd_���������na��� #��;M��;����o>����e^��sd�A�Ұ�!�|�o�_���Tßr�7��Mʝ��
KgJo#A����}}3v�u�OF�J7�����M���� ��`�ΩR@⹧��e�b��^��F?��jL�7��D��S?B�m��Vq|�K_L=������`Y�x����2r�q�l�:��-<d3�Ld��J���o?0�5I��	~�o)����YfL���.A8��(�w��s�x`��nmx�����x�����{��m�k�K�L�1���խ�f��M���ժ���H�*�ݩ���uV��8:��F�!�Ӭ<)*���K���4n��o@{��dԎ���I�3��|-[?��� �����Oٚ���^�>b;�c`j�yW�!߭#�aL��i˔�k��jW'v���S�X�B��SP��"�ͳ]��y*�p��Yڐeè���
�AfN���
�����[�>tZP���~W���i�
~��~�4�CG�����N�ܸ��mg`����>y8v��K%{S��ik��$p��%��W�5����������A�d�LĚX�y�g�?܋�������c���c:'�a;�6]�(ŗd�?�L+�&����^�����8?���=�W��zyJ����T�w���k���P0a-{-�Vm����hU�Um�ohjqF� �Y{�Y���y(����0Nۦ��Oϼq|���+ǥ�O���o�UӔ�8�J�����"�'��8����� �����;θ˃Ѳ���]E�}���#g����&*I��7�a�	%���c?��/����S.گ^L�hę"YhY�oܔ�2����g�F��0L�LX���ag���������t�Q��t�f�m;�j�˷W�x`�W��P4"oc����~��CT'-M�`Y�Ф���7�O�ߝzA��i�����!|�����'?v�lؙ��dr�D�"���t
�;G��QċW��Q�s���_M1�x�P�ӿ�S?��b�x��z�qzm�ӣ�PfR�J��$�a����~S��E��L�Z��M���n�E�s���l�G5���)����DuHm�J@B����:N^�Pޘ"���>8f	�F�������oM��\c��	�.�Ac�f��G��m�l�吤H���X����ܼkpU'��1����ze&��{
�����w�@�/��wa��t�`��>+����Z'���`U��m����f/���D�u�"�Z��s�*p~�ϱ��/"Y���ސi���u�
A�-��u��;�'����ad��˯>��P�!���J�}ۀ��$Y_�m��k6)�-�Aua,5=26�*��A�����ĥ���>�a��Ǎ��E�+�u��l6�M���i� c#�F
:iI������Ք���hzN ��1	���9��!"���2�_�����H�c`�iM0{�7��Ja����?s��+M�m��@�S���vߘb��)��	Aggt. 5�WX�@?Y7�~��KH,�zd*KZ|�x��|O��p������cM%7sN�)��9�sϗaA�K���)��y���7�H��%9e�e�	�lL�ǳ��S�F��sළ��h}���k �ܹ���_�^�+�e@)�(K�8�1�������^\�]��U�m���F�w�d�|B��M�0��D�����(}c$11%^Y����WWc��a\֡��RҽM�J�!�m'����{��Q2�XWW���`���ف[���ON�Z'�8�*W5�L0�d���tq>���o@�@��fff�I��p���!o�3�
*ۍ��)A}X���b����,_���~Cݛ����ܤ�r��/�o�@j5���lJ,���zG�n����.T���r����0�G���F�Lmޜ���f'�u�u?<�h[L�O��8
����\{�p�t50��K/�w��D��� L�'�OA�� \��o�6�'�#��ͽ�P^��]����ng����U�r�z�c@������`�O��j
�`�?_RW�ʼ#���5z��y ��H�O�$����b��_D+'_��	����)	'@0�IAh%����B!���� �7�$R��rԕ
*Pob�ݡR�� �|�fl�=�.(��x��r�C�d]�0:a�::��/���i��H�is��s#'�AM�E�Ӛ?����4e���[���HF��#C���
�s���A񤈏^ϲ;�u��̊���t��6�~T�
W}��	�O�N����M�s�6e�R�1Px��
�x	��a��$�x"��e� @#Y�*(N�昷iZP���l��v�u�[���ȖN�Z�'�ꕼ�xd_���n�;	���uQ	L�Qd���^����nu��W.�*7�w���S��Z��Nw�qA�e��q����R�d�w�OJ�;�Q� � �{��ii�
2!�Z�%�az!X��KH���a�~l��+T�׻�_��G`�#�4�"H'1��S�;Q_):Si�u��V��c�NY:g��\̫��ܰt�k���ݔ#0��@7�o]�ى�s��b���U�Wy^�|��mN�����;��o���Wk<���@w��/(ߛO"�W[���,��$��񱉣��	@}�-H���O��u}Z�"0�+[��v��m���1}�Z_ҁ���w(:ƈ�4�G��eGx�.1X�p�a��c96՞��[���Q�U��׬\Xu��H��>����J�P������gҠǘ� 6x�Q�j���=Kpz�����@�bY��'@���++�N�`��b}T�� �_S])�<��7���$@�d��޸g��}���q�I��JQ@���_�hm�f8 ����)������p��8����*G}l*^o��g[���0���\�6����j�A~�S�DmFQ#W��P���r{s0��%�������h�ԶiXD�-ۘ��ٟ� �� ���'&E]2I?���Z�fF�T%Gٹ�{�[��r�r�%��Bn�#�u�[�A���Eg�۴�Y�{�4l��X�]��~Զ�W<��bj���V��˯��!����<�\�['}S2�q��d�� 	�����DW7n��p1ֳ��80lCC�>����	��Y��X�/"V ĿuV��_Ⱦ6C��Y�4�}މK��՛���I����̡�ܠ�xL^g*�x��叔!�WRNۿ�h��By�T[�s�B:�t �������?���5^Y�)�c>��fi{X'��ҋ�=m�DӖ��;GưT���3�0UW���q���h���:�}�tr���L:@&�S��� 4@g(]�E��'��r���.�)ծ}�sJ+}: GPVnQ�v�$���I������!�ޝ���qȝ����r��ގ����µ�Zm|�a��9��f#k��5���rW�lu�<^w��h�j�U6&��2�%�<�����椖�>��8�Z�7�N6��6zX��_����$�'W�9����!h�9=�0_���|ܰdh�ȫ��Zk��죬��d^�\�|�m�`�O�Z\����<��v9?Lr;��_��E]�M��U���}�;U�>�Lpn2$��~Vnh�`b������/�2��� =W��!粦f/��$�����u石|nwVƛ�=C&L��^��₅�x�-4���뿄gz�u��m���v^�Z�4��)+�����Uv�}v�l���֣��T�9��&R-]$'m{�0��mW�Y&0��QB5Y���C�^Ub�.���d&�Vg�tE&!Ӊ�L1�
ۣn��H����N�[�D��>){��+Ob|Kv�Vu_{<����S�a��M�������Ґ��qe��OV�u@�<���2�r6e�x;p��˳s>�h����8|�f��Y3�r1*Mr?k]�dZ0b��@,�^*[����[�(!�^��>N����:fH�H�����$��iK�>�"꣥ �g�p���٣3���5K<\la���!2�x��l�4~@Ur�]T6����F�����&(�|/�r;QA9{ 
�:G³��lT�u��%��Z^�S�i���ai��&�2A�~@_��A1gKd��6�[���/�m��>�L]�/�ds�փW�vS�QC[��L)��p��	$�$�P|nH��4�H+AGX᳒Z������L�S�����褣�>���N�ቼ���n��L�W�O(��Lu@��6���䗙bZ�њ������ϥ:~Ya��E����˃.ee2����}����K��2��yJ�m�:	>�_���7�<=z����zz�Đ�K�V�j����ۻ:t�Y���zT������fg�-���:@!]����)A�����k�1E�"˕^e��ύN�Z����g�x����t�h�]t��&r*YcK��`b���m��saIA����8��%X�GDk4���I T����>���J=#��}9�_�/3�Yhx-�Z�WL8t�,?�[\�:�Ջ�m��-W�e5n��z����j���3���堞��[T��r)j�d����Az={]5C7u�»O%KS2!�S�����48�p�c�M�ǳ��
m�hM���eR&ݸ�I3$��!���w&�#�?T05-h�ط�Hg0G�,����E<�^�"�l�}Wx`��J�I�Sɡ$*T`��/��}K0���j�`߮�J�q��?l�I��,y����v���[y�����S����rj!jA:Q�S���Lf&�o	<�c�7�!�y�+����6-�	���oۍ+,=Y��Ҳ����ziU� �Ʌ}A�H'5��~1�^�"� 
{���^=�0�n6ڷ+vs������s�+�g���1��K@�'���l.������8: N����ESQ�[�
�:N&$���e�s9�o��`� ˄��a����P������e�MN��UK�ȩN""`i��(�,��@�Ȫsn�x�Rʄ�{ҿ�5�6��R��:����䀠W���l>��x�B�ۛ�Eݦ�=p�5~�&j(��o?���B�962��Hq��ۊ�G�K�7\�o�����W����L2Br$牟nnf�Tڣ0��g�y��I�f�!���S>��4��I�-RC|�S�u6nMz"~+�;�B�mh�oS����5�b~�i�Wr�Q��l�D>ǈ"Q`A'�.e�%y˻C�G��#��hݳ�_ah}���O�5e�C�ZG?�����/��.��+�IYv�Cv�L�~�4�n��hO��*x��������,TƘv���8�9���@�8���\�<��,;��HYsF'�-��8��aVT}rIu[+6Dy�~Z�]�[���a��h43�Q�v�-@!Ҽ6&>l_���b�@�˱�QT����]���5��2���1]�̡�fZ��d�3G1c�IE7PIt�ы���*0���N����"�,u���5��K��c��^t�U�@�Fֱ��y1?�R3W*�����ƤFg\��Sbki�+����K3����I�a�V�����kcr')7^^^�y�9�Ob��E��Lg�}N�8�t"1�ձϬ8�7�=��+�~��u_����n��"i�-�[��롩'�2��VCU��)�H��x��<M�ը�D�.��p>=����/�&��v��>�E�d&���Ug�38U�*��!�Yw����nrlV:�e�&��M�N�����M�]9.�Q�Z�& Zeq�����I��n�Ȳ��Ɗr��pb|����5����2~_Èف����	py��+���ݞ.��~�X볃X��6Ƀߞ��,m�o/�(M6w˸'���Q��N��µ�T��(�&Ɠ�"�)�,s4���\ҷ)u�0ik�L��Z�}�?'f~&h�=��u?ҴS
��~
��a������[���py�U���Cqz�$�<htK�p�}��@<UX� �,\;cj���*x��GL�����'�r�DM�=~���{�:z��,08�����[�� �{!�o|�H����ZK$G�%��x7T��}�C[��äo���R��iP��Jd��Mю6{�9�ZO�~@�X��|�[W�i��=^\U|��&����o	�p(b��۱%f����.H��M��Uk�5�}�ZG����+��IdVN�CeL���h�<�`�*>0~����T�rSbO�"�ҩ�k�M��Ob��jk���&��ɑф�usO����1PJ'	2�:�D4��[�S'�6���ŝF�=V�=��:N������o����y�n�b��qߗӽ�������Z��:��F��/{N�M�ɗ35k�$QyZ7��Y�<��n��p��44:���:��{+�W��<�#�z(�e��`�|U_�o�e�����X&1�<�p��.��/���{c#��E�~u��;\:e���D���b�(;6����eA��\��[c��UoR�F�<]İ[A�3�|^~�4�z����(8�Z½�q�\�l!�����}����۔��ZU{(����왻�J*���|�)�o���m��#1;,��X��~���j�C��	��^j������}�w)�T�Ͼ+�����ڛ$�϶ě�a�G�_��&��u��.��� 4-U�8zU����#�'�9��b�Nz>]x����{���;�)��Vy�tߝǾ���8RW��6&�գt����Q/�԰�U�<�ZV��%j�����>�s�������D}��zie���[�T�n�
����y���2��)�����\`�.�w��J��+5���=�Z��tǽ�u�NQ]�����S��e?�p����)c��ř�[����.�� Ӎ����E��_�18Fs�y�R�,�� KצU-3ӣ0�UD3��L��Yʺ�즬�3�9m����u_�Dl�ˌ-�,��W�P��/�&l<j�7�*�C���Ḩ��Խ{�Lw��S:(��ט*{+ ��O�?7+F�t�t��ƺ�F�7[�n�B�m���<�����3�%����訨A���嶍��1�v#U�Z8���	C�2d��Pj�ͳJ���I��3?��M�7�dD�p��/)���������O���w�j��Օ�����7�*ta��A����Fle��k2E�p��R%�PpOR!�V���*m��n;u�Uʸر�xs�͛�_�U9C~v"���O�T�$J�҇ݏ�?��6�4J��+[�#,mK��U���ޚR�~Fqe�k�������|��q�c���:�0&�qk�uA�Ã���#��2Zw��&牻�E�z�H�1aldj Kʲs�~⏣�~�}O�M�W>�s�j����g�wa�Qf"�7��ԆY����^���D?T�Rm�;�qX�W0�6	��%���ݹz����y�:���a��������$.��%���*��ȟ�j{�:OV-M���e
���7q�'N��Wͅ�ll�n�Te��9IE�*�a}k,�\�N[7f�E�fy�xO�類��=@�-N��L)���fJ#�S@�Ӯ�ZW���p��uٹg��m�k 6����;���>)�������ʔ�[��lXWTp�,#�xm�L��)�:\�.Kl����f8 7Oْ,��4D,o��?��u{��{y�Ξ��]џ�����2j�5�o�N�����*rm�XRo�ŝ}�]�Q�}��5�`2���~*�߾V���ѝh
��� ��T��
��6�!c�,��g�;�f�s#���n�j��{ޘIkv9�8�3�ōo��˱�T-�:
��2����A_�K=͋����!���;M�V�;qW ��ߪ����DH�U*���#V�ٰ�E�=BA�pc��Y������p��u����MiM�++3��m�m�����'	%.�4Uf�>�Ņ6����R��%zP�|�^# ��DW���S
w?p����h�E:��P�b��稾t��1>ŧ���݌`޽���3��LE�/v-[�����J�$_��Y��X����}�1М^�9C�M4g�]hJgTՙ�x�xb���gUs�Z�nS�K�e��/������1fJ��X�Z;U�r�?�hP[t��½�>]�����#`n;�s����N��c��~����!-�ISwף)oܢ븖��J�O�CS��/f�JF��jd��N*��?�VN���"ꃫl����3��O,#3�Z���/8����>���g�(�=�����ӌ�ޢ!9Y%Uj4���-q���n��=q����[=��rPA��C�6ϫ��X���f��1n2��1��K	z���Gڧ��"I��8|����*5?�r���j�-�9�oN�m�Nzk ���>ə3�N/["��m�n{��Y����kB���з���M�4��u-���v���w������X�-��^��gU9r2m��J��I��u�F˹o�_��fkG:֘hw�?��}_'xkk�=�Z敆�㝻��v�^�6��������/���٥�L����m�Ԉ-��w�e%wߢPߕY,S��s9Yg0O�F��z��Ú��]���d�:j�AK'3�)i<��I�>��is�[�>���JU����:���	-bJJÏ���2V�4�$W�1��J�gCݓ�;��S�#!��@춸s��Uݖ���]��J>�&�s�P	��u)�
��޴z䅂���/9E_��HH��������_eV�:x�U���c��,`�}{�2�zpq�Fs���94P\���ל�6�+�m7�p�b~����HG7R�3�^��B���4�b�B$�by�?rAc[چH����\ק��'��^oV9��7j"���¯(���[�#�{�=�c.S���2y�_������ݕq
�oH�a�z�
�����I��x������:�~��~<�R0��:�
�e���ܶ�8�m�و��Z�xL�3�_��W�i��N�Jޅ��xP`��Ʈ�ɥ?�FGm��Q�߸�l�
��Z~z�ހ|�R�)˓��k')���#��Ȕ�,a4A��.�-�y=7�3�=B�%�5�(C;S��P���/�c�'J����gݷ��+���BO��G<49i �O�Tb�����6ƙy�_�'S�����ɧm��a͖�нE@�Jc�I�v@>
�ngZ>3�+�e=����Ѵ���+�DR�>E�xDN.�K��`y^�x���
�n�D\�t,����2��^D++}��NO�����+锋B";�Q���~v���&�櫫��=Z����g,Weo��CshC�o�y���M�R��om#�eO�B���w�V�ٗڱ�+�x�������H_�|��%´< � lW����#��O+d8⬘:����a��ct�O�	�e:��fñ����3����A?E���b��)����P��m[G��J��v83�$�^i��C\b簚,�T�Ы����v��ViP�mF�����vw�t~N�K�h'�m] 6l��!��
���g������#�� ?S���/��� �N��t2��L]���LŴ�m%��&�P�|��ڷ[��6�9��:)�Hp:IH����R����?�������k�7�!�a��Ώ�@��cH�.�^�H:��G�W@U�}_�	�@Z�)��$$	A�C:E	)�CB��n�HJ# �%!q���o�{��c|w�7��}�^{���k��}G�R
E�G����k���Ն{�i��	�r��޼H����3V�Z�n��y�V�q�>���6�����ZH�bhA��y�{��m��ٍ��N�hl�7�A�)�h$���
X���Z�%�6���� ��m�s����怦�n�2�ÕZ��-2�$�����?S\��V��J |C�L�7��%�:|�*�oU�	�B��&ҽ]��HS<������2���@������3��Xj[�#t���f���z៬�GL�{Z�WsG���n���� ��ʯo�F�p��
8���]8�oY�������v�R[�S+q�pR��>f7f3��[��ʷ@-Y��o{�{�����0�Z��
���cqgQ��(y#H��b)�g8��x�t�@�t�d�=�cf	�?��.i���Pc��4��2��u��?߮�D۞�j�S<|�O8�`{q��9#�����
ZU�-ֹ%�8�D0��HN7�|"A���(g�K���@�%�vZ��h���'
��>	'�p�V�*N�jv��w�A���ݱ��}?�F�i�U����ѷ�D��1�&O����϶�5��ΆtDo�IB�/�4%�k����w�[��䌊�nlÃ-N>��I��F&V�I�o٥�S�n�1H��\YϺ�4>�����̝��q�:�uLN5��'�1q����/���U2���
�g$�Bn���L�6L�-L����`��ڽ�	��p�M��G��=��ñ�!��	>�w��G���*����RE�
������W]�a-�x��wXr��b���-ajp/
L��(��m(h��W�&b0[�ľ�6x�3��:SS6�����?�ꆖE��;����#7$�\TJ�+���ig��,��]ߐ�{�9|���qkR}�ȍVN�J!Bg��N!�Y;��x_G��p�9 d,%�-� ��EUt�-�1�1u7���xj�W��!��~�e�)].�\�#>k��B��6��87���П�c������o�:��wy~�:�%=��:��w�L[�?������`�é�����v~�j(�A�J��k=��:������i�9� >toU�����/=g������Ѣ�j8Wg���c����֫i�W���� �^@B�fD&Ji����
�[E��~��~s7��C�!�488��%^� �s���v���Kw��.������@.o���1�Hq��	�9��m��|�����٫�r��;)�@>h�"��I�43Ӳ� nɏ���v����]��\�(v�*��߿���'�7=HFnؼ���}��<��	x 5�������`������Z���9�LΜ �)qn�U�?��}'nL�@�����h3� � �7|Vk}�Zm!"��e��n��m\k"7/R
T:rjc]@�,M�m�K���o��{�Ƿi�U�t�S�~�s��즼t_p�3n��c�?��%��ܴ-� ��/��;]#�$�\$�qT�o"L���W#�1A���'�6Fh"�C��ʹw&�f	C���[��K�KqJ9��3?��q�zB{����G�F���~ޑN���ڛ(����J���7���-��D��}���1�`F ���t��0Z
_��1���>�6;��8������pc�ڸ��
nzq�]��ǩ�6�+?�E���힆�"�/W� h�Ҷs0_��v����.�@�*��?�2H�y���������[�ʌ��#.R~ߪ;�}wL�m���а:�ЏO{-�X�q��R�
�7F���٧s3���ſ�&D�M��v%� N���M��DG����Ȱ_�V��8�#\�:�W i�o�t����QM��to�,!ƭ�0@Dk�|��ƿ�aSl2s�A�����<"�w}j��@��ڒ��k�t�&s��J��DB}l�al�괲��<G�oCr!_�0�_Ť��-Xn�� \Ap�t��j��A�#R.��Q%��1�hŪ8��E�$�����j�M��a�}%��:���e�Ϙ�C��Zn&s�mⓔ�Xwǲy��j@|�ݨ''�����R���k>R'͸^PgN���א�Ƚ�'	�&X�LO#�Ú��[��i���s^j��0P��f���U���G�#������o���%���u��42���_}\�J6V��7�M_o�#=�?���~=MM�مk#4(�F�Gq��JI�p<�w����2�[K�;�R��h6(�fNx�`gd�2���,�k٫Z����¼���Jo�v� к�TA#]8��m�#ϛ�չ6�/B��;t���1���;�
H�AGDY&��d���FS2d�;����p�
��T��1#�;��̫�~n�+�\�<y*����j�=v>u+��/��U(�!�,1}�ýl�W�v�"0�\>����g>�����C
_�!7KM3A>�0[����0{)���`���p�Xz�!
��,�V/��KMg�#=[��)�J�t�'��Em�Iq0���Ý�:'�����qQ@Y��YaQM����m��^a`�5>�C�Uq9�2e�x�':a¬�̄�S�h��v6�U���]�
����\���4Hs,��B��V|��U17��G_f
_1�~��e�.�-������1�i���g�iQ�G|�?VD<��'1K?�y�!}>4�����9'pL���H��&���R�:�Ua�y�_�(�dM&AnxBt��T�ϡ����$�p�� K�)��?D��ϫx��?�y}�9W��'����/S/.S}����p�ET��;�(t���t�)��q� qA�s���f#��_���V�RN�V8�H�4�{�� N=s�X�֖�i��'����w�di���#٦g����ʳ&�l����ˡj^?Gi�$�A�a�N�g|�ux/��Ÿ�E�!_z���% ����̄�%(c�ǳ7���l'(9Ll�3P_Ɏ�L����͆?%���4tC%�Ø�b�M���I�fkd�����7_�w���W1�e �7�:-|���d���R��'��iD�KB��f�A���ql�_7�T������1�H�ɑt�1��K6���H̛^��W�K����\�?��
H7�[����J@u�-��/�hoQ�|E���:j��#2;�����X�����7�TA/G6Q�R$S�\a���� �u���94�v5��ذ?Ip;_�D��1�+,��")�N^!+�Dw%`��:���sg�@0@��҈߯�D �X1��E��?��C`�X��i�xJPR8����Y\�؛TLS�k$>�/,}L�Ql�F=Й�">�-蹊'�p�K2��^�{ b�V{~y�|��^��+��J-��]��~h�

SE^R�х3y���O�Jƶ��ߥ�2)�}�Yr��9�H��AQĞu۽<�3Q�69��	|��E1f����*I!R�G&�pÛ�eK9L��͢�5ΥY���&(c��-�/��{�;�~y��uἹ{�����O���������r(Z��kgϩ�<��\M���U������G_�x�W�g]�/��~��Q���d7���Sg/KWvb��v��?+�F,�G�n�Ir.���{c	��<Ț�
q�޽o-����`�!�#XE�|�TH~���ջ0�7U���;�"��s*�����=��zRVot�T2�&:;h�B�X�����֋�`]�4i�5�4��v�Og�BX��tX�r�d"o�
%/�p�P�Y�Q�WLʋߍ�<'�.��4�r\F�T�YfJ#�o�ƞ�����V��)N��^).�}P}kCW�S�ۭ� ���ø��~Rd�<�|��<-�ӫ������e?#ۻ�z%\�t�5��Q�^�������4����#�&��qK�3_s��{{��B���%j�����ѭ/��yV�I>����2J�bI�?����f���	m,�%���Ν4���?�,�}k���v����+O���A{�_�y|���R��m�=Z�mn���5ۢKa��-j��+�S�@�����6�xj��ZT�y�^2��̈́�e����#���u��i�0����]�q��svm���kJQ|&{Go�U���.xo�eڽ^K�jb�|k �aX-���_*O�>���w�i$�!�������F�v]c(�7r�j����@l�a*�讟?m������-  W૵J�t.>�yw���]�~�"�ȕ�W3���)mKZ���UAz�ߟ�j*�E	�ˢ#׆����lP��ķؗ�뾖,�?��*�3\�bi�Ԥ�!�__��F����"�"�2��M�rB:>,�p���XS��>ڱ
:ވ�U$����:%r�ʲ��kf(����,]~
P������T�B,�N5>�4w�y�2�3U���j��K���n�i���!ыX�*�ݏ����"�8�R�����+i��v
X��>�-�M���AF�sm�����n���>�(WYr�:���H�KqJ�Y��WL�B�\�u4mL�j��W�^�W���t4�I��9W*B�M��h[P�J����@@f�*vNyJ��h��;�#_N���fi�i��q:W��bE�����)�Y���A͏���=P�2�����DMN��1e��ɥ��O�K����/���=Cs���A�#�Dk+�������v����~y��{� ���}w����������}���B�4�i0��e��M]����E��^�y{�7��kz#��˜�/���w{x����dE��VX����q\���J��=�]�E���G�\�$.��� ������������|3+%W�U.`0Ҥ{w��*\��=,R7>b��+�
�����3��k=^�Bu�#�݈:Jut4O#�����mi,.۾��z%f���W�^�Bp{�
±��X�������^o/)��ɖ��Q����Z���T�����.ե�?`ZP�B~����Oݩ�99���Ͷ?��ֻ)T�Dؽx�P�U2$a漨�Ǽ��b�͋û����.xû7���0���������VC��7�Z/�婅��[з9�/K�ݽ}��<u�� �}��.1��	�9�Ѓ��][�&�ٰN������������ו���<���׽2�4��6!����8��6�3�h'���+A�����2!��>ՠt:>5~Ԣ���;��_�u�(�~\~}#8���o�lA�{��K���gh�m�x�/faں���������mN>쓍4�ĘW8_��p�'�O����s����a I���d����z(7m���S�U@��ޣ[��
�$��:B����Y�����e��%���_!��.�LR�@�G��^�PF&�m�!L��jb�����5P_X�'Q� �K�n���΁ �Fs�?EL���v+���F[l��߈ �5��]�Bg���;�\�O�^O0D�R~á>��+�\qjO�9b���D��ۈj4�N������.�a�'�'�!mx��5��o�!�#1̕u����d���~� )p��:#��<af�,t���4�7�p����*J��@#Dd`���L���h�<�;y������
mx�
-t����ᓻP�.��×J��ڝ�5�8��	�7�_[�/�����nrѧ��'�4�% �6�6���[55�s��㗄����C�Z��|�*7y�����|j'� 4���@���۠q���un���bd��o^^��~��	�9�Z��`���S66N�-���4Hb�3�^����i�ysV||��vF�D����S�Fk {�\������^��i0���w���y�5���:�l���т��j�vP?�|>�
1��RRV>+nr���,��4 �&/��%ke`p������i~1&%ZE�Z�#����ȸ��A������7Y�=:_�?��>k��A��
5N���&N��w)֟���Rڎ��k���y?�z��Eu�%��5���/�ɭ}[8M���m\�V��)�g�ٕ(N��6��PZ����kgo��ZM4��mSA�|:��������U�D������χ˜붯u[�p=T\�����2>&BP�O5��v�����hl8�Їϗ�����f9��de�HI"���[�����*�B�w�n��Rn�;���˷�~�AP�,ec��;wNP,A0V�.�s;�|��\�:UM=z ؐsެ��r0]Lv��W��9��=fp �o�1�ˍ\ɭ�~%4�b�E�CBE�p���:⏒�n{Vz��w�!|
��^��	�~�U^|D9�<��k�c�*\t��q��f�W��٬�UX���1�)=t�RK��e�go̓,���q���ӈfC6�(���Ysݑd����yӚG�>Ix�|'!��^�|�?Y!ގ�ll����	O�u�W>_��dv�D)�W��
;�$Hs�����1O�%�(��Q�n�f��7<�75k�U��Y}=��s�>�H�F�'Ҭ���b��������9�6�e���<��}�f5�����z��Ÿ��[H��Y���85x]��?`5Ŏ +v�S8�e��\B)��3'�(X�]ܢ�hϼ@mU\��K��Y��d����*V^�#-����~fu��<$��������6���oL�^��̡D�u[��݀Q���H�Zk��ڑqů��!�A�"�p٬���B$X������N�#=
"/�	�j��f8��z"V�)1�<�?�9P�
pЅ�G�̄>�1�����7��@WQ�hB7�_(<�&ݟ�۸���ͦ'�>�����]N�� �����v<t���3�I��/��bp���ڸ�zd����q�C{(-�^@��r��r��!v��#��}��o��v�b���/aF�]L BR�$��)��X@�p��������AG�@ੱ��ߨ�=
�qմ��-���}����_����4�l���%0=��-�	���>y7��ʿ@���=�8ΰ�j�dJF27iq#L�8氻ؘݳ[)q2��O�L	<���G�,�M?=��-�ky|��lM�H�H�3�	���%:cX�r�2N[A4�����>���S�y���'-Î�����t9gK�ǨI�
��~A�_�*��`�0�P.���E�T���2fg���X?�a�Px;U�Z�����>��^B	�E���|���l19ě������C�,�[�לAz(B���`+�9uZ;����f��S`����B*h޾Y�02iI
��\= \d(�9mV�)g� ��S�=���\>D"C7�H�U3#��q���$6D>fp��sTV ���4eV�?��"�ر$���ŉ�	I1@�H������e�}A��w������^`�,Oo�n����4)j��}��S��Mcc�q9i�y��a3�&&���V�N!]>d�m!C'����p}�f[�~F�O����?�e�}����`vd��H]"06�2/-Y~�
玾����hv"520�2(o�Q52�Z0sB���1�S�_��A�(#�/�w~��o���?��j�D�8He&�h˛.8������a��m����#�BHX��D�# A���>ǀ�{�������ȠUP�ua�]#0����S�D|���RlJ��s�az��)I�ߌջs۬�U��G�mt��/�w��2>�P�������'��T��I'H�����=��_����Z�o�Ǌ��k����A:)�	m(j�����ł߼2�uB`�}�瑅͆�L�Ѫ���R����3`!-d{�9�'��n�\V�4����EO<�T�Q��$H���� /(\%DĬ�Oa�`D�RY��T�(ʝ�j���&��WX ���Y�K�J.ê�i9���]�{@��B�Ӿ�� �(	�  ��4�p��x���+ß/nsU��"D��67��.1�j!0@u�Y�#�{rm �"S�!����� �a%���@���."�E��D�� Q{����'|��em��@�����	������e٠7�	�J�j��Y�ŷR\K�zQ]��X�}����"��A�S�nu�%�缐֭������R֦@�kيc㽩x�� Ah�lS���h�6��c���;��,Ȼ�	|�ע|ܤT!�/Q��1��y$e�!	fB[pM��}
,@��5� ���&��{�8��5��W$X�㗉�b|ܜ����+/�q�Y����3L�Fa�������Նed.�j1ό��p�|�Q�_��kZ`��O����zH��6/�+9���~��,5ۂ�<GCW(a\�����#�xz����6P"*5���b��λ��ȟ�_W���yqR$�T�Npi��[VV��w��N!cjxG�dXP�'�����<~&̚{����_�.PA�<���J����G_��7�eVo1�?L̰�g��,���oW%�<{�|����b�*޿w^1�l�������l�2�h�Z2��US����!:q��L�G3�pW�sz��u����A��Q����L���e��8��5%EQ^a\�}n�5��O_G#e�B�l��S�UH�9��>��y�@�:��Ϙ@?B�tHho�3��e0�ѮK� �Q��#��n��(�)T�4׼1�Q��5֘M,��o� ����I{��s�L`�{^z�#���%�Fc�� Ra�wo���(s���E��y<�!���	�늟�P��ҧR�c�ģ�W�O����~�AZ=.*~��w�ga��X�(F)/A���b�fY̛Y�Ӧ��pؘ������0�f�y�h��i5Jiz.j�R#���E)��a��7L��D�����Y鄲s)q�{#+��"
�c��a|��#@��+���e2��
�N��Y�ck��f�J%���
�L&vX?Pl������gr,=�f������ȣu`�l�z��V욹��О�#�oj控��Ox�2$Q7� �+ �] K7G ���.$������yKht�z��<>�U����\'�8������<�I�HP�`�1�<�X�
������xl��ag(�!�wH���ڦ�\X�����b�x��Y ��UD���F[Gj���c�k/ �ڒ@7�Lf�,1HX�kw��>F���i�7�W�k��@u
�g����o9ߑ%/wzR��M?%q�_J5o�j��_�ѐ_⥏�'�EZ��I� ��if-�t�s�E�B�l�������.�?����7�}qW�yy߿@`�;��U���{}8Rjp�X��z'eA�f����~�N�S!)$}}�O�+B:w~��wB���{����,�=[�V��:�T"�7�pYKC# @~��<����1�Œ�'�	C1�wA��ˠ��.*x�d��/��$w�@b��Ak�`�ȉV�$UET�ܳ�
b2 ��ac����>"�4��ro��D�Ħ=�{Cr��#��4�il�	�pl���F�1V1���*�=��?m=������=dز��e�	���^����:�\��N���������<�UI��)�HQ��^�����!�=��N;)��k��鵏���0PKzx$a]'��-!-ȵy�˺�-V������c��}�vL"�8���	�'���������6��v�O�6ҡ���o��K�I%�kf�n�w����L��f3��tL?�H�&#�~ ľ�S�2�6�J7m �i�Q��)�㝰Tϙ�eB�2�b���ů�)ύ�^wtX!+�jm3&<����fw���6-h,l.�͋�N7^(�����p���?��u=v�[�rV�U���D��n7�CO������d�7����t�qs��>�{� ,P�hc������%��q4�������"���X���T��O!l*��[;?��V|���.~��:�o�s��c.ĔY�I��~L����I��	`�R\�!ɍ<�t��!#��0Ւ����!MCC1&��v4��#
W�8ʓ1���0���c�}	<�X6���#6������բ ɂ�o�䢥�NO�S�ɫÑ2qf:�����ސ|�H$�'�c��g�S��ne�5������I�͸t��D��xh���Z��d��O���o(�A����Ź�ދ�����hv��N�%�jxR�7��(sHRM�����:����������O2DZ2�&���A[�JXHϹ�o���^ǚ�d��E��Y�c���炾�I,�� �?)���[�f�8�3�:B�+(`�U$`��RR�vYtf�E
c��.�J�n���Q�,�C���:D"��e�ViF�/Q��V���yFi�5��]8r1�|�9IM���A'���@��45|h�P(<�fϹw�OE��5��Otn���Ue��b���2�ho_��\���k&E'���W�Ĕ�~��efj!k*���馯�D�:<�p###�[|���|���k�E� U�&�(ʷG��pa�j&S�0�=<��k6DP�lZ
AEEG���O.@)�����)�<lrbAPrlă��o@� �2��}�"�M�{��Zd�-IG)�G*���w5A�'P����[�{��,�t�rR�E�?%W �"�����������}8v�B͙ 3=1�˗�Ђ��	G�%�`UbV�o�ҵ�BW��@��ۚ\�џ×iT�tf�B[fM+՘Zx�0E�glZ@<<T����.č4HO�K ��9X�@T\ �[Gh�%��FT�r��Y���E��g�s2᥽�%9�4ݣ��2�Bb���O��`/��'t���Ƚ�x�)�w�S=o��Ӿվ%�y0�U�0���pp�C�>�3C���_��T<y���#���h e�F
��3!z�� YY���hx0%��*z��{|Wd�T�!��kg���#��d)�Y�w�|�l���DY���;uOf��N4�uA!��I�d���g�ZK��ڰu�0Lc�S#D.�!��~>0��M2}I4|b�ɒf���9^A��d��ǈ�"{�`��T�[��E�^�L]&֋����S�?��I�")�P-ӵ�и�|�����222�3c�Yv�V�
2������R����1���X�a����bϰ�zB�~�FL`�'���K�Xm�Y��B���8��-�͛?�8m_#����3%=4�E��T�]�N��_���V�m��߼B��xv����{����{Ńa{��xNެrWT;6� �r�S�����U����>eCAtU~�ST(+Pߗ|�W��k&[��ů�3��\��#Ԇ�8zWQ\� R�����z�>@@Lҧ �+�{e�=q'��yB�#6�.�;��FG��fS�+��)#���wn�K�}�x2C :{��lZInY!2\�e��[�R*��� %��,$F�+9nV��c�p���<���9����Peљ��v{!�9��W�nd���6���O|����� Cܮ) 6�[vI�#L#��0`el�L@i��y�UڸЧ.��7�H��]�u�[�����-�l��L~ ��mT�$MQޝ���=�֙��Գv`�Q&s��a�M$^��}¤��e�q�k�=��%�p��/2��$Kp�
�$]��cU�8��G�[吽` ���BAI�'$�rLe�wnpL⧊,�>�Q����+�pGB9j M��K?ӄ�ή0B�s/~�1������s��[��!�BC�@�{�����R�*�w��)��B�t�"G{/���B�M�>/���Y�u��7���L�����K9�:���({(�|���Si�GeF+��K �bb<����X��ө� �#pSX�G�&?�5MJy2`���l+�< ܢ)��������Y�P�0c�U^j����	q��XC��J�ps�������=���s��@�숍����	Z�6�w��ت�����O$�#����ʔ�7����(�5 wܸ�b�!�b�q���D�
��L����N]:W�hA�phpx:E���6��J�uС��0�6�KpT��0�'Ć�1�����i�!�ϔ���>���RNp6uĕ�jj"�X	ǏW����#Ӎ��	�~���۠!�3�$��._&�8g��jK�o���2��'�"���ζ?+\�QJ���8jx�h��S��+4�d<��<lg-��WB^~�d�;*� VbǄ�)V:H}ZQ�b�~^��Gʌ3z��7�ܧ�r�bel{ftl7E�dDثpՂ|������ARj�S������ue��0��n6�[�H�K-3f�ƫ�O��.Hs��W�7��$�4Lk�tetkb�y`�"�/GF�L"�棂�u���A��+�nO�������a�HN�zݑDdQ��"��V)�?��h�Z�K�s�H�B��#)��W�g^�`��U����'+Zf�ᔓ�k��o�f+��Y)��0�p46q���Ϡ��z{/�6�֮r�Y������[�]
8���x�k�[Y��IrPt�-{�b���ǖ�#��κ4X'@
����ɮ�Ƞ�Pq��*t�2)�"�'�eļ�@t8]d���r�u [����쬉���^v���	��1�N���^P7f;*���j��Da;�=�=��0�G�A��+�g�i�$�'���#�[hj�-g�@�`:g�z����˜��U�Jy����\�nN�ѷ���U�����iJ�?e�*C�~��N��Q�P}�_�����@��V�SK<��]��S�Nh�����Z�I��z����P�HB�'��nw��|w������}��o1��ē����D8��b��W���dU�����~�LW��-;���T8�`�6(��LK�+����*����'L�:q�%�x���\����uS�M�!�m����v�P��a��Rh�X�8�殽!�C��ݎ���)ey1��	�����r��D���n�MFn�wsl�V.�<wՒ��Bw7�Dl�b9��i���`K7H���X���;��!���ȍ�P��6��"..O�H�v�MI���q�>�,? �Q������@���z:ޣ���O�����"ƾ+pJ����⧷(�a+�3+#��=���?��Z�M<���f2���x�|�UN-��߹�/���'r���%w�ً��:�^;u ��Q1�,l{0O��R�1�6��\Ծ[���{;�cބJ����)t"l!-�l�Io�pް�z�XrUL�*��4i�_�����=��5�q��Z2�)�1R���m^�j��D�p� �f�zr5�p���*�>����k'.��:�Mp�q���NA��h0��bļ��-Vݸ!^7k��_K^,� gU?�u��.(�b	�W&�:��ǻ������{"�U���}��3#�-�*�5Ի�����J]h���[�`������YWs�wW]],�Z��7���\����x{�qb���΢�!v7��r�lb����QnO(��˥(��dR�����!�?eZ�>y�6ddmr�rQ�*�t�J�ŭA�#��.YgF~�.;h�?���%�R���d.�L&��( �9��I?йQDO�}~P�z�#׮$�
�ȩw�:��+2ɚ��!m{�.��Ԋ���p�SBݍ�e�����sn�|�p:B�O�Ͻ \�
D:�|f��|�ee�C(�<&�2��{)��q��/����x��(���%Ѿ1�kX�ٳ��a]���p~vO�I�zT�݇��{U��u2��L^ �޼����kl��t$��N�M�%�?�+�"M5q�s6�8�������vB�$]��9�@SW�(��3N�^q�{��/_N��oX3���~��Ǭa.�786(�)㗗�ݎP���jH;b�;�����D'{`@@={��^(V�U?�q���sit��p���[����i���h���$��f僗��^m�T�a�G-+$\##vÎm���S�%�2��]�m��9&�����hp\DC8�Ћ�B ����>�=���<�����݃PJc��_�В��:����YKn����3�;_ҼI��?�_�N���v��HV/%M]m�6���OO��/�:�	0�*�k�z�Mű�{s�;,��$i�5Z�6+;�wi����:7�_h�E'����,���K`�9
]�
���.`=��v_�(���ls�_���ȴ}+�=PR�ʈUzjm��4��� �#ױ�Y���O��F��DJ�\�Me�#u�\��t����2�4u�	Y���(#�(�v���_���	_�$wb|����}��Ğ�����7c7m"�\l4r'��2��\�q��wysr2XC�Ws��DAJM^n_~�����x��<gy�%�7��pki���& ��K�'F;���Pv�ʰ�����h��Ù���	
�������;�oI�GtDW���@3�����)uwt��[@�ϩ�5^��L����}<���(7�T
�K%Y�d��r?�[�y&Hߢ���9t[(�
�%�ޙ7yF~�m"��=�yRi#����2򧥟���}L��t���Z,ȝ��~a�,�q@�=N}�����I˄�_6=V��b��t�=�{���0�;�a��佯]ع(>+/e��M_$b��N���*rm8��乪#^���q�愻�#�hO�9tX�l��m��I��p���F�a��f�ůL�o /Q'��������v�bV�Wa_�o�}�Ӷ�w�/N��$���g޵���a�����Z��M�XȘ!*1��ܐ�?~\�C�g'<\W/��aؙ ��vmIj��es�#�G��J45�Ii\��IQ��|9��d��I����:JyZ~�y���������7į��Y:�2O���o�[�9��6X����r�����X������"zlI6d����^q(��u� e�<���فrk�.Z�����p�y3qU�Fܦ;	w�O����>7��*�L�qM��p4�0�}I+?(@{��x�����z�(���$蟺o*%G��p/�㗼�al��/��=�����R������\����kA�0Y�B�zj/��o���G�ՌU��_P���7|�͵OU��B�s˞�q�vZ��M���R1He��tw؞�WI�S<�K��~eXÓc�H۳�?�C̤J3��a-�B }�N�#�uHx�$�9s��8�;�����[��K9�Stf�]���_T��t��,��eee��o�m[a8�-��I"!�w�>/���'s�i˗�I��E���e1̠?٘�i�r��XS����6\*�	�Q|��9Diu�W������~��fH��[a&�³��Ze�s{	�����G9�����iG{�q���J�p�v<���P�rW,���}:)cU�R���x�b_r��'�I}����6�bJ[OG��Ϋ�ޞ�J^����U���<�"� ��H_�]�<)�v۫��"�e �A��1KО����\�Ia��;�ܡ`�ڏ���P�����'
+�7鮗y-e��#zz\��Sm��Ġ�DUkQ��g��
�g��ٮ8��궆"�.eNO�D�T�;Y���,���C�TǪw�oGn;!ٕ�#'�Flg��8�Vji�%B5�#�9�4���t+��{�,V�u�{]��M#ps���ɳ;t{�r�!�g��V��IȌ@�)ʋ��Bd��qz��o��'ѐ��0b�{�� ���4ґ ;�ٻ u��9i�����K��m��O���H�z2R'^�Ywr��=�j������Z� ��#`�t�Z��ҝj���d�3 I�. B�ַ:�/̕�g����Cwx�xJg§����t2�Ԝ�"\`޽<�4�#>�v\�4�d���E|Bk`����ߴ�s�<טIo3���ಐ�(��kF�0��������ny�N~���B�t��,ݩkA������VW��!1��M[�muP�U@r�Z�����>m|��i�5�Y0�k�C��}
��|론��|9��Ӧ%�;3<,���h��`����Փ�S'w��������Y�yA����0�PUᚐ��2�i��U���Ѐ���_�
 8mN^��K�5
�,�����ۡ(���6�n���X+��0OR�pl�M�IZ���U'k#|	_:����U���-O	g��)���q���x=F�{HDu�b�O�����d#�.����,��Q��,4�
�Q'J�4���kɞ~�X�b�\��_���n-��
E'l1��[�w�OM�¹M��,��ܟJ�s�Gť�*�~�?��Ϣڪ1˼p��|�����`l/��9ރ^�� v͔:@w����n+�)�,\��q%���hW�e�m.���݌��1�wOW�.�eg�(��
�]}��b������NLH������E^N�x��7C1�"��Z�\\n�RL zw�8�;[y�!�p����"���S��x�V�7�ca�� +�I��W3��\M�>���^!�E�ȣ�gy�`��>�tE3�Q��@1���l�C
�gq���͒��Nf`���^j3��/�C8J��Ռ�g��.e ���`?�y
Y��_I{���d��Ί���<a_��؝0h�-�Q>`��)��Ӈ�3�d/C��*�^ԍ.�U5W�5z�K��</�W��!�ڮ���L1h��_0��9!��GdM�U�k�n��d@���ǿ>��pQ�C�)/�f(��M<[3��h�2�][��?�V�˷'ޯe��U@���I�Ī���������)� �zo�&M�G���_}LMD8��߷� ��v;O�������_z,�&�� �₊*���:�c��e �q�He�El��3*כ��3na��k��%��GRvH�l�����5����ci� �� ͚�\ �0w�uƧ}���D�繁�rd�x���o�uf�1���ܽ�J���Ȧx��B�1zx^R��t�"fne�H�Ӧ�`Kމ޽�m7���0_����j<�R����|Ȧ�����|���7��]���T{ݏ��qB{cB'�����$�>�n�c7�@�[�8�b�}t�� f�;�K�{��)��ս�Le�n�p,���k/�������x<�+�`h�@h�W��Q-</���@�׃�.��ܖ�ڪ���'�8�d�(ｖM��칛��_i� �9��0Cӽhip�k|��4����`��ޠ얫J����ѐ���b�Ɍ��G�W��Cr���=�t@��5~�w��d�c�ZWW77�����t��-���N#���W�l����h4ٳ7㺥#����E���r�#]L74̴��e15��jqIT���zW�̗,�<}��@�@��{�F�v]]��p�p�Þi���	U{�>5:jF��Bd����L7�]yש8�x~��f��P&v_E=�e��wp$�i�}��ȳ����#�/g�E�r�YJݍ�����ț�&n������}_����H0�h�z�ۂQ��x��c��4��m�BcѢL�����D�U>zMs
�z���
 � �p�RĮ����y��~{��k׫��tqR��x'����y1��wC��'���[~��$���g�����&��B�?�[�TOO ҾV�Z.:���n�����L�SV�淹DA��6]!�x���3�����5%�P�,���z��]�2U�����T�?�i����;���F2���+]Senq�~�����2S�a��̃�n�Y���.��2�.̤�g�������n{]���f��P��*�ǎ�eo�F���Y��A���c�@At����j})�z�m�D-ۡt_�	�x_'�ϳ�$����n���S� ��
yyj.p��ZXVQs6_�o��h�d������z$�G���9PL�@��]Ƴ"r~��d��w'QCv�|����G' (������j.X��?ҾY 	���{�.�h�~��أ/�f��=F�+��Yxy7o���{�A���Xo�� �;�y����MmM�h�#x^<ǣ�
X(ґ*�r,��t�(MB�%x��@��B�RC ��.��"��� j��~���Aa�5�f��yf�w�����/��ɭ���um�2��y��W�Oݫ�˴����Ta�6��I;���Vg�L~AY߇�c���U�3����fՌ���� K�Y@�kgR����Ǭ&H��/��xd�4]�_�_�����>��jnƯ�3:K�6<�F��i^�cYJF�D��Y�����)֡�����K,GC�Q�=L���%9`�f��|�Vi�}�㪱�ε
��kLW�JW7��bj�fK|�u����m>����O�<8Yw��@����^Kq��zgk�lׇV�Ƥ�����ϟ��Oʈ1=ѽ�~�s�k�qB8��6���
(b�f,d2��s�<)�N�eLMYc?��Ĉ��	����s�\�KvO�'�ħB��[^��SY����ʰ��'����xő� ��՚���e ���<�@Pk1E)SBcf�6W{b�>tn}���ʦ��ut�Ts������:P�y*3��E$��td��t=}��:R)qv���8͠�/Ap���#T���
����8?�>���[`z��W�\�Ҹ٤��I/�U<B����x��$-~�
��ީF� .t�J�9	I���W���$$FP)���nkq5�����/D��t=�e���ZXo�H�^xn nČ�+y9���3z��lE�ԥ�͛
[�Sl��2�ޅk��j�W:���SiR�]�e�~^����}� Y����>kT���zcӹ=S[�0�
z*SY��:��U���BC~D2�ڒ���߻I�ۣ+�>2P�|�-f����$V�����U�f]�+�~-('���Y8�hO�l��ڢ�O[����C6��G�a�D����x|��؛��M@;ۑY�
��!o�Pp'�P���i���"$B��[��]�����bV��ab����iUي	�9�*�<Z��O�Gj�qJ��h%5gS��O�<�������U�͒��ǘK]>B��/���f�jQ�3�A��Rl��b��I��E�=[�в�o�R��/ަg��v"�r��U�$W�ߠ��>T)VQ'{W�q< ��L���9�=]k�M�VDn�O
M�-D.�C�(����AT���5|]�Jj��fH�4<�_]�if��w���*�8�_D��ux}E.e�B��ɭ���z�㜠ᠢ�;����b���q
�X��@$��Lz}ε��J�㚯�����n�F����M%^�;�N@L�Z�Z�Rں#ս���\��*C��P��7�Sg/#ϣ)$N����\;K���T2�X,�!�$�#�%�|�|��,Ĕ���&˕:� h?�Ӹ��Y�������Z�?�����O�{u/��6�#%����>��#�>�����B�)�'!��zq
u�C�w2�4���s�7�#?ǟ6�5�������9v�!�
?�&�Z���꧕O�=��I���a�yE��HC�'��k�dq����th���\d�v��j� Z�rw��k�(Q�������2��}�V��n��旮���f�?*����O�����'oj������;�@i��䞝�n%x��"&�g8n�w�k�7=��+}�/�l�|&3��O�����8��i�L؀b�[Lj������bY)��,]��l4�c�qU�F�C�Lv���D"�����������A3�g�+綗����ۙ�L$a���-����QOKJ�R�ɏ����_|L\pc����S%���"Ԃ��\.;б��:{���޲�g�\�����H��`��IΖc�:�RX��fPc��5V��I1��^�g��n͇44�b��������lfIy+@��B��f�p>	O2�g3��'��
!�@�~����-���?�lT@	�)猈�����l��r��"^B#��nMo�84U,
*_y��sH��Q���ŠzQ��}}�E��e��)�1��ǎ�PEܶ�!���S�WNP$B���\�������-���H�����F|	����V9Ϥb����GgLܟ4�y�w�����>8
1���mDR��kBf밣:�Y*�N"N�����j!�䏑�����+C �a�sfh���s�6L0K/m26�~"����"k�}���n��M&���ҙwex�h��Q�BC�ӿ4���:]'Q��]e^�TN�q�h�`���,�4�5�tS��
Ώ�{uxHDD$��/;e�R�]B���9�nfij���sZQX5�x�>a����޾��47"[�T(+�|j �cIo}c<����^P�$��riޝ��B�1�M�|mrb@��V��T B�n��W����M�g_(%�V�1�־\����Rqfw�כo^Γ�������a�����k�D�@�&�:�l�"Kcp^z馒1i�U$�$���@sp\����U9Rz� i^�R��WG�O,?s��Nuos�K�����3�<��49�~6�A�F�rS0�:e�c޷7c�Ѡ��i�|bǯ�%��?rF
\������0_A��:
.깲�N��<n��!Rn������2�E�*G*����
޽���ך}��V*�Nٌ��^l�����G^��L��H�*q�q�d��'���C�b��L���&�f@�E@������SC3�Kol��2{��fi��H_ő�K4!W��z`u���q]i7H�����z�vcS��|!�c��0ϣ]��g���)�Y�(������U�f��g+h��ڴg#4��]r��^9@/�^t�ِ������2�
h��#������"�$��\�����7�!�V����M��ju�a�ɷ|xV��E��ɩ� ll�f�Z��!��@9 !�\���v���$r�Hs���'�X��Q�?���_���������%��3��J�e�0<������KʫO�i:�%[��<�&A-Y��@z�f���+g>�?c���r�\�d���BA����L�����x�I�Ec.�(��fQw�;��b����Wř���6k  =��D��Ń����8���s�n��b͡?l�}W~%�ר3�_��h�H0�S��U���c�,η&�����/\�-���5��!��`r�ɋ8	�BA4����W�X���4�~�7�Ѳ�?')-��'cӋ�Q�����t1E�,j��V �.��~
Qt������� �afj��_�rc���z�q��6��9�	�@y�'��B�ie9���|n�� ���}(��sm�YN�ҥǽ�+���L��o����9d%~&	x���Ͷ ��R�vV���͍�;�M��8r��|�1(;���"�?Rw���PP:f�eP�@�^~&y�aS�����쇇��J��,)N�W>%��\���%^��g�Yd�����%�J�vz�d�S���`�,�i�I8M�'%�������Ner���T�̤]Mẅ���yy_b Y�k������E�j�l@H-(q5�S���UE>ԉ$�S��x_Axy��i^�h�*{���4pw�7)Z����{v0��D+�g7��_ ��4�o���M4�f�|������[Iq�B3�\��J�R��D-�,9����=mJ������{Rn����N�{��E���p�&4O��>mꁒ=�Pd���; ��tR	�Uט8^$��,s�8C.7)���r��I���6��\1��q�oD�F�o��Sz��(r��,r��Iv����f�h��B�*�]~*��+���=_�%H�R>OɜVl~�F��	En�G�"m��y+��'_�Go	�Xz=��jES��hS��%�\@�Oи�{��H�L��R����,1akѾZ�{"�w_�|�샮{�|���__�ʝrU��������|�����4���c���J2c�w2'zz�^x帇�1�$e�'�S���K����-�=��d���d��8���&˅��F�#����)9��\J_�������'��G��4�{�L�!K/v���7�_�7h�/�ɚԥ+���x�0�Pb�u�[&��e��ɫ�S"';S'��g�of�a��A�Oz�Ir)��z�|��{�������o���k�(!��u��m/b���T�d$���n >�=�c2YC��W��ww_���#�r-�2A><c���h_�,VZ�U��Ik/��K0�,+�!\�wҝ`[�0�G�
w�"�����[�8����U��k���,���&)%7@g��vx��==��ظ�S�ԐH�Sﶎ��E�A:�l$zLVO3��w��'�s	{\�e#�zN��\��S��� =B����>��f�v��_}�d}�xSxEZN����[/S�Q�x
���M����l\�����G'l_�����"bZ#�(p��U\Y����g�T�"@�=����W{#�,-�ў$/M?;p���d��t�5aGI�l����'�S+��[�=�v��
���Q�Y�8��	���2_��}��i�y�
���Ʌ>�B�xY����cB���f�);�oOF�}/�2��6r�^.���Bb�i��w�1CÇ\އ��$��sg��RvPZZ��2��h��1:ȭ�LLj�N����c���B0�:��s���]&��0���/9aT%�4bs~�o�����P�!��u{�tW��,b�}02D�{%��ow��ښu�^N���uͿ] ����.@�����4%��e�<���[L���5�XP�.����R�f��E��}Oa�~�) ��W��Oϫu)�=Pb�dN���}__йCh
S�����*�S�A��N9���N�Pv��H�3�(qX(�8p�0p0Imμ[�I�hQ�xؿae,+�����;R����s3��y�x���D�w�s�+?����n�Q��w+�_�䱢��$n��1rC�T��\~��pb��*��T���0�T#@"���F�sP@4vm�09�q̝�<)�qs�'��%0���~��&�/�����*����L��@�;����6X���}��#@�sP�z7=��RC��O�	I����"��3p��d���Z�	V�iFw�e�z�)S"��Rg�y"�鹖U�|
"Z��GCtm�Y{�!���|�t5i$��WE�%��:=�*&QH	���I��x����`��{�-ؾ�B��v1���k�R#pg�]��Պ�0��I�
�������yʂZ���*.k�=)���΅'���4y2����~�]���T^Y?��'����w�2�7�;C��i�>']ט��&�ՁX���P��&E�M�S\b�L��מ�Y=�y!#����eZ٥m'!�?:�����#�Π"����������}e:aJ�h`��).�����|풰%���Zo0�������@�U�8��pI5��Ͼ�T�gWj�m#מ5����]	�U�q�l��@�)��;��g��KKx�F�Vl��|r�ڭXa�? Ma����t��������g<�j����H)��k�u�l|B�����Po��k��f$s�+N*~X��q�;����!�q�S��-�U
��Q��'��O��
Y�C���%69*pM�X�$̫ޔ�/�,:�rzI>���QS
:�\�����:$+&&����Z&�⊔���ϫ��o���
/�������]�Y|�� K�́��������Q�� ��k��:�a��:�>)��wǨ�?�P���;�=[���}�n�S�d�+'��|�"
���h�7�n�w'�4�;_���I�R�k	�\70ܸ�\��3`W����=
�o``��+Qp3�����ّ?���|q��[<�Ŷ���88�>�t
	���IR�l-���5\Y���ɥ���.�݃ B><����c�ʫdը��+R�4F��-���]Ս�F�+��g��]�wW��/�9���7s^���]��t�t��������2�\�>��e"�Ŏa��B���2S���ȹ��M ���C�ڙ�8��07('��a��/26;�S�����?����D�.�F��wI�.Tt;�?���Ӂ��ZQ��A��n�`����=�p�ѥ�4ԗCB�D�iS���o	��+��S�����d��-��Y6�Y�Y�o��U`)s�d�����ۢ��I��!�K��;I?���#��N��Aw���V��h��"�At{XԕM+��4W(7������剋6�}�ވa�=Z=l'�v}�D���o��R������Uy�.(������ҤW�ȥ!NEL��
@��>�6ɭ0y<��0�w����T8` ��N��H�eOh����ǅ���N@k}5[uo�j׊���X�S�O��0��5U~@�"ԩee���x���4?��i���s1��I?���**ĴN8O�=L��� TQ�[ g�� ��2fR٩/Q/.��;�ؓ`��@�=�i��&U�T��ѯ
f]���)4W�'��ϧ�!��^BW��m�#r���)������V����)��%�s��U���[6�Q0��|�~
`�W�'Ń,� �r����Jw7�|�l8�yA.4b��J&��ط��(��	����ppH�X�2�W�~�du ;(�k
Q�B�~����)��sLU|��d !�P�W�#�SJ�S�@�p;�~c9�	jv��G`f�ڵ�kW���
jSԷu
n"����:��T���q�e�'�v�{��X�?�=��r�	�o�Wl ���YIW�Ĳ�&��,V=�+\e�9 ���*͟{��	'��!����LW��l!�M��*m���P?���,#;D�F�2T����L'�yӒ��ˊ��c9�U)�n��g�K�ZΉ�{�k9b^����d�s�2��s�ܷ�8����P���1���F���)9h���y�r�)RU�$���h�tj�R��^�Y��v�MG�O�J3��w8ry��*,�Z���&��7�z�_�؉�| ��@�%il%����u�M(��8<�('�,��,�-�v��~�h9g~Y3�+0���JX;]V�o��s�c7���`�CZ�r���h�UY@#Υ�)ʆ���=o�nrO�ts��s;�Y�lN�dS����ɸ:g$�8���י�nk�؍�H�.�8R4��G�W��٘G��ߋ�H�%�VK�,F�UA]�1��R�����.�����l�ƕק����)�����W.G�s.�Y�w�L�8;�s2�t�=G��d���﷧/G7��z�rD����
��k�|��6��Vu�>l��#:�r�X�hȉzH���~�k+����V��������ߟ4Y�ٔbqy�L���;��f�*���S��i�� z���BW���w��MM���\���9U�۔�kb��,#�18<D��n習/����ç=p�:�2iQ�k����#�Β�=�����4�t�u���
�P�Q�@0C��?M���m���uw���$uŨb�V�ۊ_(r��P� 5Z��*���_g�:^y��[�Mw�Lэ���TUe?�PB�v;��jCs�9�z�]����h3�CW�@��M5���������JT��\���
Vo��X���R�~[h�`�Q�����l1x�@��[�m�4���	��������2z��Elm�(�$.��s��"T�/� :`��g�}�8���"ˈYxRSӡIx��r/	K�)x9�ڣ���-3�}YWegËP-�ve�fa�n�J�T�rC�����)��U/�6ҕ��aS}$�NMN�GS�؜[�2��\b=':�z���/��gchUE�U53�|�x�RO^Rd����Ыu����Hܝzq#B���;U�(��h�|�oD������逩�de:�N7'ڛ��Z\��Xq�(�����~�0]�Ê��_��2�{/�'�|2iH�i]7���D�Ay�����ϗc��r	�XЯ���{%�s��{*�֏�v��=��uV:��;���;��:Ċ��ˑ�c�EW��N[��y����MJ�Ϳ��e&�^~}	%�v~���e��S
��@��@"�3e*a���>��f�D��	�\M׽�'u�"����,|ۋ�1^��OW�Si�f�^5G Eǀ���/t���G�$Zz�������2,��[B�����3��^bsm6|�l�����v� ��a�|�Q��%�o936�N%�<��me���4LP��v�L�=ss��r��(����T'���|�}-��ԝT3>M7�X�*��B�ŪJg}����f?�>rV���K~�O��^N�S�5q�U�>[xOw�O@������m��>x�����8%9��o���y�d�b*�$^�k�����q�u���Y=n����r�h=W��@^r��l,7<Meκ�漑�,-vGk�4��o�n�������	\j�&&�S�'��[9�d=�$,�q [ʟ'&�[�k��B�_�kڮ�J�c�-a>o,�:�w�u��~O�wJK����~*v������Ԋ�_b
�1iI�|�$�vb�Z@�VS���>��
��u-�HⱩϕ�G)�����g{X(xoLn56�����S�c_����Ba��k�f7�N���I��=!�Z�T���#����R�g�M9�ι�5`<���hdqik�5r���y�E���h"%-u�`����i�_��*��4���j6��z+F����EW�u��2?�̅U�(�uq�*�6��`j�z�=���򞈿��K�ʋn+h�A� ��c S숖���tE���m��ZcA���ٜ��Q��!��Ό��͟%w�;��h��Gi'v��̏��$���d2*�FZ���	��d��e_��U�c�L�������Z!3n�e�k1)��E��]/�����)%�֞�3RQ3�S�$��x�{C\���F���4됁�¯���:s<�e�����ˊ�A K�Lڳ��J�ۋ�Qa������ЇV\n��[e���D���J���
�!w^�^�Y�Ў~։�-�PJ%d�wL�n?_��+�S�r��1��%F\p��?
wEˠ���@�YA\�x?�V��2��sF�.�#��0��E����W'\,�>�����_w����8����[-Ut�e��]X�&>N�-��Z��#%�*��QJe��)h-=fQ�Gdە�D:e8�������p�H'�X�{Mo�3�2�\�-�|�#��Sdw�5��cG����M�X�,s�Ƹ�^���B��rRU'IDK�VL����S�Ů�ʑ�4���_��zA�5����,p.���K��+ʅ��⥟���+��I�$��:z�($�z_S�]�\�oPl������أ�%��-m��|/I-���ˎy��uJ>��Q���i��]>����IC4�l�ԝ����L��)�7�]HY!Ng�6�H=v�>�1�S��J�F�T�OV�!.�p�hc٬r�1�c���E��D�@�Bb1��	���;�U�-//|ɐ=�y�0�����=�[����Dm2�/J顔�TNw֫6��y�.M��}��J��ܺ��7}���9��X\Q͵��������8�#�ڰ8��:i�F߯��^�NFU�f�X1�%J�}�w3:�u���\����!���V�����h��O!�T�ĵ�x�dsk%��f��f�t��4����dDt�Vj���BpיrLkk-��c�"cϽ����ٓ�B^���,C�8[ׄgk��Z�FsT�j�l���!z�E:0[.�4W��+-XxB�B��I���&�@��%���6jZ�	;��e
34A�M��{[�X�;wշKG�/8���Ҋ�_f��0�a��X���/޼�e>2s)<���J]�]��?>��&(,r`��)���\���23���פ�eհ��6N�}�*d�����	�����=J�;٢�͆2�"���m��"�""n�̽㒶�&��T��$S#�I��8H��1w�!���!c������1�[��q� ��Y�	�s.$I��{{��VmKv���;j❓[��I�0���L���r��e���?�<k'2c�sW�����x�����J�xa��^�l������%ΛbJ��f��v�綿1�d?�A�R}�0�F�k�~�pW�)��"{X�بCs���y�>��๾�t��k�3�ƽ.[D��y�Q~�LGr�TR�K����4�}�%s��~�}j*��+�1Bg�rf�
-���c�'�������=�������E�Z�Ԗ�m[�SӼ�"�VrR1^�Q�n����!C��}b`����Fs�Ub�f�n{��-���XՓǎ�N��v0����Z����f2ʻ�sX��*B�|���ư����H�;�dkTs�K�'�j�5��uj�`��?��˺��C�%�1�]3���A:�ݚ�~��#���N���eY��]X�j�@�����3�����)��:�Y����	��7�T�<O���"�k��C[��\_�f53�.�eco��z���n��9Z��>�925�X��5.;���Ǡ�ޫ"��3�T��K��e�n�b�~���wWR&B�&2��Ѣ�S����7[���_�փ?�����y{(�G�)p��`K���bk�Rq���X�V��>��э�ޟ�P�߬�Y*��h&�	�̿i��9@����^
�Ԍ��KYN%���q�p��4�mw�X�\��޻.��9P���+إ\$�(�%
���m���҈7eb�qxԦ�����^.(b7�@���Hܞ��1�9H�i�IRz�0꒰�y�t�����Rz:���v(1�����m5N����L�_m�0J�b�]��Vf��Ւ@|ޒ��%*+[�i��}�a��B�3yl�5�j�����'��W�.�x>�]�l,��M�t�er���"�5'�htKQ'�r�d��N3(n�����f��+�a�ξ}l�붟�g����������8\����魙^.E[Z�
ڡ�|��5}�cl,U�u����E^E�s��R@�'��F13����e�b$�iM=[ٯe���添�ˌ���(S$�$�)o��f".��>@H�?��uf1�T [���b�?]����ѨJ��]����{���2!���5�i2�>aR!&C��b���߳9��Hqi7N^4��.y���h����c
�|�!�?z��1IkiIYm�|�[��������HlM2ٳ��4�� ���+�-�c��r\��X�f[3L��p�;(bv�kavQjT���ǻa��!���a+����[x��;��b֔�_����՗̱�x��v<��v���\D�j���xg8�d�ѫǚ䪃�q�����>���=Yb>��B��dX,��[*������A��v�莨w]��p��ǖ"5���a/���[�}�Y/�3��8�FpfN_�x�;����&�_K��d���᜚��	[��E?�=����/��6WN����UX~{��rw=v�1Ps����h0��i���d2*�u;֮����B�vߏ@���K~�U�i�U�Io���%	�'�D.����A>8�p�	Er�%>�~4%a�YX����G�~��mwд���i0K��Ihzx[xRќ{4���OV���WBn�X�z���,���U2�&��2�ɸ,����ڋ�慅��ig���f�(?��*v�y_4��b�n���?VF>}�rާ<��UH��Ug��w��R�"T�'qT1C�jI�Ӣ7�ʽ��ߖXqkQq��D0:X*��봳�ވw�����v���Wq�WAnr��aC�J�g&p9�JPF����Ut�+�������F]�SI��Y���&��>��7�m�w��M�;�%�R�'��;L+쭧�$Ó�/�mkmM}����'��^J��\��d�_Y�V)ݕ�S噾�Ǭ��O��A��;*��C��c�~|�	j/�EA�֓
=n�c<<R��rH�����e�ЮP��g0C��n�V�o�������-*������`�l���h������B���8 �Ǔ
7�P�5�Ɲ�������=����Vf)��4�������~��G�~ :	��S�ʅ��XGi��Y��h�<oꇸ�=q5��1���F�GF�����������C,���.]��'�Gc'(m:*󗹾�=s����ܸ��j��wN��S������Ű��X��/I��	�0�����r;�_Ɍ�&d�8;�~y'�)��ocE��;���?=�rvo���H�t;z�)s���c�D4��J�/��@��}VQ��B�ʱ���7��E=z3��ٚ��8�H���a.�޶fc�5�E�9���%��8(rkV�s�X���cJ��Z��~zO���3=+ l�ԝ��c< [����j��辕LO��8�,X����r�B�u�u�R\�fO�z�����sf���B��{X�	��!��G�U���E���U��f��mDf��5�Lܽ��/��-5T��o`�t9�/j~�h���-
��΅��z�pv,��4V\�����ffl�4��a�Y#��1��s쮀�C"���s�
Ųm�M�Y��Б��9]i��"x7|�r����w�]���������Ǽ�������������_O��U��-�=G���E������N?$�ȯ�3ʧ���bk��}�i�0"s��o�gu�obe�CoGE�4PI�A�t^��vo���wv�hW�a�!�?�5�CZ�Mȍ�[9y�ćp���lTK�v�$1�n7���4�*�Hqơ��b���J��S��z���)wo����&&o>�V��mf�f�#G50�+�	�q��G񲃚[�0�7�g�M$�iD�<1~���I1�w����bb�d�E{*��*E����Kdajxӱ$N�p�,T��őJ�J��g|��:��rx�Z�ƪ���*?�հ��l��Y��;��ZFH�D������n��[���͟.k_�j��J_��#\����G�/~��9��ymӚ�7`�6TV7��2�4����N1{�5��JL��#on��kj����ᡢ�&�P��*A��³Ғ�_F�|����\�4R� �;��@"U��N?�I��*�r�?Z]ɸs�@�����>�F��vt���Ei*9�TS'�0Ƌ'I�m~L98$7�TC�;��{�k���r	M�Wlo���pH�j}L����l��	���c����|BT��b\)��װ��{V� ѕ���^k�=��_�AQVP½>�RF
��qݖ-��ƨN��M�]�vJ�"xX���P����s����ȁ�#�/fd�p��P;�S�5��	���L�[�@&я�,�t��D���0��mDt��!�6�W+������S���^��۾��\�K���B�e9rP�7���$�*uh�1��GC��]XW����U�Y����@��O�rnU����r���+��:X�e�SJLWcc\�I�S�8zǩ�f��W�B���U|[|P�q��90rV�x-*��U��n�J���/ݣ�}��:�*�ۉ)_"j�2��Q%��+��p_#Y�����R���+��	��hu7�	s��l��a��(a���[�K�q͙z'��>�c\�E�<^�1I�m@5,�18U���W�-"hϳ�r7m��9��`TI&�p_¼�����<e.���:e��
"ˠ�jF�<�4M������F����B��/Csl0T)Y�_�]ϙ���h���|�d�a.������;0��_蠴��8���L�\����:{n�L����]Y��.W�Q�k8��&�A��㼴�[F��-���lܮ�����g#���CO�:m�����e}��0�|�jDf2'h,�w݋\)wV�:��mo�b��~�.�[<�m��5��$�0�-�@�>��WH�i��.�WP�8�b���l������f����1^fb_�7��5=�A3D� �C�����#��K_��ǟ����ۻ�\<%3C>9bCo�mˈUI%̞E�_�Wu�X�G�"���To��O��VP�a�A�*b�"4প��-��{����D�r�Q��f�f�!���r�DH�j)P���_�E���T��4�9�̩����!|+��}��L���K��>7��gI�O� Ύc���>�q I�kػ�s����\w�w�}�EUTn�r��S����$��m���[�T�v����Sr��=�`���MO�%�oU��̔0��y�2E���[Y)��JU�o'���:���o�4}e 9����X	)Z5|`��w�^*��M���������0R91����;�{��_����
����t�,jt_��Y��A�0�a�B��r��+���L��l�1:Dm����12n�rg� �A�ۿ���|ퟩø�	>�$�M4I���XDp{��:::���/��@��{c��e�U�K�c�ۛίzk�v����9~�*�&���u�F�-$T�@t4�F�cd�BoGO^<tx%U�VI������3�%��2XX��Rnm�^��JM��Q��jȃR?u
f�)�K�KuB��#�����݄O�/++�}w�[�ρ�A�Ɖ��8�ǰ���Q�0��V����)E~��E�з����;��Z�0�M�`$�"�x�e�tu� �V���a�h�ذh��s���W���N%�о��*��p�c���G�H����Z ��"���'��}K�0�(%a�Z��uy@������
6�H��\_���?Tgdd��a���C8���p&�+�MX�[�׶��}��\���p	��[����= �=�!�,%�
4�ˣ8d^�5��ϛ�,���V���"��1�r��u��-F�R��{��Z܉X��*�Ճ����}�;�po���\I��g�)���������RUF��"��Bㆱ�è2��=�_C����Hs��,(BNz��Ek�4��ٲ�h�‐�J���.�y�꠼v���F>!���#����V��L��ԍXg���!숗�.��$��Hռ��H�	n�Xd�9�r���m�gЧΆY����;}Ō����-(D&��:�	U<Vg~��n���{χ�,v1�+�5��*�(,�0�/c� �!ܪa�5�Wb�{��,���%���.�{~���-i�ְ����m��xZ׽,��������_�V�[J�Q��rN%U����Z�)\o��R���ZC�>�9Y�����Ǉ��Mվ_���WK��ZQ'M�d�}?o0�?0��������ʻb��s����	XZ'ki."����Bw�tu��5��v7�H06�c2�4i7�q������3��m� �.<��<�;Й�����C�ɁZ�#FK�lP2Jv��Z?B��] ��k�(7�ɡbd�Bm��:k�Th$��8�L�)N�k�� �Ĳo��[������7_�&�qI`�g��ώ������j�F�'�K�4��Ƞǩe��22Pz�����|�O�RQ�G^�tčZpuD�$�̾�on�PL��2GG;8׶H�JGY@ ��4���4�;Mu\`�V�$:/�Ý4�f�J�=������Lk��d�5�uվ-�p��%�LN$5�E�U��bϯ�ӛزՆ�gӔ�J��;�ƶ�L#���m�j��!��o�$�_�Y����b?PT���8h`u�o�`�_bYJB�i�?�9.�\{�tw%�Zx^T��;7�(j�{�
S�Fo;$e'�$���I�QOi�q��]i/Lmmj��RgZ������k�b|7���KLz�m���)�.�ڂ�w俿H6�K�y���x@ZC
��A��,Z������^#c�;J���*|:>,j��	�3�Q��EUMr�0/�}�9�z�ϳ�$>>���Ϸ<El�0��*�x `Ƹ���l�UY��@�c��*��岾��3�-����(Ki��1A��z����G=oG�T�2�Cs��g�P �<xS���|N<�
!L]��oV��V��<��)ϨO��a���m�]�� r�'�F?��!�8���~FHXQ=} �s��]d�,�c
ך>�I�i��990Q�V��t���[�.XwSV�$[^��8g5Gdn�*��_6��)�Sx��B!���L)���S6q������"�>�v�vc��)����
z�����f}��&O(�@���J^��4����d����vҏ�u����k*b)�u��elD����ăhO��㙚�b�����̕����:�Z�(��R�&����g�Է��T-�P�9���F�[��qf�	��ᰂ�p�
�ж��$�;A���ˇ�=�U;ǗMc����uהX�\*5���I;#J�2�z(�i#IQb�]C5lQ���k>�k�g��(iFҹC����
��pN�7Y���Em���70xM)�; L�^HM[t2�1M�K +Q�C����Z�E4^(��̦��1s�?-&��	2/��F2�M�<0�A���&	������wu�y磌�R�!��q}-�IC2O�'���tW�z�Q/neU"����p��2�T=���Vŭdwk9��>@��(I{?X6�5��OF�kD?21[���� ,���RRx
u�2]���Y�y�$�v����XI���*��|\³^�V��Aӏ-�e�IjJ�o�ȿ�)���5lv_�ax�VV
�Jߊ��$�$1@"�p�{OѸo��T��4�O�^\uHT�5�T�{��<-~��X����vkP@\�e�:�ފ�v�b��o ߺ�>2�ٌj2��d��ET��Q��'�$�������px�(�(&I���M0�ǅw��Z}��kJw�p�m6@��X�+��J���8&�X��:�%e�0u�{�Vk!�`ySоt���]�9�=��+_�u���"Ҡ
�0�ˉ�[�sK,6n�	7�8�a֗���~�i�1��Nw�~�}����Gף�Չaz���ݢ��O�Sfޅ�L��B��2%J�c*�(U)u|�N��_�m�1>pb-s�@�Iuz�4���~sm߶��afs���\#���Rm�w��M<J�K��/s��qB8�E!r2��,�a��}ȑ��1� �*!?v�ܙr��	p5�))�c��$�|���'U�V��Ҵp��Ju�tYOO���K$�u
��c���Wf��*����'�I).
�`jW�APS`L�%�dXK��[�U�b#^�P�}���M���t�{��1화��As�F.�ݓ ��������|K�kb�#��m���=���K����]�c�_�mX�^��0%mz ��L���r���x.w�J<�c݅�b���22Z��?��19�YQ�[��f$�`��I�����!��}&���]�Y-�:a�beͯ�����|Qnfj||��b��x�f��h��Ԥ98��Ql��zmzg>������#�ǅʱ�â2�eg���چ��|ô|���2������m/U�s>�޺��a8�t����^/��vwc��������GyOi<~��D��k�Y��n�.��j�؋�5[|/��zL�.3�\㊇�#�΁�,��o�q}�3���}x�0M�	�O���n��[���ɺv�yU��>"�B���YhÈ������_	��C�ċ�#sg\�_���Y�L�w��44��%�QV��o�In��j��T�\;6����2�7���ސ��O݂zρE6�wۖU� �������F�=�m�XŐ��Գ^�͸t�$S�VN��o6����D����a�=ϹMJf�|y�0�k�W��;�/�^����T)�����x����#�toESB�.�$���X��A�4��#dɾ��)c���Dcߗ1L7KY#��F�6c��}0��=�=��k���~�����>�s�	�\~�Ϛ!�� �}�O���R��dyQfz���]�'��LW���5�gE}�=����&U$aJK�\��\�K�!�X�&X�����?iI�T.��J��ϒA�űI޹.H����}Vo$���w����o5��,=�W'�+4,�A(�~=ۏ�͢���������߸ʊ���[�^�����]rFs��s��>��t5�2��F�Ks��0>q�,��Q�Eӽ��}]�c��Y{w�"z[8ո�?/�=�����V��piN�# �:x�������b�'�7ƿ}K�G�}^a�2$)��Χv���
���c9��D�jC2�/x��2�Z�ܪ���1��nt�w����OrΧc�9=��oz��E���4$�Z�3$t�w�E\!���M�� ��1uB��ϟ��3zRb=��ʜs��ejR	�3�1ua5s�.�M]:|�|�k"A�+��Y�2*��� �p;ZϚv!��� ��+�q�ݙo���ʯ�ҋ�(���sھ�̴l���<������os�Q�酊/���� Q�UtU�绯�7�Z�+��#[g_��S��ٺ�;�jMr~J����
r�W+�����ޒt�|{��ٖs�أ�:�����1�����k3��eU�d.~�3A�N�ִ���Â̞O�C3�g��q����ГNp�0���'>0��"��ᥒ}4������pâ�!��X3ʱ�2�>1�/�K���4�|b"Z�G��d���7��|Ce��-�U+�N،����{��_�E��~*O�c3���>z6POeM��AU��x��V�OY5Ŵ�z���BH~���2$%����ů8r�ɲG�(*+q�$ܡ��q������E���p�8V:hT��P�~�=,��忦�,��Sy�U�,Ob���aMaP�N~-g���W
���I拷Iʔ��PR�|�cI6kP�nv��;]r�*���z5L�Ny�#2	9+C/j~O���1�4�E�O�֨�v&�*�������潘�x/.f�<=E�N�Ȧƹ����5Z:Q#�턬������/a�'e�i��iOY��Q9�%^�������)��O7�Kxϸ�hqNq^�����n�H�4���5���ϗ)xC@�_�"��R>2z���Z4�A��`SE��Ňg��.khE���͕G^�O|O��60�'^�V���v���$��Ii!� ��v%0�1�W��2��©b1����&�9�<3��S�z�����R*�7�x��ܖn
�bWex��=��U32�\�5�o�W������(2ĕ�}�^��n�։٥�	J��\�
�lno,5��!��z�m�����TA����%Ӗ�
�o�>$퇈d�J�����������9U��cV*�U�������	��WZ1�1�{���C�)�%&��f�n�®g��ӽTPn?�CF'��kEҎ�wFX'�v9n>�i����������MP`-?˅��H�-B>z�.���;C�g��C�~^o����K�7A��|F�%�.͍�>��@���6�9P�D���y��^��(
PW�DM|m8y����-�~�D6���'��@P8E�K��ceޜU��A%���v��/�z���8?������D�N�g�H�����������R��޷�������ߗw��,��p���m���vx�N2�s�M1=Z�j.�J�>z�+>��<�x���:ZQ<|� ��ۄYj���j!�ϙ����u{��`Ǘ�f�b޼�����퍼���;�ʯ�L.Ȭ,Cվ�yժ�ɩ�V�E���c�=�=���;U�-W���K�?�`?��#�P�z�տS�IK-�V����T�c����� �4�"o���!�Rh?oί��tN�٥`YژVf�!e=�N���'�n��KJ��#s<
*>+TÎ�W���e���KS7�~��2�^�\\���Y���U�%���0M0����CdШ/^�����xE��?�������y/r�ŖcrIa��?х���,��
��eX���WϦ���+�<�_��LձX��ޅ����?�Q.��ڿ}�JqԻ��O*�Iȅ9�������`m�M��h0��'b�����G�\ș$��8~�J��*(0vM��y臙��#�K~�0�gKs���m�B�7H�{>�����u?	᭸����f���#��_��\�G�<��˅�s0r�=X:����#3�9T�g0�,e�'�_�H�`(GG �z�f�3b������r#�@yiҥe��]����(�
;r'%W�{�~� %�J��/߹P�R&���^�S{C�V��W���pE�����z�a��m̓��s�f�P`�N�y&���ax�c$6p���ܷ9HCߓ$K��d�K�Z���������Vw�%�>��Y�e� �%��X��ޥ�6���z� ��41߸��݄^����W�,�[~�s��3ٷz�*'��{�8+S�0~�
�Y�FK;ާ)�!��I1{��hM
��q���c��`p3.}�R]4IYf��YK���
��ER.���X�7=�S�J���
m:�~���\�|?H�1  ��%��o-	�DF�Zp�:{�3R\6�L\�f��] =J�=Jrқ7��w�I8��qC�_$�RP@)v��X�������]�^G��$E��<���|��H��b2
��y�}xZ�Ύ0r�nډ��ö��S���r�J��j��: ���\PD��/O�1�F>D��uϒ�������H���]v�
�ݦk�����ң��
����⇡��L%=i�����GA y�t�����n*B����9� ��mc/��6+��f_��������kν�d��' ��b���_��p�^�,zB���\���*�d�c<�D���5�KS�־���4/t�{`�l�8k��ci�(BCv Z�
ɀ_����R��ZL���腀�x��#Z�ׄ[h��h�f����ܿ���rL�:��Rw9���c�[!�lWq2.T�>�j{Rl�ͻ�HP�Z(>�a�i�v�F+���<��r�n��u��5�9v�I,:��1{d��rj��ndj��r�-���o�s�� ��o�v:m���Q�r���nhB��9������5J�{
x�?��E��� �	�:�+W�zד�%��j`��@��YYT��..~�d�qáb���0Q�E�9qԅ}�5��D�y��.Ҹ�#H&�9	%������B4ib�:=Ĝ�ӈ�<����t,�\�Sȵ���xuҼL�۱J�� �R�z���<�3��-	�Eq�������H�ǌ�\SD\��X��7���2X�VQ��x������w-'����R�0�)ڸ$�SkB9��`�A�0�:�����D�]O�.7���S>�X�/P�nC]jn=�����ɵ���ɿ��3X�I�U� 8}�X�v�e7��#@设�+��;19�ۊ��tM꙯�l�i� ��S���,ڀV�*�����jkn>��ي$���xY�2����AE��E\Y���!������f�����j�!��IB��}�u�ލ;�\7����Աw)��rJ�-pf�1C0�1i$��[ik	�������F��	:fS2}e�{��AX,lݙ�����_�]�Ox>���
H��qs����c?�q��x+�9�
)z��ӟ$�?�y���A�F��N��CWɋ�Uy/�է���&��v~�f(
��	g��W���j��3N3X0�G���Dn.�SB�B�?�����M���e���@D	4=���� �({/�x�I4A���~9��>-k~���:�B;���K��5��^�tS�S�`�%*H�;Q���$�<Y��ʙ#?�6��衚�Y��r��^�kE0ךlu�?���ޗ�8�,4�u>͟�������e��@�/��,7���8�2�� ��dLC��V�p}L��X�I u�4�O��ۯ̗��|k�����ЏK���j=�W/�@%��		��<#�&��!�uS�Ŗ���o̊6$���kf�ܐ���|����]�j��$>���!��9n4���b�;�k�+ �s����F�[O,"�eM�@��V���Q�@�R횦�� z�9�'*p��`~��rfL�]ٰ��ռI1����F�+e �
\�w�ڃqN_?���RB��9O&H���ƀ�Ύr�⋔3K�u���Ę�B�&��V���,>Zq���T��駓-�
�C�'*f:�z��x�O}0M��x��U�h� ���D6`ј��O��D$�J�h�9>��aJ���,K��)���x�s��yh�A\s�㉷^E�W���␡6��9�-�^F��2ʋ�<�i)lÈ�����8���!.�f�T�ςe�x��c���F�}[�U�"�Y除�YW�+�t3�G���v��i {9,{ι����o�s�h����!Q1�.KX��1(\�&
?�n���o�<�i����Փ�Jn�ǅ0,7؄�N1W0�u�P
�aP}�����?�KRf��픢���]'rD���j�Z��?֪��k�r���+m&*��Y�� �nf�:L�g����[�}�����h񉷻�#�g�Jd���s����ꇉ�V��[�˪p<A0��o'�����\���g�Y��$�~�*�F&1ut���� o+���jfu;`���ݬQ�������9%{H�<F��6�l�3+wً1_@V�"��r��-0e��{ιx�۔���EJe���cR?S�c�7�]��ʀ#�M���LZH�LE�L���`�A��6&]���ߦ�ʆ�����T��8Yx��xGx�8 ���5����!R�	D�d^� ۞�c���|c����]��K�d\跥���G�]����
�8OX� ��A�k�R�����c��!����U�R�x���h'v��G.��L�C_B��7��0���� ���*����,�P���]�+��w:��s�i��K�S��C�$��rE��^�U*��]�o[��|���Ǵ�*#�����aG�J�'8�岁2�^WӃ�J�����k�eE5zi�U�t�U��*x:	V�#��[���
ڧ�$�0�y
y�ַl]�Xw�V�Q����?�G�:Y<8!��S��m�f�p�� �yDԘAeI���枙�|4�{�P8�x�R���7o�ϳ*zGlF�4��d��虗-:;f[<h���@�|�<~|��Z)��ڤM�Q���"����<�5gU�����\]������ʢ]���Y�g�@k~d��nvveS���]l[���~e@� �4���DVU}a��5��&)�!��`C��	�%�ρ}��g��H{���+���0��+i�B�D�)f��
b���!�!
D���6gw�B�(�R�|���6%.��5����UF���_4X3�&����O������]�Gi����A��d9�vw��r��z_'�g1R����]�1���n���"�:�=F�}���5?i���s��O���l�{���=6.IqV�ٟ@0�:��IT��2�ww/���2=�5J"�c�T�k�Z�����a�A����qZ�Ni����[Y��tI�199��ix�o��7w�U_��\���ѝ7|t4��t:��]�-�}�q�O����3g��봥����/Z=;	q4!I�_�8F1��l�ؘ?���׬��9�l�<������+D��/�+m��ʯč@�>�r�a�^�-����y+<�q�'�'(�cq�:�D�PJa���y�`�r�����s�i���,�S-k��X����{*\�.?�}G@�RAOe��g���d���A��)�BZ�*};��V&���R��؈l>���x����˞D Z�m�C�Wy��\�Z�\�Z�^}6U�N5�����wp�uPa{�:<���g{��;q��	0��?��Z�AlO��=D��)?MS���LR{�~mB�����@���L�����d�v� ��A����S����I�Ei:��W2�β��姰7y�/�� f�ݡ�i*Y|h�"��]�� ���۪w������5<�^��|�]��sύI��,S"�y�HZ��,z��D�պk��y�]���!��L�jZ5���J*�&/� #0:�g6w'�wy&�ѓb��5�7sy��8�u5!�v���K�����u�'��J�2�������҂��7>.8f|�Ͽ�s;��m����W��@+:`��k�~�lX�L�і��჈U��ҥb��2�M/��i�㓕��͸��%����T)�fmUsCy��jmk�TA�4+x~���e--U��<�l�4�O�u�����b�廔�A:��rd�[$ة�ؕ[�2�r���hta�g<7i9q��T��Z���h[�]���=M�Uv6���2fha�HE�M��y�M9ޔ��_.D���8Uj�w����O�&A�� j���9��ު���n-Ҷ"Ezk���N|�p)��$�rnW�E�|3���~�w��U��MY	C�9�_n�9�[�X�J���|>g�.V�Z%��6"�6�s�EׅU�w��$jq�,�t:� ��8��1q<.�jд�jh�n6���&��l���(��8�9����8���u����̬�L���L?������U^��ټ���DD�����K�5�*>Z�vuf՜��W��E��4Ld������|��M?�f|^�AB�_6���9F=,$�=h��m�H��RVMt��54�\��_���.���'L-2/���͙bUf!�/���ȅ*��#_~�& �0t�(�����7@Q�wK�#IW�a���׿�n�v�ru�}LD�o���)Skw0����!:���I�Pm�Y�x�̹�v.H@����[X����+�vi�;��E��v��=���Ɏ�u��ۉ�u���&qrɊ�@�v�=�a��jhͅ�RmZ�e���}οó��Y=h?ߜ� ��"hU��3E�*2��"��|ҰC'����YR�d8��ޟ8��C�U�u,��?��M���k��^����P,i���Yu����S���Nf��4.�zS�,���N��m�Y D�,̇���s��� �E��A�P'ZlZ��I0�������\Ȅ(��d�X�z#�Ͱ���ĿŽ`4Y����#E���{55�R��zY���[�J➿@�Nv;�Ԑ�y[���~��.>�,`��D�UUԸ�ǬէO�1ԇ�<�d�ݕ��\�q�����T�XEO ������DW�.co�wֱ�yJ?�;s���*ѯ/r��T���Ͼ�����X��<D�@�J�T	5�M��H=��i�Ȋ�_]F�'+9M�$�x��UUk�Մ�\���ߥ���/�	 i�����p�]i�S��z�n��+�0/c�W{��e��n�	Q�ꋔ�낥W�����nM����g����BO�,��ή���iM���&�z���:VcS�+߆7�N��}�
�Mg70]�-�ﷺ{�X��2b�̢��I:�Ĝ�}��Fi���¸��װN8u�oT�W���_8��lH�׵9!�?������DGZ��o��g��7��i! �@o�Z��%�\�ʻG:�EhH�Hl&�6!����=P�0$�˷O�\�+�q򈦘<�uSLC%�E�����F9U�@'�1w�q)~z+���7x̥���k��vאU#&���${����ⓛ�|�i$���SG��7�v.�p����q��Xk*��c�$�O̝�ٲ����Q��-�By{���_t2}]^�7��	ߚz��_\j��=j݈�#�������Niq��V�������ס ���]$���B�k��P�(���6<��p�����>	[p�-u��d��nn���݋������W��R��#=ཌ��S4K��"�v��E�^A��f�
��m�X�4�W/ h������;����� ܤ�t����6��/�	&����/J�R��wi�j�����9��!�ꘈ�'E�)��"_�?�����!$*x���bN{2���V�ur�&�C#>y�r����,+�0���E���;��~��]����ϔZ�.� r���|���"��L�5��WL���5>��,|���4=�tY�~����Ö���Y���7�W�ߖ�V�����]�F::�bL����nށƥ���v���n7�'d�1�F��"Q�$X���,rp��}a�$B��e�����
��+�T{�X�q`!Q] 斦���]�����,c*O�N�сϚd��g���H��҉}�*Y����̌�ѣӮB�xC��MV��&
�l�
����K�I�U�?t�]nP���J��AR\Do�qf�xp�q5x�d�k^� m"��q���zZ'�w��[o�m�*���o�Q�q~���2����y ���@������	d��m���.z�G'Rp��O�-������	h���&�}�� 0��%I�	�j�&#���sN�=�X,s��i .�)"㗇�7����%�(��i�e�Eg"9TFA��E����=��l��U��6��Q���5R���K���N��>��a��d��6����|g�i���v苧�i���*�g�L	�g'��`�~l�)s�|<|�o�۫��,���8/�v�@9����#�ΈЏ�@�~�q�ǰY�i��̉ZN_��Kc{�	���˼�S��B�؁��:[�?R@��Iyr66<�΀���H4��P#^8@��x��|}�̌g�����T~)�:���s����;�D�b�O�m-$�=�>,��r��Z�玪�a+Z�瘠'7*�S�[�H~%j�o��}r�+�°)��:�r���hx�)_�2������U��l�a����y�%��aO�b��Y3��
����x��y�� �4V��2�cj������(Dˋ�?�f����g��Y$�:��eWߑ�~���i��_��W5ե]�*IX~�9���-ڤ��0�^�[�`P���L�l��G�]����L֧)�Iqr����L ��)2}��c��!�&ʵ�]�����-Z�z뺻���ؒ��U�eT��-��pݱhpC�B�o)�+�W��[��-��3�?*i_X��\>VnTs��_  ���+) ����t��°<��k����p��l|�~�D��C͖[�  vz#��ed�]M�a`e�jD�p��뇩j��2�a�Vq���6b�PL�s4���7o�@wh�ȷ*[��G%�u�#����.	=�}J�XU"�ov��ā$��[)g��TQ�X܊��:d���ѠV��X�Msar䃽'C'Ƭꦺ6<��A%���-s��	�Y��a����ؙN{��E���O�4�ܧ1Y�p9�c�u�%�R�|��&�զ���W��׽�E﮼��(���	�2�������yft�!��3�G�mW*����ߔ�TU������~���c��|`��N�����5Sl�_JL�wm�Xf����lkk3-q�[a������8���I�� �#�G��)����h��C�DY<�?I�V]��ٻ{6���9V7����$����{�]L�&]fJ�hψj��Je=�V��A��v�4W#*����uP!����V(V�zm>���G�ؽQ(Tm�enS�5�,���hyg��zd!A˟���շ����$1I��@��ė�Y�����Fh*��$=D�bg����̞�4b*�#�J�Q_pK@�5�[K�vhf��O���'R�F���@����|b��X.���6��L�y���a�^^�/^���0�J��ʛ�"��itO��$�o6��% ��gv�x�-�Q��&ʔ�(����b#�/'��CTҝ�֎�+����u�߇��3��w��O��>�B�D	�����wB��=v�萾�3�Σfs��Kl�V(,� ����门�qu��1t�1�ux�*{��5��X�B�p�h����5�����0#���/���ԫD��?{;���\�R���W	��;�m�/�
��[-'+K��=)(�C�G�r~��]���_3v�U�1YQ��*���:ni\֟U��מv��j��]	C�j���.���~��j�K)����/�P���'��C��{f���wYШ� �=���]����UV�F�����!������eO��4n�.�<�{�O�[���D+��j�iO{I����0��p��U��_I[}=��4��dWu�8�V����t�O�+��%���KU��<0}P	��X���Bf�Z�n����L��)4�K[�`��3m��
�eȂ�e�
sH� V�}�B�/�M���{��!�*ꆬa��zb�"7�q��'�n,%�ڬՠ|%x��SJ~wu��mvA�8��)�N�@����:JJL�\�O����T�E@���2q���O!���&9`�6-.E�6s���}��3�6�1�8��d`[� 7[�s�n��	{N�'aT�;:.���:�+�*��yF �h/ԓ"�;S�}�?�2Y������L�o��bC�3b�˴�sV���=&YU��=��8�_��q�)b�z����z\(a�'M��D�.�"}ݫ�w�����`|E��P�\f�6 �&�%�o����?_�~��,tI��W��jm�8~�픍��ջ��@��OV4/D���\ ��Ehv�]��*H��P�!�^�¸��Eoa��&��?�xC$��WV�͹�r� �),�?WsY��#��]�v�&��ļG�F�X�\!�Nl�R�w0r���Uh}�����O��tzz�,�!��c�/�լ�8�%�ކ$�L�G�)���}A-w@&���7�Ȧ�l����٫Հ��?��������h�Gӆ\����?b���+_Mj��@6fǬ�a�$�Po�#���d�ݲ)��/��l�ɝ�O1]}ZN�ZV�1{}�`w_;�ߦ-�,�̨��iw�NF�o�~�l��R{��D���H��̭"��uX�ҫ�ЛFװ0<H��ȶ�]>z�
���j��2�ۨ�y%�u��R��¤�<��R><�A?z� ��ߢ��r�u�b`�;��B04�I�A�+��a��'���3��y �ֵ�-��Ū��Q��(6�qz�][�*�����\����{�k����>!������]\I���r��MJ������tN�h��x���b�4�+�FKx�S��,%�M�_�1vm�]
++��]޻���"�#�O�sC���U�U���b��i��<�v���b�+�N�>��a�K��ij��N��z�dg��f*������?BFy<� ���m�I��@k#1����P{*���R�����e
z�˾,W�Z�G���>��9��򾠏�b�5�a��o���G���Q�);�f�\�"eu)Ucˣ����ن}%�|�6��}�L�)|23]Up���i�2_�uU��k�&G�) �D���F��=�|�>M�k&�P}�YXE������.�CӯsoO!}�u�-�c�����1c�����5�"��*���@��޹����A�}���]������\v�����9��N�i�֩*L��p� RH@`i���!).bn5y��w샹W3��7�9c$XPw�o2C\�MI�]g��PX��0e�:J7[�x�,��,C.��6�\ґe����مAʄ`��^I�6�{��l� ����	��ȝ��߫n��ڍy6��D ��+6GC�S-�'����^��G� �p)��M�[���)�BJ���n	|�~�.��t՗�j�qm��)�>hSd�� �4��رQ���i�8��ɉ0�+_/%��22��O�b:���I��7���Q%�/h^��u�(Eζm��٥���O�˶x(=~��x�tY���.������������'~}׋ ;�U�g7�K����P0��3�Xߛ|w���gh�L����ď�#!�t����Qt�O��������1��Ha%^�o��f��g�l�y���(Q�b��/����������\��x�A��;`����>1ː���>�,}�1�t���Z{��뗕��yj4��&����TJ�1N�^�-�I� �ׁ��)��#
�����r���� �Q���ӂK���eb�� ��  0����x���̞��?����=i�t�mڠ{�֦�E���TC?(Z���j�S���P-�7vC~Q}��6���-T��N,�O�_R���.�8���xO��Y� �W�W���L�@��A��j<�ā�V�P���F�1P����P9�s�z�j��n�vé���g}�F�;_У�QD�^~��S��څ2���o�O���1G)ڛ>����ȭxO�X�<:�hz2:���]K<6?���A5���������D��D� � t�!l�{"wk]3������f��w�#�sr��̾��m���M�H��%�cZ1+�7�X����g��D�����h�L��1���!X���t������ ɯHEa)���-����B{�E��m��F�����o �SB�5e���o��[��o|Ȭ�I	vf˃���cc��A!U(�p�^��@�Ö��C�t'5����Q3�U�۽c���G��e~�&ml�Qpsb����J�hf$n��Z�L͵�f������Owa�?������0l;�}��L��b�O�����%�{�
TN˙#����(�<�?r�]�LU]m��40�k�1NY�/?n��j1<H���jQ�s=�u{!�>D;e9/az��L�,Hn��މ	�,�ns�^�޲��mÕ��yEhD/��H��@i@`�G�$n"���ښj�ѹ�@�<dzI'�0��"0�i�/A�0��|a�7��#<�6A#���>
�K��a�p���S,�H��m��,��bA��� e�y5ڪa)�\?`�ڤV{zx,a���[{�ɤ�������bv���Gg�MĘ�̋�����ۄȑ���ꎼݪ�l��Z��c$��ݱ�֧m���Z,b�����sx�[��̯V� �;�5װA�M�Û%�Fd�A�����NA�H���8�g
����bqnN�� ؂��rT�B�O�(�z1*=�y6�80��}p;S#�=���B/�@1�+���d���"K�f���Sҿo\~8�HK��g�sv��d-}2����@�|y�N��'��E44�l���?c�����K $2^ nwj�����/��x��r�~6�!�`y=�̀�?l *_�_3΃�__����(>�6gVU\�K��2a �3�j�e?�i�����`6��'�x�6�r6+���EW�o�d����j�$�4D�2S�[����|f� .���7�2*�Vt�쟽%�e��@���6 
g]�9
]J��������q�a��NM�����Ksﬔxj�c�Ŀ�+Z��ڀ�W���;e1�4�S�K�K�-��9y��w8l�s�4m�YnP��}	��^l�j���fS����Z�Mj6�3�0�j;��bY��wL� ����NB������\��:�:��#]�m����@�l�9*ө�\s՟W��Q�#�S7�G�n�s4�� 4|:�����hmd���")�fo�D��?goO��p"6�V#���}��Х0@z�Ϥ�{'�������U�.�S�vw���[)�7ܟ���������5_�NNjGW�:�����S�Z�0�m�odE���˹�t�G�����kx롲�i�d��V**/S}��p���Ҋ�Mz/��N�f��a�T�tb�M�}�0?bfBy���!\֞҃�r�~DA�N|Ed�vE��~��PY�i��_����;�f�U�k��,^D`(i�[i�O��G2%�Wy��y�P���Q���{��	2;�!z�����7:�/.Ø3�8��_��)��EZ�S3���hVt&���}z��O^���E.L������:�Q{��ѵ(��yD:ʓAtf��g���DZY�%#.Q��;�#��ZnnzC:�����&E��,@� "�O�~[�Y�d��\or=q�:~�S�#�U����5�4/2'T�_�33��5�$L�m�\��.y�z�=sx��No�D6� F��%aX4����}ޡ���P<]Iz?]��`�s�;n���H@�v����omC�	��ɘ�q�R'�d��Y�O7�����"0ŹC܂&%C��l�@��]���	^�$�S�q�[���p^M�`�}��K���B���^�� ,��SE���}��VP�*�Z�R�LKC��;/�'�}��ku����__k��n��12�����%;�N�����w�`�P\��gKǮ����'S�`F��$��;��P�\�=
�F�F+�z,������@Q���{�`T�L���?XĻ=��p$�Kٕ�}p���6�=˯�������4�h��Jx�'?H�=�q�5�%ΐ�)5�HF�з��|�@���L������"��p��^+��U��@[]ƙ%�Ot(1��Hz;�x_l�#R�m5x\"���(���X��Y��y"�3ۀ���/6.�����5�I�u�h��!�)^��ڙ��!R���ys� Z���]�xң1�:�,�CH� נ"��q�K��T��
��!{�L6C�����69�~���^����+��.��?�e����tTϐq[C�m�3}��vβzʐߏ}z� g�^=��r���I)S��鬮,D)��Y�)-{ʌ�~��1B��:��t��Zޖ���{.��ݱ�11|�X�6
tO��@�_��ۯ@�r�kИ�s��/���!:� T+b'����_�whs�}�!h��R����$?h�{eR�b4�Fd'�����r�C`/hМ"�v�%ғ�
�:���m?��d��&�`���%a?�}�Un�9�o����߉?r9i.����m�\qρx�:�VM߾I� :}]x,�ZV�H;�e��,����X n�
.��ͼGH~�-�k��y��*}��k{�i��ˮ�AJ)p\��7��[����Ҥ��� ��N���Ӆ��y:���[�m�wCX]���B��.�=#��͢��J|��Қ!Y�^���&\�k
��-��X^BZ��+(�`�m�E;��G�
��c��S����I��FDۓ���z��;�0��_���.O�Z;#���9�5�0I"|��|�b������8�lޢE)��r/�7�|b�o����,y����3�b�f��q�' 9���i���y	��XKc����(^�#���y���&��|h�X(��q���	�/X��(:S� �<+m*<h�?n�Z�����r�7�a�]XN��t�EC�2�@O�����֤�?����<l`�t�=v�}�����e��)��F������p#\����ܮYQt��Z`�`�m~��ψy��Rz����S�к����.f�7
�Q+� �
�Ƨ*��ð���^0n�pJw0��e+���	�M�&�;�\�Ε�ܒ�y;���^�_��:=�K�#@��<����)h���i�r
o�~�C�6ϩ��`x��(}F���@l�e�eq*j)����h�yk��)%l�͓�}��t6�<�Y]
�nZ-��}�Y-�i�6FQy�X�����8vmq�&��v��8e����`��.$�����.&��ZM3(��a�C�>9Ȑ��E2H.7����L��#������`�_�)���m{��pw����p��;����V
��T�5���}�C~B�,��&`)������S���v���T(���sN\Q}k�@e����Ǐ��̑g�vԱ8��QtF�#�H�`��n&�g�:���pG�ԑk��͋��zR͝�T��7�N���W�vAB�?��-��H�Tjq.�Lϼ��_߹��6�"����oA�lx�]4�H"9Y[c�}�c��ボ�P�h���2r�h�����M�׽ǅC�����q��/�fzV���GS��Hۈ?���9>c�u�*�y�@4`��~X-5���f���8�w���Ķ�vL�k�OA�w�f9<;��+{�m,�� q9���'-\�۴�1w�T�NtGߜ�@���=�;��ifpϿ=��s�����^	D�S�a'33C/3���F��,%*��^ƚ�%�Q���[��K{�fI�'�ؙ�^!�[3�T]O�@%�F��%;ٝ���)���"���냞��]A��w>jU��N���v��~vI���L�،������Tg�7�����#+SP�Vd�:�=0wL,�̬Q]��;�50���d�p��H#-�������R�ک]�RZ�.jf.�H$鱱>��-A��G|m���Z�;�-:Cf���%�np5�3@��jA;����oO�m�*NgY�(�F�^
�9�����s�$�
�#e[�?��Ra���Y<vsB�L�}��W^F(I����?�%E���D4��,y����SV��?���\q���'�� ���e��v��@2|d"�p�ccS������zjjj�,��K%W��k7�Ϗ��ֳ����2۞��u�D0*Jl]x߂��ơt1� ��ڟVې�-��7�������?��ܨ2�4�ɋ��hd�̋N9.S-�nr!�ӹ-i����i:)%�	ʰ���M�
y�lݼ<:�<P!���ڗE�~g�O�k]FM��dۨrq;��gZ�F)��
���ڲ#��}cv�s�N�XǤ^��ɥ0�'(��(�����JY*ju-r?�U������I|�]��"9Sxc̐%Y�����
�rI���'Jto#�n<o.��y8O���b��}%�X�����$0��߫,Gb����
q��c�I=���`*tO��&�	�X��K�ֻ�a�{�u��Tc[X� ��m�G�S��n_l��_a�$�V>�.se)ӊ,�6/��ՉX#�u_�_W�q{��pf�zƚ̊r�ԟ�=��>�9��y�3=}��t7ͣS
�'����"�L���w�pb���UɅ\��Dכ��(ăD��k
�k��-D �_�YG�:��4L�����l�ۯ���]�e�;��Uz�S����'+�!b_�ԭ+P�{pY=W�j�ꖮ�������R[��tO��7vJ�ͭO�$����^�u.�3?^:�mě)[?�>������$�o|g˽ݒ=���j0P���q��
��4;n#~�h%���2([�Zw�w�G�����^�K�R�%:t��gW�4���O��O}MMf���-X���YE����%ڬ�J��;�=\[n<Y�
�1���<���-wp7ï����K�=xw�s0E���G��[�_�ty@�5�{[2��M륀�}Ѷp����K�@�����fU�].���]/%��RK%��N44�ͅw�sv6��[��C�>��BݼׅL����������;)Pi55�$k#���I.�&�wY.�=�� ^Y\�K: �\�u�
O�lƾ��ܝ�|�C>��4���j����Xo�	t�<f`wC�m*�� z�7;ڻ��2�D���)��`6O�R�L�*j������8M�����u���ڲ_}�V�\�?q�{ӗ�M�V��J�J�t�5�4/��E-�mEJ�X�<��|�ŭ�j�"L� w?�rH+��s��[W�=��38._?#9oI���a
9�s�j�k�Η�!�g�{F�f?�O�����>�́��
�ܷ�|*&C�� <0�Y�˹ŗ�~��\�{����*�/�ᶃ��?�l�;Ky�8B�i6��i'�~<'����_�{P�'���t��%������S<��'~��ƨ���w�+�S�mCI�M�o� �����R���m*Sp����@Mf�h��kAE�.��� ҄`�AAP��K﨔 !eW#iJD�F��"UzU�5���~_��yo޼;���3��9�w~����c�uxߡ����ޡ����{�@���j�,G6_A�}H��\�8x�T�ǰ�G�umn?�8�ʽ�Xy<�5�߶RZ��Ri|k�����BV�]\�0&
�#pi�/���|?Dq�b�/��H`J���j3*� G�]�q��0��Y�
��5F�ֆ��:��W@�Z����[����""���H\�Y�T��H�`������t�6&4\�u�3�3b ��z奋�l�g8t�~�{C�V'
 ��m�O'C����t��J�nYS����] ^"�q)�4�H~ e�@ޡI�+�� E*BY��,�D��	W�;����1���]Ǭ�w���F����ڿ�?���m0(�-�C!�bh�X�t�2� r�5EYa ��ß�,K�����`�+����� �"�ҨT�Y�X��c�Ӷ�;�����,t��i��C����޳`��!��w��iJ�H�n���yx�[����C�@�n�>����g�|t�b��D\�^�I=�d
�Ko �PT\�
(0+NQ�1f7L�QF`��D�R���޷A�ؾ���a���?��!�8�u[2MX�T2s���d���`����D��%%��5k!�M�Ï sM�z}FR��̕��eǵ|��C��i��ل��(�W=f9�:�U�) ��V��^>^Ul�V�8_�[>b�hY)���C$�2o|���|t;\�W��t�\'�qb�Z
��w���P�� ��-�h���Z��R���t��Y	Oˌ��9���d>=�˹�"G0�����7�c�\}K,M������*̽Q�R8��v�EE{�Z�Fnk�)���ݼ�S�gH�S���&ӝŚ�^�n�v�����CX�|�N��A���*q�����*�Jj��^R{�čY��㍟�f�m���n\�?��y�(�d��Q�i�g��i�9��;��=ʍ�j���Ȟ Y�y	���qz�,$sH"�x�)��ܷǩF2�A؊�j�v�E���e�CD;���某�h%�vr��F7�ފ=G���&zO�����|�V�(E��1��*�`�[6��>��a���^a)�E�y�g��K��)������.�^�l�*���Z���䌛���������ʒ��3|�+�>oo������w������%�N$5�$��]�L ��E���-
%�*�S��� ׉6�OÇs��YB���Uѳ�-��'��A9|��KZ�Z�׿u��]�
%�7�������9J���[�zv<��	S�Ǆ�ߣ��ĘAN1�[��̨��A��\ۙ�������*�w7I��~wj鶙�E�fnoظ�X������XǯVә��u�U������f�����^�S~�4��O@�H��7W�#PM6�J��^@�k�N�Ǝ���,G�Z<�?��=v�~F�{����Qk�n�{lw�mxU�g�\?ˏ���۝�NZOK���S�;�`�b,܂/�q!d���Y�4-���$�ob����b�63V��K��{�փ&C	$ww�������s2�Z� �}l?B��?�n�=lZ��F��r%;?@o����[̰q3k����@���V�|Sr� :��5Q��@�#P���D*'���m�ƾ�)e�b^�wj	ZE���B�6�8���פK�9���R#v� �����cK���[�f/��>"���L����z-��#gn�6)8B�8��2D<����X�����~9h��;�d9�Ŷ��<�x`sʵ]n��f`1ҪL����\.V�YI0�w�]h�k9���i�A��3�ٽ8@�c7>��oח+���H Ԑ�aO���Kf��)�k5�$û���V�egb���y(DX32pTw�a�܅-N���o�J�<��ݐ06y��
��}1�v$�o�&Y��+�;�Ln��p��Ţ!3	Q���3M8֡1��b�Ӑ�J�i�B��g��ѻ_������{����m�t��XG���]��th�Y���&��k� ��҇�O�K����{<a�L��۟'�¼�S�ma��e�5D���]\�?}��z�`d�֭!r�q{�/�+A� 	@ (b������SD��cT�+A5R�w$��ڼ-���"7��ɱ��<��(&�>�?O����T5B�膎P�;� 1����#@��[Q�4{��Zh����C�mf�_��_�=.���2�(Y������~���/M����q���C�6o���ţ
I� �]�=�	zy�Rѩ((;Ϧ���w�o���p�{���u�\�\\���M�0�j����#3Y����.���[Y��u�u@�ƕ^��A���I�#�S���D�l��ǧ�PG?u1Ì���c�[Ua�2�����������Zr9��!��Q�u:\o@�,�s�>�ƴ@�_�0<R�v>��Ḷ�)���ńK�:�y�xs�H���v׀�W� �C]�K�%�dm3cg�ou�(<�_���,���PBaᅭ�H">�X�#ʧ�lQ��j@$��hc�rv�=-"���g��t��IDy��s\n���` �M=f?���F9gsDMa��ݵ�9�8_C|����l��'�9�pn���+���+��)J�:��ryO�1GIXUл`�QH�5F�&P�T��>`"
d(�u��A��#�,Z�}��m�:���i~U)���?<$x+6���~��ԘG�q��b(��*��KhmzX�<Uz?�S%�(���r<�v�k�=?�i��=�T�����V�����O�d%��HL8*=���� 9hy��+�0^�X��M%_~�G;��.^Ґ���?y�VKy��@zL�xL_^�cw!k�A��Ϙ]z����&���]�K�[5W�uc�ki���C�<����y�����X�NEi�#�.j��|���v���V���Mʏ*��f������wt��`���Z��^cT���Q�����S�Ǽ$vl9���E�g��#Ϩm˶�\86�z�=�D��X0OM�̀R{���{%��U���-c�8i����L΃��JSӂq-���h)pM֦�ƿ���M�oms�;+|��X�a����'��hxgQ�\9�]�� 'TʼS�d`�����7�;��*�3g�.4KN�<��p�Ja�RHF�?�6�7U7vV�������mSbV�V*�㇃��OOM�h�� ��"/�Cg[*�}���=w�\;���B�uJGuYC�	��Zh�Q-_��q�������"m?j�o�Ցjm��ӝ?��㾋V� ] l;�1��
7[3�I
TKk%N��Fn�X����G��脝{0�U �R@�矸~�.7���lՓS���K�ns������*lpoO͑�Z����G���Tk�AM�&{��v���M3p��Å�ǂZ���v��+��WF��震4�	z�� �A���
��ng܃��P��ҍ�٥q��<_R��>%�ր��$�(�$��p9?ɯ�����-r��3�`�JQ5R<듩���	0����A��Q��^��r����&��U0���!Ӑ<��������|�Q�������旹�>�j(1��+K�~���<��K~��SO���p���/f�����I8�����͡�"����; �:[�]yX�������9K�q
x��u뎨�9�P ����[@��n�Y�@�P��q�KRpQ����%����z_' �#�~�Ti& �����M���Zz��L6��?O+C��mG�g��TB	��8��}Ѭ�.��ƾ5�յ�$�/���)���������ު���dzoΡٲ�i����Z�Rv_�����эDT�}	�%#tyVcA�,x���ٍ	��<��0��(�pz��L����d�b�B��'?��F��Ò��ҭ��׍���s�7&S�C�ƀ�0��z&�4��cGδ �������ߒ>���Һ)�<���������q����U��$�����圷>ǩ+qK���um�;#��K	���?�zN�b�|�Xn���QrW��ax*�ކ`�p��.��Yn_���%�|UeU�ij̵E�(8=N���q�Co��u����J|S�I���L�����7b�B�4��v���D:)gy%�js�m���29]�@��U�x�鯅�����k�LzƷ��{*�9C�s�k�[ ����Ť��n�s�վ��<�{��*��򍛤���uu����9��& �nuЬ��|$�_ l5��c"]���ZT����:6��4e��M�+u�!p!y兖�ܦ#��O�{��Amt��*�yQ{In����@�^�4JN��,�T����ު�j���Z�� џ��q�DZ���+�)��"�v}XyD[g���]!�v���7r0����Cܭ�"��;�ծf>��P5 �O9��R��M��G�s��pY�>My�gL0���ƷS[�q�H�Є�,P�\mT�7w�C�E��:�`EBr;��a��N_�|��,�9ReI�Z���I�Ifn<F���.7�I�ۧcꮛ�3۬�̫�T3�C��P,���ؕYt��᚛x�T�J'�lW���tv����ZE3{˽��Ty�	���,��M�n�k���l9\'g#�gJ�.ׅim�`�+�A�z߱�^Nu�Yz9$��Pw�M�b�w�d�ne�T#�m,���:��-�	(�ʚЎF��]��H/�i����@>c׆�ޟK�Zz\vm���3t�o�E��Ƌ�z]��C)�F�,:�Ұ���~���q��	��T�ۆ�j�ə�E�ȝU���)Xh��v#W��!m�wb��E�<'�DQi�o���+CCI�=�B�Л�&U�i:�2x�\Y"DA(z�Nf�$u�	ښ	��������: �l�Q�<ڞ�\3��0�|~����ZռY����ɍ���VT�ϵ�~~�Ck���K������=�7��&�`�E�3C(k;
 ���=����3���+r�m�T��]�3`�tj�������~^��̷���y7xMZi;�+�C�eA�W��i����r{�#I\}X��{ɜԇ�X� �G���c��}DV����Da����6�^�a溺*��o���Ǥ*�tv��9J�͗�f���e���«�	lM�.���u�آ6�[6jༀW���RSX���[&ݚU�dA�uBɥ$<�
��2���V�����$��|0y��j��
���.lZ&�I��[z��<�fO˙z�[}�I9�ܳo���'�w�'��Öc�����m�t;ס3C����i͖r��΢2]D���!P�	�����o�Ik���B�ˊ#��߲
g�7�r��Q"�՜'����4/rڋ�����4�
xx�RZm7�6���]�p��I�7w�6�rO�#��[�ZC\<�[��bs�@��,o�`=|��B�~�
Ji�Ra�@�܄�w�zf�,x��k�ly\+���o�ʨ��>W�^D���������7ŵ۫8ԅ�r-�bl����b��uE�z�9�F3��c�[���p�t{|e�}/��E�HIϳ�)I��ߞ+{��۝�IY8z��w�`���7Pi#���ћ�]q����fX���'�~��eRnW��b��2��@�U�{{�#ZBT��ـ�􄀨{~2:��uq{!$��h:���D5��6"�,�T��T�]�OO��X�F5&����yc$�����}�[W&f<~��+?W�?��K¸�n�����B�}��O��k�.כu�%��ĸ�?_E:�;�(�� �/����2����N�J�)^�6�/����F�Kwr���Q���*G6�����Q��g�dE gf��l�X�j������sm��)����n��_Vؽ��^e��p���>9�J���s�����gs��`���&�`lS����/�8�mV�b��_c�E�xd��Mgg@�@**�����;	��_����"z�V�h	�
��9�ă��;�T"0[xי	�����Aw?�g>bT���~��/�}~����;߱wˁf�\oSS��_�zU��� /�@>��יc�C���H�U�kB�^co�<�AE�Y��'�Λ��,�z�ri�H������C�6/���D�̻?��_1�F�dz�-,� ��P��*��������M���c�^K���L���^6 T-um�JF�F�w�}�4oI�����u��b�����h��ӡ��]vlMU�vou'����2����rY =uLa�戄q���W��������!�(H(�<���A�GB;b�� ����	�)�'�c�7�����)�����&����6�6�	�x>���^�؟ն��sH������E��]&� �����y��=��;�5��_��d^�N�ߎ�_�8Y�1���#�j�i��/S ?+Ӿ���&�⮖JΒH�,��T
�����?�C;_�(��,��B51�����h񸊘�c�nr��<�O&ƭ	��3�J*�� �E����-���zYP�ԋv�m�N'�tr�L�-��<j��n��v���$�mz���0V{f��k	D�-�m��c����E�B �:Ɍ�7��K'���KC!&#������?�d����AЇ�3`�~"��h/���*r����z1�1�TWo�hj��g�t���(pg5�p�bY�7��խ|<!�E����jb��j1��;zbt�&��"r�3|�33EBoݺLZ6*���gl@�&�g�i�{�V�#�s���`��N�u.q�Y��2C��S� �*�g�s{^02:;�h&�`k�/�r��'���#�>�2�#e�;��w"�s�Y�� d�2�`3�q8c�@U7�y@3py��8�$˭��h�!�A�Q�S�-7~�I�}�����B�B�}�����\J�����%ʻ�)�y����E9�&�{���p���ĵ�c��� s3�c�p�Á��q���R�R9c�Z�����+�
�vQt@�'u��$�B_Q��2O�h��ԟf�ɞ���z��W7�h��~�����j?��H�d���m����!�J="��Z�� :)0���7�l;�0��@�
�p�e�_ ȟ(I$�{]jmrI�M��L"\�Ǉ\��3v* ?vy"9�=Ma�y�������c�e�D~KcG��#f/P+�^H�h� �_ڼ�O����p��b��!�m�<x�+���un��fG��ˋ�7�-��X~�hc1هB���~���.���E��c�p��f��9��^���Xu�:3�E
pF�{��p�ߥ�YA"�����.��uk���-[SGZ�6��3�h�*��������6�WbX %� ���[l��-�&Z���QZ.3�`�iUN���w�I�^��X�X���|w���AE�s�K���i�3�K��k��d��K�J���bKH���c/���W�
'߇������쟇BM���y�πެ�r�5�X���	�:��2������?D��ʕ�*��5R݉��Y �F�}��7gLj?�$�\^��4�)��9d�w[_b`s ��~aRk��(�|��S�%�0s6������C�;�t��������|Mh��B�-7Px��C�vY�@\ה($��J�e[��S)����~R廨ʧ�"���]�c	������'S�F��H���7N���G�x��Esk-��![�|�Y�8�n)hTY���{>�ak4��G�`�)���F&�l^NW|�S�J��> �%1$l=I�M�h\��ˈM�a���
��S�B@�PgC)��Nd����-I8㼔��D�:�v��Er��V��-_�h�V ����﬘�%��@��ڨ([r�p6�5�mr���MR�����R������sz^!#U�������`��a�~�XV��T'�`yz��G���^�
�j';:��8�=S�o,E�r��-̔:�������<��'�]���&���b�,Ԃ%W�+h�U#)��cf��V#Z|<�t�Ư������Ϭ'���+)p�4/l롻��j������c��W7V��Qo��ۢF�c�2r�`Q�/�f���L�s��r�q����~�h2LVUY	K�j�f�Ne�ƚ ���zFi�o�zV�N^?�+�$���J䴾B�^G;�0��t��T@A?{�9�� 쿸X��>�Rl��Z��4+ǿ6{]��pD����'d�.�5���3ڱ�j}|�\��n�ys�8v��V�� Z��8���e&���pp�Em���'��_�A�+�c�NO�F�Tȍ����*&G�����C�頾QN�	+z��--��F'���D��7M�v��6^Cz�Wl<��Z*���8m�O��y�K�g/���
�?�S7{� y�;#�Ժ׸�p⁨��_����O��{�,�S/�5{��8j-O��5��ӡ1�^��P��;ݍ��g��>�1}��1��J�Xt�7`?�x�o����4FD�qg�	�O=��i���`?a�QV�y_|QC�Eջ�Vv�u�^P�鹲z7Crd�2���񈪛�}���w�y���� (��60��[`m�yW�������ms�ػ��4�~I-��=���3x��*<1�٬P�n"Ǡ�ݳ��%[nW7	-����l(�a�t��,�H��V��35%�EàFa����..�vD��Q�I�LKn����"�}'����T����f ��0��%�>�oz[Ɨ���\����j������g4m�Q#�&g��f�L��)-[��d@$,_��z{D�J��v	`����{�����Ȗ��� xY��f"͝�6K$�\D���u5c�f}	�P:�mQ��Z�j6�_30�ӡ∕�u��TZ�ַT����
P��ע��%Vq�����߱������[��
*�����=�3�R��NK�}�^�h��W� �]��m^ќ?���Z����\�V�R�Z�s�-��!��l�X>(Lֱ8�DLDc�T�P�.�a�<�f��INn�!�D_�l�[��[ AU��|����Pn/�:���H�����/�N�#;�E��F�d��|	�@�����h��Z2K�^��T���R4�Y	n���]/�?���r`��[��<��Ht�q6��o���%	�^�2cj��捈�+y ��*1�,��Ъe�V(�K��j����&Y�T��B�8ȧ0ק&�[�Z\p^PQD�9��Ŗ�M���/�lz9�v ���L�<�t��#�LI�B��5���!T��t*�BڹR�R���#�h��kZ��k��#OK�yN��Y A��/{��� �S�X���)�ﹷ��ܬ�o*���"Of ��k���
�6�n��8}Iy�(�^����C��D�;<�>��I^@��i`���$�5���OxnL�z
H��o12��� �&B��c��Vf�9��{V�T�w�^-A8y���^���8�բ��ia�
��������Xօnw�]L�t��Mj�U����8�G��r�bX'>�������7�q ������I3gE*4�M�2;w�U�uC�y���}���3��qy�Z����&�Iݮ8��]4Xx$J�l���S�Z^�q��I�^&�6J��ή��Y��L������i%i�����AX���8o
����`h�ZE0�+wT���a^�뫿�~a��J���Rﳡn��_ݨ%� HJG���t�s�l��#sM��A�u�0)K�X��6��´�aw��'�)����s�s_s� ��~:�M�4+V��?�������-��Ϣ.#;��d���(�к�Z� ��wqL�}e/o��/!ǡ����~/%���H��a+��o
�Do�-B�k�$�y�_���C?"��o&��ڔ/���_���Po��b�6�� ��};!S�ũϹ̫�hk&h�~��PZ��#��"+D�&x&� � HQ��3-r`ޫX���W�$��yƉ�&��d�p�u��IH��Rϗ�h	F�\���s4�J�}��'03��@1d����|���|ݬhv��#8'��
��(�}���P(9*�>P��`\�z&� �w}e�:3.��X��5�K�X�{*�C�{�x�N�W-FMF��o.{��V���L�N�U�XoJ��U+�qG�ndx\JK�V����H�ܿ��6� ~ ����t���3~�;�B���J]^S���55�5%�޹��*l��U�"��^��z�Z�tא�CݨEՆ�F��8Y]\�pk>��~�����F�9Oe]����ɹL0�x�ܧ�U(@�@�.g�]�-X�@
�:P�E�����?sq�m{E{f~Gm�_���3/�:8�k4�S�N�_{��ZJ��z@	��TX�-��h�\r�7e(`c,![�������H�78�Aί�p��{:�s�>�5���0$����w��}'�Ԥu�\!_M�j5&��!� ϱ7R�s����0��ot����]�֣�\��p"��� �'�D�Ng>Qԧ'�~l�6�B���﵂龜mA��h��k�2�Ǚ��jQ����a<s�Ũ��&�H���������W����3�ȍ�E������[	y�)���~t��s�l��l�]-,xSQp�ި~9; �++�m۫p�G ���y�m�#�Q�HHP�i�d	Q(�n(�EЏ�OD6$F�E����~���R�s�I���J�z̀���ڐ��1R��lK.�{F.���Ԕ���6鲊�?GZ6fƧ4[їU�_*%o��4��U�H^ڥ�z5�MC��}�;1���ŚM��:!��ͩF�yK�c�d��-��R_U0����2~�Q@k�#<��}�fSMUHxs�1=Dx�e_r��lQ���K�ƢBBl��ф�)�$���,��/�J�FW�^6������W���`[`�&u=W�\6�&�Qpx*�Ulr25Y��I@��I�������t6G踒K��h�yqP�j�]�	�]�3��.z��+^���J��{�Ho�?]̃�b�+v�\V"Mݜ��ѴT�N�lv�� �dx��YaL�M~8�Jw~��G�̍VL���r*�M��r�6�,��d��M5�q�L�M�c��3��@9[b4рz!Ea�-���W��}`���Qf����Ⱥ��x�?���E~��u���˸���c���C6��Ja��^�	�J��۞�?|�w������9����&�N�[PEJ��7P�0���Y�[���o��d���0����g(+�h���_΍��(�dA�F��7�}C�n�GY�9dEəEr(�s���r���6Vr�K}�mF��wg��kL2�<B���Go�
�J�̕��وn���Vq0�r�ne-�Kz_��m�g��愝|u�KF��kAV�m�\��YV�B*܎re5˶�%߳�V�4J��Q��Τ�+9���6K��Y�͒��o��L�m���y�M�MY��AnE�D�k��w<�k�-Ϛ��n�V�׮�NvK�jx�Je�$���W0��}탵ɡ+D�;~��v��,~���Gv�A�S�(�	�iw��G�U����
�z�`�!�g����1(^Y�\�u�a*���]dV��p�=[x0/�W�RY�gnL�<��^�M��)�ӛ7i��V}.�!�a5���}�lS�;��)} -]R��~Gyˋ|��R� �y~�p�}}3,zʘ��t��r��DE�
r�ס�9�P��m�䇅G�zj`+9Td�?�Å�غ�5�6���ԕy��f�viPS�4�}�`��E��R�Ej��<��\�e��l���)�J�}���R�`��K� ^������jecl�8�2'	|�B�)��s� �n6�h��~*��콚zl��G�X-#�������������,��C�;�ġ=���'1dMqna���Y��3�s�t�O���w^��x�����Y�<#v,�%��s��WL��J�j�z��j׆/�Sfр)<
�7@N�������ZHҞߎ}fv��NRv#*�F I�0M�g�J���\E���2��Eg�2������sOȇ�+H�ý���S]�؝����6��Q-h�N�BҌ�������I�M0~�a�s��^2Z�(�W��t���J�m�r���fQnj~v�׸�ӵb^���TOSQ��Dt� ����m)In��t��s,p:{jO���l�5���̳�L�޴]�ö�M�v�>(��K�z"
�U��{Q|���e��H�����_�����d�?�d�e)�ܢ��)ɣ��b���]snv���h<���4fR���uj�����8}7I�g��*i"D�H��?�ɕ)���3=���lh�e;Cu��4m�H�r<����ƀ��#��S��'��T���C�mc�|Co�3n�$�sw��.��k#��x<.��h��e�φ�^���+w�õ,����cW��5mJ�i��Jxݓ�ya��w~om�jl��|q�CG>fn�I��t������K׏�%��*�M��X$ұe��G��oW�3����Ty<����~�5J���q���1�?i�T�AUE!tJ�k�ude���$.��;����q3����vQ^ �'E��Ez��&��N�&�rm!m����5v V��	�)��5Ɠ����?Q#�;�^�x,�<$���E�e��a3G4p��<꣋~4�
�z�k�sf:y��YL�ԈCg�d���#0��My�i��t��F���k�Q�N��"�tc��N�+�P�i�w�@EѽU�c����W�N�J��zg�%�&�{�'�� ^ަ��-��Eŝ��-�KTU����6s�G#mx��2 ai���Q7��[{#T�G�KtYt���iojx�N���y�?(O}�w���/�1�1�I��W�ѯ�Z�i������,Ĳ7
�W��>��߈�|��LR�����>�
]��c��ΩZ�HSR����BwS?�O��S�ّ��!,pт']�x�!,�#�D����}+i~Y��Βq�N�&P��Q�׎��� u�ٗ�)��?�~����@/�(M�/�u�v�Tv�?T�<BW�"�c�7s��1���(��G�y������o�+Kr�/>��KwG��(}� h�X��H_z������T$��7�X^�xޥڮOw5�t�����,]�T1ѡ����-�-TY�� ~h�,��Ѥـ�,�A\n�1�2�~@�*��%�P�Ł���\�pzij�7����Mu���u�<�pf�f�v.���
q:
:/Q�ȁH�E����s�e
H���8����3M} �L2uk�6ߍ��H��H)n7p��f�w�����.Nii�ﲙ{���g�8���%��3K5�x��Cm�K/]Q��@��J�:��!z�ӄ��G�(NS����^u��0� i��@�SZ��R/�s�
���7��|���h���M�߰�
�ǟ�^&u����N�@�0=��ӷ�;lǙ��PM���_ʩ�]���Q�!QQj���v*��Q@�eTqD��8l�*g������h��l@���x���5zᡧU8I�%G��:�w�GLN�ݖ)��T�E�Rj_��|���c�3O��MNǟ+��~��|0�@����D�0D#�)K���V���fX�S0L��Vv��KU�e"�/vQ�8w��KV�Έ��&�L�?�Gb���3-��]�Q�g;�KL��q�(�(�i����ڞ�������Y��29����û��A �������Ϭ��7A�&u�oѼ�GLa����������ߑyձ�A�y�)릏�8ʒO�J�Q�Ǝ�] �����թ!B���}M�]��^ZI:�=@O�3�)/g��M�����`4,Y��lӨt�nBc�����C�����?���0�s�}r/aS�� \��	j����Lw()
�߬��e�ţ�
�N���\����d_����wg���pI���(S<"�9�{R����X6�WR��	˼hO�sh1��4�G�U��M���3D��98vZ�r���<u��2N�HWx��"i���4�y�c
�_qَN���������;���T�z�F��q�(f���d������Oe��	�L_��/�Vy�w�vH�歯o�^�s��֦�å#ػ4y�I*���ӾT)|S��cK7�e�R�ڎ��9����O��\�b��&7���E�Y|���w f��z<�tn�0���AN�hǠ�� �=U�MRfɧ�EEMA*��rIz�å�ٵ�T_�*PU�T�m��zk;(��+��.[�A���e��O-����U�ӳ'�O�������j�pݕ����*�u�m��lC<mB�A��xe�$�C�aMܸ�3��U�ܟ�)�>�so���?�'X�V�+��Z%qM���s��lu����0Ov�����
���y6/g2�o�U�hqE��s�¢I��� �:���Ն4�R&�\O�N��3�yD>�jV-g��6L�|����5$���(3������~H�]�L\�\����w������LIIab_���s�_M�_��ܗ���������A�DW���OiEΜ��'��u���hq(Z����{�������Wqs�[]��g��_H�x��:j{�Ez�5!�6��Rԯ�<ˠwu�֥��h5iL�h��gJ�^k�U�O�oH�P�4!SE��)��w�>�n�� ��#^���@,O[�?G�'>��P�-�1ku��6��&lB�%�E!LJ�����Pa�Q�?�?��:�-���7<�7�R��f�E��d��.�}~Mj���U�P{=;Z3� {$�ͤ�܁���X-7��Wm(��0ZS�r6�n�CkȪ�2R?S�f�4?O� ��_$�����a��3�zz�㐇'L�8���EБ	�`�e3�� J��+W�����6M�ڳ�����k�N��|��Fs�^D����"��C".��q��Ϟ�q�ʞ9������\��=�E	�g[�
�����]_�V$��eѿ}i!��:7K��Xj$��qB�R�:�[����O��فKUß1�Sm����MYp�J��p�l j�����܊�É�Mz�X�Զ5�~��D�e g_�u�������N��P'����k8`���?��z����?sAd����B}�xl�.{KD��^�\��"%ʒ3�|%�YӠ���bKJ93$��OV� ������nkɿ�r��fy4�N���R�~����pIW���c&�7�
�곡�<|3ca~�PM�
�nz��(Aw�G�ߪZh	A	#�f_��B	�xh�W��r�a�������^�r�/�Lyp����&��?F�迿�Yݮ%�Z ��Nqm�tQ�#���'�~g��Dֲ���uS���ك?V~�  �?�3��U������/�w���������9i�G<��z�ո�y̓�~��c�#�^��_���i�-� �"�8�<Z����ܾ�����2���v�)�}��=�#7s���ȸ���Ť�il?l���]�� �r�wa��7}xo���* *.��s�N)���v��W�p��$�����/�r������M��NK���ߙ�JW����Ɨ֖S��ca�r���Nq*	 �K�
��e��
N0����Q��6�&$�.� C����k������O�·���Rƹ��K�����)QՖwէS<�K�k�ʛR
�v�J���9r�!��E��V��I�|�@"�ن�1�wBz�.xhG��dZ���cW�e rO7Q<�x_�F��I��Ley��@0(⦚�˗A���Z����ڏ�?|:f!�����G���'l.���9a(1�G��x�J�q��L��5�!�P� �ͲNH���ف��1�?}�񡱿	k����6*ª�)��o�S d�LL����fi}���]�K�@��4>����B\��M���(��y�D�gmB@��<�2̡[��U��*��`���ǳ�xo���o��FZTF�;N�����6O��e;;���� ��5VdI�s�r�Q) �	������T$Rk�߾�cC���0��"_�g!rA�;��A"�o6W��=�#Cc��JR���ykW��B�/��G���R:��w||�W��U�˷�E�'7;�/D����rz��`�߄�C��vf�b��ݥ�&ߩg�J�B��v��]�L�&�1bv`��/jք<�4}��pqc��T�)I�l������^u�$�r��ed�`�,����:vzW�I�Н>�W/_%6�"Щ+�ا�v�1�;oW����e
����A�RC�x�d���v@g=�j{��=v:`}�Az[ڗO�~i������3 �m�nH����W��Eq6N.s��,����-�iƋ�+��~�D�!��F�c��>��@AN���$��66��UT�8���ͬN�'���Ҏ� �(�vִ��.���? ���|p��/��a�ۦ��YY`2)���/�	5ɝ� f�������ӿ�����"�mZ�
�ޏ�.eK@IE��d�ľ��rY��^�i����]=���^c������ǰ
.�v���F.��p#�����gt������9��7l�NO�[��e~؅nHm�13��)�@��M=�S��m}������$U��R�Y��b@Oj�ڙ����~�;��q� �u~68�������i�o����oܻ������ܛ.@�ӌo
�\[Q�Q�JXٛ�^й�%�G�l
N1a׮C6v8�i����y�|�������E���E�|�F�EF/��7�<��ow�Q���t��!g�"�o㲿P��4�>t��u 5L|\��!�m�*v�	�O� I���Y+A��+Qr���e;+q��k��Mk��$(��o(d2�� �A�f�ٮQ�g�
]t~���b�§�]0���WE�߱�Q�<A�E����.� �Nvq���` |��������##����@�A�6%1 t �������'w���	� �@�VD���y�R=�H���K�=&�;�^�n�.�S_��%���{�y3�+ʘ|T�#���-0na}���~�-@wF�	�L|� ��M���2l���:5�]�W�e��K��}�C��Cru`$���z:������~
�=/�)��r2��2��x�h�t�;� ���x��5�*��\�Ose�$���Ǟ�� �<�sbqG�	F�ɕ,~��\N:�w�3�	�;���;���|x����/��o^*��f��V��N�Ƙ���	 ��	{J�j�SH��Oȧ�m�{����Z�c�xJ��O�_Ew��쫡�Ɔc�/^�}�����ӵߛ�Uq�:C.3�����A�\�ځ����*q�lU����$죈�������L�>�Ǹ�`˾�2�R�De�-k��8wz�8ƀ�V�l*�͏ ;�Pv��I���}�rSX�KoW��P���Kc��[�n��@S��}��'��`T��Ӯ�X�2XY���ad�{��F�� n����K^"~�b��j�/rۼ��\&4n,J��؍{{.]+{Љ ��o랴���%ȺG��F@+(WY�ӯ%�Ł>�ޞe�э�_e0��C$�C����7��F��~���1d��K�͖�Q�� �!zE�蜝���|�����6b];�]W4����?Gd�� t�-FE�	t��U�r�B���d����l]F�Sb��j���Xp���,+:�!IC.Ȁq�L��~��S��8`j��~� ]WnO&�B#�>��sY:�N>��� �((�н���F\St���EC{kk��	��I�{5��h�Zֳ=:��()��$��ܒc�>������	���'�["�PDc�>H/�����B0G���c{ɜ|��~�c ��4�)ū>M$&?�����/4����2t6�e��>���|���B�e��rf�=wZ�����\��h�b5{�Όww}:��*A�l��`�X�|�j-ɢ�x�nƥ�~��܎����pEA��IF��}{0�� \6�8��A�H*KU�t�`f���E|!;�^F\���/U����Yϛ�:Ƶ&GA���I�TT�΂G�99}>���>�q���k����;k������B�O(t�l}y<������n��n��H�,���5(��}m����WeʖK�*;YʾO�f'������Gx��}<���3����y�g�xfn�*�-i����O�d��d�9t�ŭvB���S7��L�\������m�%˶�*�[�r�̶�JW.p'ik��7���b��������Su�
������G�K� ������ь�ڬ�O�pg/n"]�)X,vj쨍�C��V��8�{x��N��o��>|�a�$�����8tY8R\�W0o$��r��cp�&Msl��_Vh�=�rT�z����2{Ƌ�p��+Z�!��+��RS@�����6�A��7ݐD$�b#����4ǚIn��_�������ۘ�vW�\N����KE��[u�iƏwH���k_M�l�h�a�k�]���TnG��f��+�؎���"뜶�Q�U�����ü t#K��?tˆ|.Qm�[8��s ��+C��VkvUnb�$w��Y��=UA$�[GۀP?��J�
TDٽ����KJ���'�NU괧��iQ����@-p�����I���4#~޳Y>��|e/?��=�aoI�s�.�a?�苾�N-�w���t�;6��s*�����0�W:6d�J��{�:��h|��'�)o�s�H��k��\�|�&�V<�l��/B]y?�Tae���8���0�.��#��؆�O;,NB�������B�;�?�gO�a��N?�n;��`\go���ʒm��s3�5�.K�f���u��m�����lz��5��"��Y7t���p��ħ�Kb�e�Gm(��/}��"�芍t���e����o�~��d�CP �+�8�n,K80j���n�o�tz��T4�����̹l2�+�➞�|�{�g�&)�q���a��v�d�a���D/ǿ��G
�f̷�I�f����ݪ��Py���������w��|����:������:�rfT�����?|,u������쩺?I���@0Z4���"
�iQ� �tC�i[���Z�1x�� M�捙L>݀�t`�^�lL���*$
�.
�W-�6��Yoa֙Y��EZ%[Xr=�̣�;l���΍�X�b
ȃ;�-	�_�oԎ�?��]�Bq :�����6l��̥�I^ݦ�K�J-%D��m4PB7�[��O����x�>0>s�ze�L�F]��&�$�䓀O6egd�ob!��*� E��b�7	}3�����P(��(e���NC��Ҫ\ƨ���ͭ"�.�¨` ��᠊*���LAy��?-EK$��YC��R�m����^�v�
,�y�$؜�P \RUxUȧ6��b�5�rk�ĸ�B�����;�j�=2[�c+�j��J�a9���D�5��P�}������MA�_BF� y���
i��	�&P�P�pڵi�%t��nhftg=j?݇I��H�� ����ݚгqG䵝ə0F3��մ7
6#W��@~p2_1�EY�6[�1���֮.yn�m��Գ,�����_"������4���e����,o+m��ϥ��kf�71�mL߷��ߛϪb�`!Ty�U_������j�w��n��u��d+yZ�H��	Wu}5}��E���;����X�_�y�j��J��~<�@�?����_��Ɇ��['M�Ic�C��0o��Z�<���f����w/@$I�������o�إ����E��̆D�f�R����;DME^���l���P_Y�?��W��P}��ۺd�Do��x`q;!n����ڄ�KC�o��q�~��)�6�W�pi�� �k�	�(�P��Udppr��U����Fw��:�k�/l�XX���M���_���n�Y�����v �v���a��;��y�-�`ڍȬ��*��[������5N�C|{��A���߸*�n!9Ԍ��`�;�6{}�!ea���ŏ<�8L���U���@��뇫Ng����j]��Q�q3��B� �77�0��#��V.e�@���Ϫ�[xD��'vG�����4;?{N�=���(�e�H�r����G����UzE����me�/��������ќhrǙD,�V(�m[�f
[��o��r�Դ�O0����C�(����6ow��@�yU�:Q�*�)�(;7�ޫ>��31<3#�b$m�3T��)K�����c>�����$���8k���9]�6��mx�;�����#�UT�l��{2J���<�+�ױ�W�/�6��M���|D���(Eo�
��1x-��]�E��K5/�wR�q%E��$��ӆ")C��贴�K+i:q�"�i\��&O�����m�+��/)J���'��+X�Eҿx��k�Fڔ�`����c ��2�R��t4����������$�a�@h�RQ7���Q��۟�y$g�OkK8ľU<_��ZX �0Lp����[R[���ړR3�&�C�'��U�eo�2�:�]��=>���B묬�,�1���Zl��ui��~�6Ȑvg�ٌ��,�"C�C���������
������_I��3�(�K�f O�	�&���W�AŃ؇�6���q���g&�����2��辰�[CB��r�IwxA"|w�֟sfd�Y��v�����aS�3gzk����x������
����F>��/`W&�b������{�Z���p�ܚ�i9ޕ#_��Tg���I �u���܏x6�ȣ,��Bb�3wވ;p <WCS�H~b����݌xR�rj�C���4��]�bM0d_Z�Zfgwr��xǖ-s���£���]@[�ob�'+�;tl�8w$�Z�͎�8�o6����!�z� �+��� ;Y� �A3�Z����q�!���v����ғ�"o�I��Ԋl�_7nؕ��s���	�Kٍ"�*\R]�E�S=̩�;�O�&�V.��b���\|��U���t��g�ݕ��D3^��9�FK�`9�Hڕ���h�L�P�ڷ_<vf�w�9�ʜ�Mqv�F��k������T�Nt1��;<�Pi�����I�Tx����
'�!�M6_���Lq����\sw�*�U�f�'�N���{�Ivk5Jo-|�]�F5��+\ý��T������-7�m�n2`e�(SX�E(8��?ޑ�bN��c���ħ�)f�~�����4Yd�.��~���-󔊷|-��K�*}(���ii�*R�nK�̎Ō�������jt)u]��.;V��0r�*Բ��U�9��t�io����2����v@4���S�M>g���4=�˴�j
���霦A�j/a�A�	y'���	�����	�B�r�5~J%�J���A�j�#�%�yR=`���j�Z��j�Iu/fi%��z�͉(��0A��N(��ve���'�#. =��sٺF�C#\L�}V�a6�xp���i��=ɱ �i���X��&`�lOt��^Xt�m��Y���8�����o?�n�<=(dm�@<���`e�Ӛ�gZ7���	}�ϟs���&�ff���/|N��G�Y�0�5�|q>�ȱ������V��dH7Ӡ8ˤ��-���E� �E%�{'����t���W��g"S�=i|��O�<&��O���ə��_���AD]V�R�����,����Yd���?��ؗ~ �P^+�A��?- �-���7���mM�HS1�@��y^;0�ce������޽4�!!�-��gẰҍ�N�};;B�}	��Q\*�g���W����'��W�a;sx�2�-�P}׍��RNK����C8LS���ꜙb���!��J�� �e��2t2WS�����旁�bsCv�[Z��ȥ�X���ٟ���n�H|!�x�*_�
�]Ö�q�_P�(i�������$,�<"�~/!K��բ�_�_����C�}�\�ۺ9��wT�M�5�����@�W�N��B���=e;p�<�S�0z�,�o�5����bQ�v�|�s�]A�?��U�-�2)��\iѫh�\��N��z�UA벅������瓴M� C���g@?X?ه��~
N�.V��fy�k8���'T8˳���0w�*{�u,~gC�C��w�9s�G
d�
�g�T�d�g9��DG����ò�C���\?�Q=hь��c����0w����Y��z�a�kh<]턾�N�; 6���[��ނt�f0����(����󌤇v1�03[&�]���E��9���Ho҆\���h���V�f˕�����x7)�)��y��u$��ts�Ɨ��FQ�v�6�ً�\o='�̼�/�l��Z
>]ݧn]8|W]b��J&���)�kwp���sK6�6���V�R:Ս�cdT�'����D��6�9Oy`�� �]���%�����Y��N�W�h��ogh�9		���2��Nn�R��O�fQ������kz�Ef"ŷ��Rh�U��K *�d���М�X��#�����j.���7J.�	�k:Z�O'��?h/T'�����S��>.8�8AZYF��,��T@�N猙����h��G���OLd�Ep��N]�A�ҕ��z`KX�;՝2�K�nR�pNhK�E�>��4�	�۸�Ӽ��_9���ci?vO�j׉��z����u� c?�HP%�f�{_�&�!\����̽���9��^Z��O欧9��Q2Ni���W:�9o�OT���s�����wꝫψP�<�M�`�*`�|c�@�n���be6h��9xVV�L\;��r&�n�B�ŅN���g�@��5X�n@��ST��&$���>.��9||^�S�6,�"�[y|5{�s�gƝ��q�Wq4�ͦ��0��T�,�?յ{_־U�)�[*4�����v�e\�H�5Q���߶#&75YCF� K�J�bG)ׁh��Z�,�i:��u
�\
C�*%xP"����iۯ���>��#a���pw�����7y܎XM�h}����=?���uѷ�/�@����5�w� �Շ��dq���~��6?�̛eǽ�g_7ˏ�ׯ���8�^Y�B"S���8^y�4�� +q
�L�X䑜�s)0L�G$W)5���3w< pn��:����gq�-ݳ}䪾�51mr�>�Wc��!��1mS$��`=��������(�V
f&'�k'0ѢT�sj|��|}�"���?�B�v�/[�=	{������6�h���b'wIY��wnI�f�#IX`��i��`���O�X~�ܵ��lF�,��-�3A����8%~����F�~��������I7��`���+�m�j��#�R �t��:��V��Kf��L��3��A�9���Iv�r�_݀�*k�j:���"�J�5�����j#v�F%Kp����؈��Vڽ�Cê��IW�Y��q;P��7���>H�'I�A�~[V
���84��-%i�MTbpL������~��mu�MS�մ�������Gj���8��/l�GZ��S1�g�_Z�4�0�LC�'�o@]¾J��
x�w<�os��!'��?��斖$����NؤFn��ɭ�p�V�@���'nD�oЧ{ߏ�07/8	[��M��0�X�����f���	Yr�h a>l��F8�*.�mw&���-hcC�������;�X��T��pd
����<��\È?�-yݝSg�N��=�`D+����"y�{����ok��7��W��t��m�c���I�|ŷ8��i�R��&**{����I��_yf�6�r��:�ف3�ގ�Q����3i�i0Z�1�L[7�� ��D�;gT"�W
�)���'�}�@A���7n��Gv�1��B�
�F���N���b���_�B�NG5L�C�p娾�5%u����O_��
�����QO-O� �9�����/�^�mf�'����M�M���3��Cg�\d��OX�9��Í��#�����V6�tU�j�����9�T��V3|(�Ǡ�q��Hwg7q&ŧ��D����Q;�+pSgSc��f�}}�⁢�ax4P�,��P�C(��'>�C8�T�$�k��	�F~��@9�4/(��A��8w����7n;�ZB�����z�v�!��Iz�t�Lr?���$H�A�/�|�2��s�F|�Z��Sz��4`Dc�������'��i^_mj��Xs8�/�m�-Q��drZ�XC�9>#5"g-Hq������W(9p�W���z�4����P�9�
n���x���T�%1ZC!�Ձ�/yӗ0�O8�n�}>����1B�ڦ�|�� ���Ž��{�iG�c4��|��FAW���|<�ǹ_u���C����45�Oݗ��LM��}8�A���rQ���0������"\Nr!�k���k�绛��M�*�c��X��䗞�+"�zfeqf2_���bnN�\�tOgh�pM�������J�HB᪷�z���0��9x���`:�k�~݋y�����+k���sx����n�ب�֤�;��$$�oi�vWD)��6/�j�
�Ҹ'�R��!g�"�A	uk;�i[�#*א<�9q�)�L�>��DCx�֨��b�{/��e��dN��s0�UB��6�>���Z���OQ�m���>3%'��u��H�%
p���r�m�oi5�˾�A�0���;M��)�����sh��mN�2��?��ćиó6��נ���<��-� \���[����|P�@�޸w�?e�7d�(pղ������p+��;a\�P����y�����㲻�� ��0�� �m?��+�g�)�V���a����V�f8tr�s�����:�Wt��gՁ�}A���2#��+?��{��ni��cQk"݂�(Tv @���16`����`�.���y�qvl|,�ߤ�rŌ9�U��:��|��/����`|4��a�I{��V0=�x.�J_�c��.�Y�+��A��i ��1���v@�xTbG�m��Q�7�v��z��8���F�Yl�b1`��t�}�AX�Wb%Լ�C0���[ڥXjb"_�{3���R�����ZX"=X��K�s5��PP@�0ҋ���
_�s��W(��f�ὴ�X�q>O�~�!g�0m�swSn�}vAf�l��} ��z����%���Q��;i&Qv�߿�H���A�G}|�Z����_���<��\�>��:
�Z:�)̲�0B�t�N�V���.ˎ��z�ͯc5���l%m�,�&��3E`��,7���Cx:��Iǘp /_π���F�/G�]��WRv]�k�[Zvd���d���g�,G\�`�c+��P���m�5&Q&穳ީ<}�]xX�>�tW�,��j]�!D��_}L�R`��殂��%��f�����kï��$�ēL4�y{�-�.�'���?�+}�;6-hU���q��ب'��Xl%��D\8L����vj�9�+�*R�X�w@ t������ؤ��չ��JeZ��
�\rf/Zx0�:�{�w�<c��PREǉ�{4ܷ��N��g����|�j l)���Pc��L��f����\2��q�L�WK�����Pg�9
x�����BJ�n�6簗 ��xU%([G�`�Ţz���6�&�g"�nv��I��<]��_O�J�-S�QfY�l�/�
K\;�%H:��U+�QD�͈n�>��t�ll��f\U�};P�Z�W+�,��8�4�nT��As/�ݾ�O�g{ǁgv,n�g�u�����	Tp��������R:*�<.]�,Wy��b�f�o7�?����9��iu�b��W�otQ�.���e�>�(���4������k��F�m�-��Kx��Y��9���vBUrOiN��VZ��x��������S!c���8�_�M��#�}Dx̯t[V.H�����Y�n�]q�����M�k��H���Z��������d;%9P-�((�ܾ;|����\q�>���,�ȫ���>-}4 �,r~:�
K���$�f����80mѶXv_nH�nv6$���x����.�+q�j��j�J��A;���Y�	
����`�`Sf>��ǆb�Kۤ�6o39�kɦ	X��)*ui.�/�o5���b�b��C�jь�<����/�K�?�+�ރ%���=�B5�9�T��4㐴7[hK���8k6Po׊�� wٱ��1ut�.�S0���Rz�3^Ld��1�q���#v�-�7/�����g��e.v�U3�R�;`��"�-��cu�ͮ��WT�$����Lw�6������]�YZI�����i�z�݊)v���Y-W	�o�����$:Ty�b�;4Y�~}� Ň� ���9��~�ߡ��Jͱq*6�h�̞���>���1�����$ԓ+4�|��h��\����2���C�è�>�MП5�ּ�D�QÂȔ��2gA��Ǡ�^���g��"�q�]_��j�%@��3�����O%@��J��Z�W�t���@���F�~{�U��'،컡@u���UY���0����"}�z���v�-v��&�x-z>��(?�����ˊid7����c�e�,��)�L�,�������Lj��U��#l)�UIX�n�H��	p���#���p]��*RP�u-���'���(����QCE������	>����!�w�.=��im�����Uq���ń_�v��2��w�7�#[%��G�5�P'n9� z��F0�=-�p�����a�f4z���\��\�q>Z�d��sJ���D�2�,���+��)�F��{VBGM�,'P�� F�8K!�ޡ���3i����d�+hA5�U��F�s'�,�l�����y����\?h�IB@-x���8�[��\�?;D��HnH�ҜoܧZ�N���B�R��:�E����4`P�����{�Ê.ptdp��v��o����'43��a�*9;t�r$-���ޥ{����y}��=Q�V�D��{]�u�w���3�T�r��@���ipX�}�����
[�6�.��YQ�S�S��H��f=��kϽC3;:-�t����]��:CI�55�N��pw�A����o��'a�;u�����ǝ!��w8�#1��#W�&-���0�B��܃�:C_U�r�~p�~Y�Ǌ�6TU q��+u���\�/�$�j�sBW���Q�Tj�}#�b>����\@�T�X}g��on�"-�&t���~����� �
@[;w�ӷ�'{�"%-a��������*p�u��I`�|�P��ޞ�U�l>HT
��F���������ˎ�͇&z��V0;�G���19~o��jB�;�a3F�!@��h�p�TTû��|�6����	���W�O�J,;p �Ȥ�������iP?���.�y`'G���:���m��_���wf�-\��t�Dd������Jߒ>�(7���`m�d;x�Ր\��ww�kQs��9�B<*�oڧ�/ -�Ai��N����z�s�m>��$k���?��=��N�� u׶�<���s���g��ڟ*Jӎ"��@s�`���6�YU��2B>9�W��������eg�A�h�d��v����l���>`�ׯ[��+	T�z^��~���d�5.��^�3^��V`{0Y�x3�jXw�I:(�^B̥q uo��4l�E�����$f_!$��?(z�t��|���A~���C az�^[#NʳMz>�v�<�܃���\����o�&/��{�Δ�q� 
]{B���#a"�|7���\W�Z���E��	A �<b������P��M��
|ba�P����ǖ�60��w���̤�ױ��F} ����f<b��
&����#S&@*�h:�	����6ý�6�1�*#���v�$���\��Rҏ�<T͊�MQN4�e:�e�A�B� �����FA���!:�3��CCcAOq8��4�geDu��\��E;e��c��	p�����Vo;�T�KDЇ�n�]y�Q��|��j4����#̭�tª"�SQ�a���w��zq0^ǘD)va�`���P�k���9�^ܘ�Fa�N�/��N���p�:S�q�
�1�pvw��e
��0N\��J�7l��v�\k�MfƲn7�4 Ǯ�͈�b�n��6�g�uX�7��鯒'��o>>�n� R[���
C��ם��y]����x��Y����u����E��g�f��+�c� ��_���/d�T�Z�J֜�6���;�;�;ave��7�+�@��Y�~��� �m�)2qUK ���=��:�+�İ-�8p�uLH7/��y�Шo�H��$N��dK'*'���#��y��{hWPw!~�
�c�`��#S\��+j�QN;-���H���1Em�
��3Ǟ�r[�V~u�̽_�vxG�\�3P������⍝TT���V*lʦ�G�a�o�9(��:�*:��
B�;��Gq��<�Sț]~���i��*���s�*q�j�[u��D�8�v������$�n�S�*�Ӻ=٣��ȧ��^}��
�q¸/��H����p�_KkO�*)Q@��1�&�L�W{����x1�J���\���	8T���~���L�0�N+ḇ��z勴G�mXPj�Z�<�(v���*GB�p��ud�����H������������x�A���0�iO{
ļ,.�D��|���@�J��R�/���N�i�Nf�Ò��hgnk���a�*�-�!�.�wd9i/T�e�@oA\8d�ċ�������H��.�]�UI�Σj��8�6E�1ĕ�ۊF�#K���U��a[͝���"oow��5.�Dg���4�>�W�t��sƖnD�\^.YD�[�F�!���^	Q���n�cs���$�GÄ�9=�+��|��$���7�gȴ�l�m]ֻ($�T×�w:�����}D�2�_���`�V:NN�/��F�2{ˌ�e��5���4�15��o�)}1��qtI!K�ݐ�;9�F:\c�@����|�1b܍����Q{��:y�}0B��X\Q�!�s��By8�,J�����%i��g�aR=Uj PrKQ��srt�e�r��H���p62�'^�,�q��N�Ve�EStz}�ACZ�k=g������K�����u�]��w7~V�;��و�o�N�"�k�ŭ�����ŜR��/h�ן�t{i�5������<a���ow�W�j\��{�����{�ޏ�g���"���".�.��A_�b�x��'"c�����G�lQT_i�u[�k:�Ql.�i���־}�JL�������FA�d��Gt�B�y95��l�p�ڪc��l�?��;�ޕ"��_]L�6��V-qw��%4������>�79Zo�����o�T��	u9��FQ���>�yi=$�ӠT�ɻ�q'����ҍ�T��!{'6E��U�ዾ�_���M��Җ9��U-�~���ǳ��j�(�1���������j�\�9�[�D�vh�)�o�G�bg�E:�I���uF�h3��j�	�o��%���@�:6ZĔD�f�궡�S�_Õ�ܦ�8�۞���z����"43��e�^@\'�b#������o0З[/t`�8�U ����z��ߴ��A��l~M]�1�>*RaK������ƇG�rw��A~=�8wa�+J�S�2%a+�*̓�'�L:P���n�A�2�(����G5Eik�� ҭ�&�Y������yl�b�U*]HlYJgqX��XW�<�%�)��Os�*)��z�Y�V�|���z�K�F��LB�r0b]�%��/�~`��+�NƇ��+���U%9>�ư�4�Ң�8�Y�=��]"@�X�Y����N�_�/��ԝ����~F*��6;�qpАȰ�D��z}�������������P�E�n^��
~�ӏ$�A���$�?{��֌xL����cל���جSRq9\���8�Jd֐�H
u5�q���N��G��Լ�8'D<�fA�=�b<ͱ��a�^�}��jb������Z��.M9B�c>��_�F2_�uM��'fQy+���.,m��6�ġ���Y��<����rTm���XU\6ΰ�*���1�g��<%%�kv�4���������~���k}���e��%�����/�t�5���O��π�|�_�>W�VEpq��9���F\��UO�&<`��B�Ȅ�Ԙb���_�tt?���O�!�Ƙ�9�N���a[&7�_�Wj;�9���k�h�0U�̾�j��f��&޿��8�Oc2���*���1p������O�{�b��w23��R�������U��K��l��G��Γ���Ջ�(<}2G��pj/^��SAh��U+������d+0���!z�u�o,T�z��r�;����L��᜖c�o ֔.�^��]|�>s��̬��⭝l�;Nւ���^�o��e+�!l(�x��11��L�'$�nj�׸2zV�F�����ꮝ׀��A�b�fo6_F�d#��U��wie5Ե)=�7��AW�.7譔��D!�`��CcW���B�&����|}0���X��Eɐ�H5��Z�48���W�H@D��[s�;{K�T�k&:HX%�
^����=c���N#,� `, �}�gb�tԔ�O�m�z ,8<����Cf6�)A~;l��F����6�2�͏��q/�x`���^e�j��a�%o�~h�TyVJj?��6zN�2��S5�!ș��m�w����=��	T�q>oUo�����W�OG�8�����xi�d��gIgR�S������ٿ��ԊZ���ls���x?d��Js��v��j��z�Q���ո��>���n��@I!䃹��/-h�|s��BB�U�;��~��9h^�b�w5�p�w���NG�RX��1`��EeǇ��DD���kP	��}K��Ց8N���ͥ�+�a�����kp�4�0u�[�=o�'�����98�a����\��C�}���4 �z$J Z;j�������������Yo��H8}����5��c�k��������9QI������K�"�s�<sA�E�x�X�>��"[�v4��t+My=�����\/&�GL'�f�����{�`����N6Tg�|A��B#���:c�)@Y`��� xYŬ��D$��(���jk�j���¤�l#}�ʠ���D�|O��^�c�( �����a�d��KR�Q&H��9�������{���u�E��Ѿ�V��.B[���f&���5���_�U��S}�4�D�T�ߋ�_;Z�W'�s���C�rz�?����
= ��J@�e�w2Q]=���'Rs�u+8I�Ѩk��*	�D
�T5qfT1�(���|��Ϸr�ěO V�S�$����ːf&xr��;h|�i��q����I�utt�iF���Z�5O�XQ����� �	#� �I<5(r���@��'��h](�}yV��֜v��[�������^m#�1�b�x�?}a�E'�5�q�-@�Dob>��
̷�7e�F�F����ݜ!Ȧ	��O��p�DP�1���:��~�:�]Za�ʹ��J�v�KF+��d:��D�����eiK�E?��?T3�`$H��՝���"�P�jY��h����8�����)kk�g�V�u�e�_*��3����޼���=i)m���a�-442�Lb=��Hŝ�}��+ (����H��H�������sz��S�p�C9��DDXg5��m���n�Y��QK��%�����jͿAj��B�{_>fo�N�T��ֆ����գ��8�S۟���5���&�^���d �V
=J��n�/qUg#���uk����Y�夐O���ȥzN�\]��(����_c�@+xP�V��ޫv8w�7���?�땇�d䯙�h���%���uiQ}�
5�?�7u(e����;ź]��L����1�w�B�;y'�~p����8�'��l �j�)������4vl?�	X((,m�Z����^�_~��*e��a0��+ P�������H����̚}G|�`@���GN�t-�/T�N4�g"
;�L��z�����	� P�-�H���}B��-�\�_Sc`>����h饹*�A3����9&��i������A�y[&0��a�
(�'S;��ّ�g �f �8���p0���	 5�T5D%��c�� �.A�J��e'�Sl��*��P��D��R��wʅ�`��Å5��� �"䌾}�����#<��G�� Cuʳ	)�$ul="%��c-�>,��q�۫~����!�I�2��O�!��Z'�*������%�66�H1!�$����Nx�u��}���k�'䋎���e/ �x�k�}� �@=����Ϛ��m���ƣ�k�����w>x��L��|��!�VD�V�#."�OcŖ	t��	�j�(m�|l��������$t��Ӝ9�'
�k��]bOt�>F/,��ҁf����'��2�zB����!0]��;��:{����y��ȌXq��ola�������9χ�4��x/�}!�����K��)����l��0�r�]|��P�*�]���+6�G���)(���a�2��	}��<�3��j�ל���|$E?̻���R����N��f-�{Vᷖ⸛��ɞ�:5Edx�E� !��D�%�lo/c��*}���Ed�S-�j�#
���UB�j\O~>��h���#�ʤ]U��[��@)�[`u��&Ӏ��������%��2�ŗ"R��נK����Τ�G�;ckr��⇎G�Gn �<��R���P�������ݠ�B�f�7C�����cƑh�(🜐���0�x�,ܰJ(�Dj�����5{�.�
@�(�Jl�0hHlX�,G4��蕵�����2��>��|4���)_�-.��+v:Z��-ǲ����(�/�
�d*�Eǎ������Is�^����ʬ�h�k�G���!�R���i�V"������Zdf�:�j)���:��y�q-Lw�DR�]�щk�?s3Wʁ���lMN�\����%�Ʈ>+&7���g.87k�-֖Xn���B���|m�/>��ӻ��� \�J���������ŕUuX�=��-�����)o�47���-o�1.g9P�x��3�9�b�}��V<;S�i~�.�LH���~%�շO��K�a뮯�L���̅���A�G��"�+1�+����KQ����V��nv>�^^@����n2M]��6�@���he����d�"�G�_�T�]9J�߆7�����ʺ�om���|j��F;�=Ԍ�JR��|���g���
5hk�+h�$g�IOI��z�\m��BF���t�|��P��]�K`�4D@�i
h����ŷ��$���G 2��J����TC �Π�ů�6t�>�^3���*K�#������_�্/�_�l���r�K����@Y�,��3��#D�l�L��g�Ǧ!�.�r�a��Ϡh���J�����8���L��k�T��3P��sZ�I�%D�BTJ����.�_������5c)�8{�{��a[��9���Aƅ�^h��XGd�܏B��o�J���xg@	ՠ7wEl8}+!<����s�oױ�'�}0l�N�ޔv���s�}'������ׯ�G�ry
 ��@���c���x˱�;��_US��LhE�f{u����;�q��w��}�7��������<�d�ڏ��7�Y
�)�N+��7�B)i�6��-�J^�7c�?���Y��Ƣq��
tK
��[� )Ն�)(S�8Oq��?kkB�9��2dh� ��*d1�Gԕn�^��g�)d�	hL@�5y��%�J��}���l&ps�� {��D=�IGN91y�T_�s�n-�q��R��SNF���(�](+�:PB���n��[J'a3�|1y)ׁ]U�M���,���fN���a##�<����7�ȕ���\?I9�|_U�/�9io �9������]ƥ���q�� Z���ӭa>%]���'���W��DGw
�� 2�����;���ʛ8w�ٿeJN-&��9C��-$t�,G\�sy�¯\K�^��F���<+3�t_��҅Z�_紈%�7	n怖GHg6���|��}����T����7Փ�r,��� mx����m�D	Rk�i���w>��2 �����t�sv����_��@���J]��
r����.�}]������~�[��I�<_8�H����'�M����~'��a���c�L�����=�"H=^��������f��Ùr���p4�(ed:t��d�u�Zߪ���]8�Ԯ�G7��1������;���@�/0 ������XQE�fm+ÅZ�E�#?�\��k�������&��̔��9O}�Qt���%,�+��2'6�ش��ާ��Z�_�����K����?>AK�)�qL��vQ
��</Z"��G:�j"q�UhBB�C%వgmc� :����L�1./jh0�p�o����R/i��!C&�(���*�]Qk�~��9A���九,e=�z	�����c�oP���`g_*��j����. (*d��3�V�I���SE?%����!��9�\��x�p1_-�3����Ocf�}��J���@��>��
���zg J����� ��C`4��t#�gг�e@����l9 F% ]' ��!1�+ݑn�3�e�^�����x?�a��9E~�(d˩�RH�G3>hb��?�]Z��m1��3��薻�f$�A�dW�2�0	-�]�ۉ���rA���"��5��P�t�������Xd�F5 �b;*�(6�@��{l�����	E� >4�˰5���n����V�f���"Nd�����1�[J��E����z�R�X���ۏ�p�/�,�Y�K�Q��3�z@�z�)zL��?�U��}a������2}��u5���˚�#���[n9N���7,r�y��� G�?���U��CS�߷ �M��.��&Z�D��[k<o��п1	�.�W�~m\^~�r��܎9ԧ�T?�x@B�HB����\��@#A��Yz<A����?���s���ޤ�ѵ��{�a�)�띒��=��y�OfKo=����[�S��A�*�6��;x���j@�.cc���rd�1�s��'���ݬLFF��8�vn;�A�������	�x'������.x�w����|�%�K]a��4�D��.�oJ�)��K���ne��������չp�\�R�Y�/
��^ ���|�?��,�l���1T�VP��,�	,�q��M)�d3Ǫ'���S�P��;���V
{@#���wCV-�_����kOC[[��B�p�PՓg���w�Ԏ��X2��r<�������t�����,6Y��oCm���I����f�^E���o�=�
�UxW����A���eOKr���$Ȝ�ﳴp��S�T�?V���9ZC\���;α渐m?SP�"{��?f�]�;�.%�9��Od`q�zH@���Z�2���H�hk�����5� S�"^K���hiG��C�6�
+��I�Ѵ�_��1�(�yCY'���3�a,��(G�ɘR����+(�?����DI��}�jcO���U͖yF��-��������ݥ�����)��̗��և���Wg�r�JHL��󵘹�g��J����Wu�I���?�������qt���T+���\������zr��%�y~���z�]v��x��煋�!CbL���r�;B�����x��<-��`Д���L5��s�������4��w�6O6rRvR�(�\�M��[K\񺤦�Y�Jq��s�Vz S#�r����I�*JIu�`��E�6s�X�"Q�f��֯]t�����o8ui�r�:��oI}%��%�������Ck����o~�OW��7���21��5�0��<<ĭ���ґF����x�w���7��V��9�|w�~z!�������u� }a��h�A_��vG]��+�B�/j�Wc����7M�&#%Q�w���f�m����1'W�s׾�jz%E5M��Mq�/]J�>/ȵ��@=O��0�UU�ڥ;܉�oI���M���t��V��gYOTy�w����nńgؿ���U���=dh���_HjU�C\^��z�P����'����lĪKr�!���CCk����k���@)�PD�\t#���݈tI#���f�����A��\�{?~���w�������<���,Ŭ�� ��E6j#��%E���m7�8"O��;گ+�Q:��Ȫ2�6Df�R�����^gS�O�U6�����f3�m)zfr)�=�;JT�sƉ�>���N�F��h�o�t�B���	���1�s���Q����|T�(A:�K��Y�F�r���1�8���Q��`���[���<�#�҄��G*/C}���qS6*h���`���2nP�Z��O�V�c"��NOSF��
H�?�:[�Npt����4M�5�+Xu
(H.�Qr|�Y��ĉ��V�`���bPg�������?�y��ؤ�Vs��B\���%nw��6�(x�[���B�TF��`�?g�
^Έ�,���3%3("���J���Kuf���,o�#���Ģ��r4��oq�%}[�#�+�����|�M�F�4�Թ|T�a����/8�&��7`-���x}J.�}�h�����؃���f��)q�{�}���*ܐzPǜ��3�R�p�C�)��-Ng�?��~Mu69�4�oFfP������[�A�}�&�?�6$����s��|�n���\�W��������sx���A9FI���6(���R�?{_��/��\�ӂD�nA?_ؤ��/�����fGZ|ޔ�uf��ݏ�f����"�El�۳�t�k���@q��'e��E�s�B����$&,���g}�xٌlI{�����JM����C���u�1I���|�:J5�ɧf>>���ļ�����}y��DGǳ��\Eai*"�����֕!d_�~�?k!�P�\_��?o��lz�	-w7�ٜ�-��t�;tj��� j�<���Hu��b�����jW�����@+H<މt3_�Fw��'I��?Cq�M۵A�||X6�-V���C$��2���{��VJq�N�<_6pq��
n??��Ζy���ks�>�.5�S��L<=5
|���ж�[1�bcU��"�����^��3������W�T���]�w[C7Jmo,q��	��-GQ�f�)n�]�J��OW���W�K��ҡ��Wa������U�^A�6�h�ѹ�	8������i��.Eףd9���i?���țN�i�l��'SJĝ::)���i�,�N8�TXp���,�����=��_��N�'���1�3�(�A��;�16���D�c���_O|�K��t���b��6#��\]�i�T�&���9t��Z'[���p�o�UO.����[���J})؋���3�bv�q�!~��-�x��G�	��c�h7Z��Z���`|�=c�D��F1Xeǹ�>��&�&�ưh�6�x1�\Z��gvj7�k�]�$�H'\���\:�M���������Eޤx��*гDe��f�g�����f����g��7�u�6�J����
	�Ƭ�I�R�"�d����w"��]-U��g���e�֊�C�"I�Tg��m���zn��r�H��qsfQ�au;Sh~�:�=��HF:�<�	}���E����\h�Q���%��ų[��z6x�_G�qjv/�;-�	
8O����∬�".��y~;Q�m3��t�a8u�.m��Ԯ�gD\ `��A�Vmvw�~�,�r`<�ct	L�9�8B�o6����p��}�5F?��$����㽵�6I�DF�(/�����wW����3�̈K�?���D5�G���f��2剢+&?�yu�d���փ^�ꅑ�G�E'w���/E��LB:��~k�q��(�L]�M��t]�g�j�S̈́�1�4w��[}Pl�L�T�J*��l��Rӊu�@B3ЪQ��^�t��u,��O5�M$n�2x����'��1J��R$��ur��r�U�M-SO����M��&ے�O���l��@���"2"���Np���ǐ��
޾�ǵ�0����wv�#�V%������=v�9�Y�y�j���*�p�?T΂շ��/���*	��R����"���?�C-}F��)A��Jo���L�b>{�wCd?E���j��f��K��pY�8�C�"��px�wT <)b���OuU�s��Q����e�TՔ�J�%m����)�P�h���Е$0>�?\��|m�&���s)�BE����86�Sf���j��А�1���c�$ؿ��F���e?1 >P�=Ղ�[f��>&z߷l����|��q뿐�Ro��ȷ"t����G��ݔ��ϷX����>����.����.����.����aߠ���w�?�@Ng! ������	��������ƪ����0K�Jcc�[��p�s���-�2�@ �L!�r��+11���a�/5W��,����Ё�
��ƗHV�ժ�vt��
**Lvm꒒�����6�9
��ʬ��Ȼ\ll{�M�%d�����k�Z��K���Yt�E����zVm���;?G�T5���\�Z{���h~y9�����]�lR����G��", @BK+��8��s$G(�t��Ѩ��P�DY~>d1�:AK��U�K.��U�U}$�
ӂ�g��<��<v|nn����i5���p�@�9�Z���+�-�cUFa�����h�G�͒*,���P-�ِDR�c��6׋��t}�:�P��W)��\�"m��c�u����3�e�E����^��Ơ$ats�\K���R�V[50FPz��6�����'��'�y%�$H����||d3���o����l;�#=%���G������\/�����|ae~[��f���%fl��N�qu�Z��@ꡡ>{�"��o��b�z�"t(M�m�~��e<�ネ���IK���|ڛ�s�oL����V�������tW�z�+�o�;�gԢz�Rv	W^�Au�t}CN��`��֡!N�]$��Q�R>����U-r~�`22����!&��kc~n#ô��-��C;��*�7f���ӭ(&~�o���)1��Ɠ��,�w���./�Q�7�	�����밌q�#�����Qf�a�˅�V��v�#������_L����^GD�Q���Cϖ��f{�b�+$��1<�����Ĳ5$��"�z``��(t;�>��
)���MF8�Џ�n�O�%�\Lk��	ߌ��k���TV#!�"q��Z���-�ðlE�<BX�Sc�jվZ}�M|��z��XnC�-��Y�՚�ݫ��Ý��a��PQ֙~�	�o�!͌*iN{
�!!��q��ߣ���-�u�X���%��
���'�		����Uvo����!��ټ{'Eʃ�N+۶�k�s|I�)��'��\#����k��}K���Dڼ����ڃI$,%�s>��qI�������@xnm|���\hO��1�?���,@4I�%44QT��Vq��%�Ҝ�l��q�
5�!�4�,`�IxO��y��jf�c��5&����'y���l>x����#�S�<!�3��LR�����褽x�H]�
���Nۗ�DH���G�9�
���Zh����uv�~,�A-�he�bHoc/\,õdڇɭ8��y�	M�Ί͏E+�.9 �0�$��$�c<'���-0~ga\�	���<��k$$�m�؛�8"��=]KEY�����qh����<1>N���;��Vhh(�R|�1��8��շ����7G1M�E4G1Ȧ��l���\uj��G�5��z��z�� ����%6�'M~�煼��v�����q���ut(��~,�~�&K��j}}}���� 
�t7������^hJ���F
�YWV�Z��	�������lَe��6)��0~�HcSӠ����x������?��ʃ��S�����/ۜ���?�ۿ�Z�[)�hɔ�^�?YX�ґ81�\�"������+	��=X_��lh�O��_�ǱO9�����rՏ����7/$ۊ>?:��p��i��@w?����T����N,	���'*_Y!s��������<��Y��3�?aD#+))Y4���!�h}Y��i��'V�;}�矍��!L�8/�bG��A��Ǐfg��1Ȃ***�MLccc�-,����ero<+/+�ECC�[����F��)��r2�z/�����&�Ze�6��>�(&�Sv8%x�$i�4Q�4}�N,����O[������-X���'�� �_���,�[�㑱��|%D�1
FY��p���x���U�(��񱱥e���h
a�4=l����H6ICMS�n���̹.�vHݕ"sK1d���G�S��-چ������;�q�P(�fp<���y��ő?������z�$))	}p������O�~ϲ�	`*6�;^	��V-��<��C��T���@�E��6
��c$2U���%���+{�;:O����Δ���x���=>nC	���q�����������3�����S&��^(������JE��)9��=�+:��y� gE��/�Qu��j������"G��*vyg�|���hp��:k������B���������=�LyO�1�����j���%�h@[���3b���n������$����*+E߽k�Ȯ�2Ih��`bbj��t���CĘ^қ�����RP���5r<1A&��� U��Z��������߿����Ϸ�sIn���2��Z�i��yxxL�aP���@�sc8=_�S33B�ǡ�>���)I399顷	�J�+��}�VQ/��Xd�7�@�"�#��Ǥ��5�Q ��s{���bw���i��술弹����n8�HԷoߪ<��+Pwf���WFT�+��o^ y�Y�x:�~�^�v�:>���
���������pp��LYM���-������r���g��{��E�^��JF�qWS���� Lv��ήA�������A fOK���!�kE�.��t���D��*�;.f�)����|�(��h���'�㍝��t����/�η~�^�ALBB��~�^�L0%�`}����+�8�-�����m����,)�dS�s�#���_��Z�98n�8�0�H���O�'��.kXvL����{����f����nVۚu�z9���'���;+wm��G��A�A?���H��v����n[��5bg�2�o�G�!Y}x&����r�j�����.S���8-;����+�k~&h�^XWOOO,�A�ĳ��������%���^Wf�<�Y�?9�������=o�O+-ewqqI������v`���_Td�R�����MѷQ��G~֌���8[��.:�Z��oً��3
o��#A2vWx%/8%�N|@�UY/�LWYSj��Шit5e ?��\Xr��[wF����A��c�3w{��`�X륟�2���5���|@�hz� }s����.p�����lSѿhʓ�IF�a��ؙ�L��zzz�c`����w`��,��okk�HIK�{�7��1�x��]^�<YI�����V
�H�*��{����������R���6HJG�٘��)C�NcCf��uz�l���7����8���3��M�y-���Y�Hn^#22rZc�@B��R������%)�v�f#'�L��o*:��:+U9�!Qe�쭬
P�P8=dX�܎�DAAIol�i�Y���6�����g��J��	�:#mO�?��ZR��.d�qJ�������+͍�Q__����Ӈ� =��'O4���Pvh_[��[�<i�N��Ǹ<�٬��7��RY����`�pQ��*Kǥ������Đ���\[��_����6�a#�Tu�!���OZ$paD�d�p��3���CҪG�)Y�,sin�dhd��`��5ⴟ���ψ�
�I�Yr��Z��Pv�?P?�0Ր���{j�7&+���nn����]3P���}u��t�w��zO:�n|�Λ�a+�iMNM��2�7555�l��Q��(�IK3H���&�c�_&��W�XKқ'�n��6���4����4c�X�� 8�^��J�������{z�ޒ�.��,ܮ�H�&:�Mȁ@�\s�H�0�78�B��xp?���P��/q Fd9R��[�չ�(cb��@�YE؍ɇ[�9?��h��S���W�YoCA���!���NT�{��N�S��;��,���.Z[�[��K��ᥘ��p= �ON:~��T�%�r1J���. e����2���˙��$]zH��+.���t;���c##�߿?�?~,,*�ANS�Y Bm��>i	�y��\ `'v�qi<$�/4���Ru׾)�����G���}������S���q�G���;yڻ��4ȆΥ^~Y����s:�`6�%�~Yu����B"�@�����хiG�Ң:�j�$�+C��A[���ggg_;l�کT��x�*�+j6�������x���IQO��>�k�gӌ�t�\w���8��$�5�Ud	T���<h}��Q���r92�V��>���:��ڿ#ȍ���|���F,��N���r�蘘��)�5�ܗP.��F==����_�-���og��#=�@���jrp�,w���ea�o��E6{��"�j��?��Òn�&_�r��W�l���B���@H��w���ӸQ.---τ����������̵r�����K�\I��_�l<$���z��7W|b(H�nkru{��@}���.� �H���p��n���v�N���z���KGkQ>�$��ܐ�)���%��\_53*� .� ��$}��'�� ��ϝ�ʷt�M>;�J�47����XѦ�t��c��ՃM9o��@M?����w`�f�˫B�z��ug �Aٍסk�z��H��`"m�g�2�h����~`Lv�;��u�@�4X����r I����;�'�nv穵�S��Ĵ��e�5� ����慔j3�Yt�R.����"���sZ��o��ܸE��7׀�$$&����_$ƫ�O@��4��1�`mOO�=���=�Eב�s��%���(A��;:�h�XJ%999 �b7�����s.$[ۉ2AY儎ix�����z��sr8}4�P����,�1.$�Ԥ�l�O%��"�:.�~w�H	��u>_w:��=c�����pM�Rk����E�NUi��ޚ4R���ζ<�O~`V(G������\(䗗]�H7���%Owy�9�l�9�N{�S]�F�xf���)�g���4�[%�%&ݑ�K�ŐJpV�Y
�J��ڳ�g�g�%|��m2��S��H�Y����o�5���2�\Cv���D-���؋j�2n';H�Ж�g�D�����3&�p���!G�^I�2�ׯ�|��L�IMEv�iN�yi]�o��.��HpEEŦ/ �Z6��3��� ���������>̶��A �=��C������V�40K�蘙������U��}��GGG7W[K.�	�otG��c�'�Ǝ�C��������݊�0����K���8��� q�a8��{�:!��3���9�zi�cq򣮎T$�Mb=ڱؼ������Lv���-�_k�p3� ��� Ʃb��yGY^锡�#:VVQ]]J�)���/��57~������wS�睋a��All��;IF��>a��ؓ�!�[4��Ett(���t��}��c��������'0 `�YU�ͬ�|��@/3�c%%�b��w3.��@���P?kp �mo��f��ؿ�XH3��B�p[a��H�r�Ӄ}R���H^B$e��P���8V�j��ao�+�'^y	Q��N�q� ���FH PMK�7�D�լ�u7~���?�܏�٩$���h��&C���?���W��Կ@����G&;X�:2b��y��w���S��eݼf:�ߡ���X�^Y]L��]f�P��Ibjj�56?Ӡ�({(pvV۩�bo����R��b�m�⷏(����"��EQYy���p��e ����S�'x�^{��['m����	���nV�o�p����v�P�mm����ѱ������^g�p�0�w֘�Yc�����zr����aFv�(=�'C>>>ՙ4��ǧ���:e�Vf@`�;�I��e-��rź-������P����ʆ���~�O�3lo|/����P���l,M�\%�*��\���jn^^DRܮ���I��ྏ��!�HU��Z�����,���x���z����R�f݁}rv&���Q՜�|Z�_��"������m*g!⏀�w�4��>`,���92ǘ�$�GUU���,fl\�{�ʴ��^����	866�@�3I��9w���C�TQ�_��^ZZ���}�g�&$!imjB����i�n_/�9�����UO���	Y[]e���G��}�z��
�����G�Sd{D��z�T�
]儧Ň��R+W�������b�]�!.>~ZII$J![���du������A-�V���M-���o�u'�?��������cv�668�lP򪄸X�YϠ��� �j�)�[ή.������N�DEDx��8�˓RP��||n��f4�O`��xubqQ^J�;��G��'�oٽ�Z��h=�7���&'}��W^N��Z�m�1?e���Vr���AV?..����b/�~�~ʢ�P�>2�1)���N�
66<�����륨]"t�q`?��x�F��tt䪃����/6S\=$*-�{�I~YS�Y�m5)~�c���B �ڞ�j�i����q�d�U�������C�U�*̴|�+��P:�hݎ[QI)����A�k��yyh,*K|���-d�g���@��#���]�A��R4Yjjj�+����!����v�a�n���wVx�7����M�����&�n`���ʚ��~���;�Ӫo!j�o��ިEZ��Ԭ�`y*DO#�\kk�`�B�܎��%+�j*��3��~O������I;]JD2�(R��WNɫ��GGG�=O��\��I��E��Fks�%�4X�0��L4{�ik謡adD$��\"�dj�

:yo�s�"��'�7< �N�3�;
��%�����C"*��֌���8�����$�(��?�y@�*��QQ>55�kv5 �)�؏�"���q9֏�\���'��M�]$P�,%de>�v���d"�Z�u������-�����wl����X�!Guq�i	%K�O\�4��;s[���2�r*u~�K~�1������]��'�;�%4��iƅ���OXL����.���y��Q��+̆��Q'�h7�Z������5��ԿM�&y�28�K�9 @L���q�`59��7J&��{���$��ށ�"�UW����\l�Y�����R���@�����{�N��U6�����de='mGd�Ӝ���� tMט<����\���^$�HF�W�EY~Q&,Iiix2��פ�ޅ����_�P�z�p_�p仳Ѹ�O�-0�	�� ߜ���z��LMǯ�{VWa�Sw��9������Io���[`�x���nJ���F����"e��2��ϰ <���V�X8�ÍVJK��ԃZ�=���|�p� ��ΤS�w:�v���ʛ��Y#��h��f�C��Rϗ����Q�L�+���]�O��=,�z �3,O>~t:8[����%��k�:�VU���/�*Ef��+�+�(*�[a�Is;c�E��؍�/������mN���?�҃=~ힹ�P�"����r���/GI	*�S�������(*�v
==}s_O��Fzlpڻ��!!�I1z��g�M���Q��ee�F$?y.!���)@�]�o�Ci:���&�/$���넅9�ͻ	�q[����!��j��t�����ձ������$��'�P��B����x&zkO�2T�d����Kr��0�
(��)
�Ʉ/%������iن~�w�շ㿼���3XX�F94��ڀ���� �0<�.�i��r�'?;;�u�@o����U��z����Tt\kTl��fAN��TTJLܤ��`�lB*�">��" t��"�#���ߧ���m2V«k��E��I&�Fvff�^��*>"����߭�E���w|/��t�9�?�"�"��ьATǅ|/�8L���K ��de�����?�:j0�C�o���P!:�7��Lp&?�^�7И�^���8���,�/�+���G�y��� O�:
��/�q� /^#�f332����A�����L_�����o�;�u(h|�t2�1��вa73`F�א=
�-�HK.�V�]�\�]Y�3�p����΁�^�4о ����K++z@�����F,�o���R��J��AH�hEޜ�����ݽ�\ġ�&&�3�6/���y�ƪZ3H�}!T���@�!U�c���{�D���x��ІGG�rs�Ƥ�S(��8�k������y��ꕘ��s�n/��yiq���	s�f�A��@ڋ�ⓒ�̟G\O�><J�b�H������<�%6jSIII�Q?9�h��Q~��-��Ю��OH�NO�g�gF.�g|�n��X,(�"����x�A��û�;L8�����wN�ML�͵ciBU��0:�2@�-��͠��)\�U�39�u��oԄy��w�bUmm庄A��*���E,8�}2'�I�ig��Z�B�rwD\������]]�e�[���(r<�q$S{2�DC��aVRE�x�@�w���ۀ1������%%��=o��O>fҭo�*�&(P&*�m�8!��^��&(x�����A��H���҇���ts����E�D�`�����歚�9Z�(�y��l��VSS���������(���ԝR)�8Ԓ�o������U>Y]]��R���\;"�������ǫ��u��f�4J6��(}����o�	��y#���ӺRC�b7N�]�4��@Z�02�m�K}��>�X�O��!_6J���A�t���766t��8B��gTp���~Kא7����}�,��ۀ�Zm	!n�//-}�� ��-�̅T ��6O�,�Bv�Z`;��x�V�E c�`��z�C�u��`�0�Z[2�k��B�#�7��.Z��"_���y8rX�nfn'����׷��r�|�������W�{�����<jt?VC���>Q��l��s7����������v�u�9�yed��06��8��-�99��z��Xw?~L�¢LI	@01�4�����
m�f"d 5���m�c;��W��C����o�#���)�4x�����rtt�e���$��Q�Ĉ�ls	��RL,rw��_���(b�|����7��==@�@�t?�|��=Lxw�?��M���g��Xcc�*.��6x ˜��Ѕ��� <X�FR??�R��o 4ʷ�VV d~VVƱ9SK��C��I�����dQ�oh(b}϶�����"�K^�o�m�;x
���5**]�eJ$%--
hU���f/u��H?jim�I�C�-' 	}8�R/��u���:/��J�A]�}U\n'��US�]7����@q��&y
�"53���1`QV�O����z������+w�w���%T��=��Tì��� �2=1h!��v T(�i9(�_�$G]]`��������/� x��zi�Bh����mT'�9�U>�$+S�7P
��`��o�C��9���?MT=���`��kޮ�R[�Fd=���:tKa'6ټ��d�b���T�O��up�����e����)@�Qk�ka�<@D��/M)g��P�D���s:�t����E��t�� T��
�J��pk:����ײn��E�\^Fx�G�d�y�ί��7@���J��#{�Ally�����3u��}������}�B~���@��sM�w�����z���@��xv�t ��Zd�5w��zba`h��5d!�u�-�xz㉴̏�>ߍ����g�X�����*������Q�z����T3B�z�z��(�Z3X%�BBTTA���/j4�V�D \�C ^IX��<�=���??a�|o����"�
����%�|�RymM1�p������z�s�TՈ��39��?m�4�Z{����@{�fjߥ��b�(q��d��%��"��_�8�8|�r��J)3(�����o����0:yα��s��K��D)��JWM-��OP�=3K�����=C�"..5��tɟ��J�?��W��ځ|��L������`�:/+S�������_GzLD�dk��>�9����;��������~��QC8�����H�<����f����a2b��6���(���D؈)�TY��L�D\��H�F�2��I��P�%�����!+�L��R �Q�U�z�*�E��ݺ�����|�~~�b����J :�>����"�7o$W�.�6�J���<][ۉ	/&jG;E_p�p�x����� ��z{{y��d����%*��U�-O_����`é����ٚ��@�Q�&ѹ��i�8�..� �4YTƧm,K�H��(!��Yp�b6�:��tZ���e���(�n�!ˏ��4�e��_gn� �����u��yfʭr=B�y�������y��Ey&\[|ܦ�
��Nq�H��쑠1����t&�>��ϟ?�=á�_RZ
��Cj��Y��`f�z���v�v/$ M0o�eފ�SUG$/Onr���F�Q`E��6~����V�USSCG�1��>��ty�6>�����3555�<1���)��F�Ё����-J��? [�����)uKC�����X���"M��tQ*�_W��+�Þ@������WUS����1��� ����K�[ºt�30�~�{�D5#�A�����l�X�y�o��	cc���Z�ݡV���6�b򈁛�{5؞n��/^�H	ޙu9V��˹j������T+�����	sU����#�!a��jC]��}���EC�:MA-1� �\O�}�u�G���dde�>7��C�pq�@��ֲ֝�Y��U�.��
ׇp�{xǿ�Xp���Z6e5��Ym±��D�uxu������#���hC%aGº�����8S�TB�[Wr�=:���Ti�D�����;�qT�����
���¾.�US!P�� ʋ{2���zӗ��a=!!!����m:����^���z0g�\�x��na>hN����K���/��_�
��W������W�j�@���J����Y�Tt���Y$��;�hh�JJ�BȀ���eggzs��A��TtL���3\�Jf!Ê�m����Z]���i�(���9��;����t�9��>�('��u����꼞�/ �$f���=��z��=Rb%!��`N>a�����@`^���K/Q���"�rƐ�G���sI	9�@���J%���xv�!4��b�T�2㥇@,nag2���r���6�Y�?+�����>�,�aKx��L�;���I��/ �j\w�0�f���S�/e����Ӛ��~�����5l�5Pk0�`~�g���{r����?@�SNN�_�X��@�:��7���o�UϷb��*�|��>L�lN#DM��RƂ�fd�_	9y����=�|��ja`d�WU�j"�	fI-򅶼�~ƚ�G�����̳����?B١���g�I7@�l����zq�p-�z
�����`��p�=����:��V�	q���"��#^�9��m��E�M�ň�]ja�
��>�J��<��۷��wl-n(�y�&me��0*��Ǎ �?�8�>V�v؞Ωr���@ԙ�5( `�,9�se����.�:ff%J�gy�/���um��I=���y3�!`I.�=z�������� шCE@��AA����yRؤ'��׋�@�������YY��E�c���X{����7��l�����pm�u"�o��#��RC�6:l��UѺ�Ǐ�����2��@����	Yo�����r�Dv]�{����;����x����j�A���v��@�f��{�xS��А\�� �E(1N�H���.	:C�n���Fp��y�5�}��>p+�	w���8���~Y�������'� T�@����fc,�x��}�n�s�����>��NA���^VWz��k�TXZ:55�����P��Nryp��}�j�@���Z҄�yh$sk~��%�	�� ���B�z;�bg��	����qrUS����&_qi�{F}����;j` ��<|�Y�kxun.��~����`_&�9W9$�3�?����y*=Q�@��m�3C�!{�%��I2�I<���*
Z����+�22s���� �*2O�������WtC�(N�ܬ�#UZ�}�^@�=�)\f��r��OX���wT�8������{�S[t��ti��6����5k�Q�KH�@ ��D���|&\�Pˊ��
h�(�	���7WA����u�#�>�����f�l7I	z�� T%6 ���m*���hd��r����,"2����rӄ�<%66���\_aA>:ɘi9vc7����:1�u��&Њ���G?A9��6�N^~�J�(|�=�n��˗r������w;R��z���> ��C|kC]]}�4h$�=��1o��T�Rޗ�=���J��`������:U�''�QL �=�����b�<l��|�?�<;^�ffTi_��_-.�`��� �ٖ�D���3`-�It���Rbj�犡�T.q
��r��QSzVV���$��ً��'"X��d�t�b�_@م���ql�ݷO#lFx� ��\y 
?

B=��1#�M�����p�e�1�+�Ҋ�х�����x�_o�k��Vp2���x�yi�Og�)i��@]�vR�2L{�A��+-p>�	n��;���Z
����O�=�`�L��KJJ
�N�O
����9cZ�<���s��	d�ǿg} ��)C�)JČ�+��mu�*��2MUyt���0�?g�ſ����E�	���^�<���(�{~>:�i���iM�͙<�i�j���x����ۢ�Rk$8�O�WB1��OE�ZPE�t��{�k!��ԏ�|EJ�Q��Qz��{h$�����$�>������;��耴�����iI�����"@O�Ԕ����'ȗ���f\�Kh�,)�	�!ʊ_BIBE�k��} �'�u)��	s�r [�ro���ޚ�*��	�=umm�����w��fZ[��� ����㵊�Fw�(�x�'Zv����x����$�/�GFF�N�KL�s���{ ��-�WN�t:q�p��
��ɯ��ZÍ����æ����PC�5���||dp8\w�N-E��/��.Okڑk��DwX�7o�0�Pհ���EgǻelҌ���~�X����"!1�������|��w���P��o�����$�fP遝�[/�	�~�^��a�L�h8�d���	6�<���W漴�(��[.&OGN�[ ��ME`뚲Z���x���<x���nQAAA.��c֌��_0�VI�'u8ܜ%�,ېO��H����0(�����_�^s ���sI��z��x&�f:��Ƞ� 0�𲆬���k4��S��
��NWO.���~;����>Ej�����(N$��\2{H0}��Ë��^��~c�wCU��;;;#��h4�����{����h輸4���j�AL^3�����p33�݋+�0U�^x�E���}�7"�7���+�M��\~æ)�.��s��[_�Nw��w��	�bG�Ƶ<|���/�����)��?�Ϲ�-���:mV�T���M#:%L:3:��c��E����n��A��lo���Ę��22�i+�}N���Dt��~�?�©f~a��D��������E���wO��wXӏc�y�t=�����3:&F���k,�c8}���@Z&7:�<^2����hB5ϭ$�s��u/�W�<_��ښ=b<(�����ᑑ���(][
�S$Td�>9���*H���N6^�C�ӏ��������	�//D\$�����-#�@;'4��{JNM-p}���]o�v�Y{���$���{��u�3��.��N��o��-�p[q4YbccK9���ꇈ,2��ސb� ��2�
X�;Ӂ��J�S����R�������)����c�a��^##JU3�-��dZ���QS�1�����&Ɵ\������	�^py���* ��	+�V��)��/d��A_W������K*��nZ���r�-�|��4Wۮ&aݥ���|~�4.��{/dm�gI�v���־�?*凗߾�a		AZ�Ŝs.m8�۴��������c!�S�k�&������De����Lp��p��?���~�P�ٙ33���N��N��>77*e��	�e�8�LGg��V1H���;����sk���_�^t4.�y_鮫g,zzz7����\ZLY4��� uww���#y�� �a�S猱Ќ�B�4�%W�"u�j}�#�¼k�b�.����i�����}�`Q�mt=<���<�F�$WT8	�(����HQ?{�{S��Ӱq�!H7)�"�x�����ǭ4/��-4d+�$P��4��#�j�oII�>n�ȿ���jMk���c�a)��:��ȃ_$7Onz(O�%�;5^�s;7~���l6.._��W��F?K܎��A�"y5��5���OS�����뤾�j��m��j�_����2�dM�EG0��5{9&�#7o��p'aHKK�2�`x,�]D��ɓ�?Z~����Ƿ��ZV&B����;0�Q~AA�1�͓n�lCCC�:�+���w�E��#>Isr��70������mn��KF�Ή�>	���Q��ځG{p��u�%�H��;�%��E��ԓ�`JJJ��\<F��%��Ή-?M���
dBK;ȳ��|* Ⓔ���TJ;;;�Gtu�JfdR�����%$"j��d �ch;��������y��(�v��㏀�cy�3�]�������T<P��UU��j��=��-�/""R�Pf�	�W�i�] ������+7��\d���M���0l����kb�Q4l�zB"��ji���������/^�+��)�GL)�mƻ��0�"U��#���f⫘�M_Z^E��-�0g�	�.--u���!��LF !v �B|�jz� ����gp$��֗��*s��O��4,�6< Ff��CB�)�*:�ZQI)'�����%-;%))	�����H9:��ڋ�U{0
d��uڍռqQ��CFO�����?��=6@�U��oE\p~֞?7�)IA|p/,q���_ �s����$$#���?4\PU�۾*JK7HI#�J�t#R���������K���p��n.�����ctu�=�>�{��6���(?!�Ȫ�X�Z�v�T?�v׵}����Ā|�D�\h�ˠй?�<e����@*��h���"G�����5��g�^e��1�h\Jj*��D 3a���
�	/ٟb �=���l��F����CY�=��
1d�@�Q�I�*=.nn��4>�aI�T�Oe���d��ie7[���{��1��j6++Tx����~?�F����kKy�o�'���<�dڃ�o�D�/����-1�.e�?��ȀI075��V����ݵ�^T�`u�[l�G�5՛�=�j����!5x;�=��u �K2�V?e���v����5P��*�LrRܸO��ǥyns�wq�FQQQMO/� b�?H*$$$V�IQ�b����+�#_�Ȳ�pe��g��0��ŏ����i;Wd��^���5�����p�kVo�"d��-I���������FG5��Z?���0����f�4ZorXwx$�a��C���4b�E�n��
�H4O�TQf��ly[�����
����8V�ԇ��Gȗ%`:���E�7e[PZo�26����Le�w����rk0��9�G��75E--�))+�x�↬4T�W�,�X��'~�:�a�J����#x�'���RWW��7o�n�Gl�tt�����z�Q	�7=���j����V
P�����п=� P[��gdt���:^��m�տ�gP�P������$�9���K�Y�x��]ͦ�A��`���3�G�������Ԑ��Mi[�"*�I���y�~���}���XN��꺒3�G~��<R5�[�Q3�}z6\�g�`��f����K6�w�+����n��IY}�b��W����6��ũ����DEc���|�B�������3�cޟ��p�Y6]�������$:�O�>@�66�+++賓����GU�����_N�ۥP2z�\I���%���h�X��[n�[nt<<π�W�ބI�/..�쟺������gAc06��p�+��}["�7�vr�%(yttD�j��<p,D�-\%�1���E�Y�Ik�r�A�Esomm-�~J)V�$Z(�5$��J_?�[L,ȩ ����^�L8���3��Ȉ]/���D^K�&r;�[��,A�̞��69��A!�R�<���I��-�;8\��&�T6�?w���dW��f&(AsVC����j�똸8s{{LoooR��3O�X93�qp"�`�#�1W8⡴�����L~ޗU.r�xxx��� �cB/�s������p�<�G��ݟU�`,�&ҷ���J��I�;��pv%K^�=��`��᫷oɶ����|�T�1Y��$i��v�~�s��"7�}�Ӈ͝��*�DZ�E˄IW9 �mmmM�Ξߏu.�v�+{�2d%��7wf��	�B;�:��^瑃ܮ��RVV6��j� 
����Ps����,��F�y����xVu(�G^�:��~���_�A�ɖ���:� N���G��j�#,8��!��v"L��^�~��ʚ;��(�3m����qT��l����ކq��܍��N`TQ����a���;
�U��b���������dѹ���ݥ�8]��y:�L�o@tQoU�@v���F����`h---z�g�X;;;^���*���+5�ה�H�.��7�r!�x�y3��e��C��a�����a��\݁߆��1�J?�����o�"E ���������5ɨ��:�x9��^��������.t��"�?U����;>9і�^�&�\`~��&(*�W�Ẍ́����ˡPP-�ˠ�����D�n�S�x�P��I  ���)�<l����~v>��{���=�ݩ��*�K$\MMM�)�}-��`:��w`V��n&��p�df���q>��|�H���R�������zY���J_ד{6WW�l=l(���� g���{bI$���_h�6t0>���)�^��n��01;.w�/�F�מ�`�.LYRZ�dE� x��
���ykK��8�#�v�ڴ��bw�N�#4�WP��j}ccY]]d��;A��>	�m|h����9���}"�81h�?[6��n��>Gn�OJz�U�������$������O�*82r3�0�9klK8����
�TKoY�#�0�;1�0/���2��&��TP:� �fnF�Y����[l����S��RD'�$����G��k<����u��gMa���!hI��

��DLP� 0���0�y���='���uCq#�zƧ��>;;s�PW$Q�N�i��i5�;�J��'tB�C��(�V|/�edeß|2��&����k�T�.6�m�/hC��gR@��5�Gn>��<���DnY��~O@D$���M���w3BB�J��Xx^W0��A�C��������^�d�T@�@T����3��f�N���N�I�!�J���q�%o|!��g~���d��f�d��U�����W������3��O�$nB*�@S��J��DYp�=IJ|ɛT��7�p�z�,��B�G����>(�m}���)lll�V�n�&��:���� |�@<������Ƶ��"\pxE	�|�D������ʣQC��XX$����mǨ�1���@�1[��������:L�����-~T`;�]+Mzik*���WKV�0���`�r~v1�ȶ�����d]c�x�:�i;���;-�#B�#T{�����m�����-^��7q&��XL�%�u_�#RLD�I�i������{�b����)���H��4�g�����T� ���.��=���}_���=9�ʢ؝�z�T1~~��"���������5L���xAH�ڜ��{д�<���?qdp�H�+�C��Hx4��F`S;�U����;�t�H��*;�휁��9ƛ7m� W�i�x�J��V��WԪ~02��5v��]�3I���[_�i�2(��������$p�M8���\v�K,y�$'��ǆ7���{�)
�qKdqq��%����}\�;�TZ�;~6��<Ƞ �m_�b�O)��#��l��ɟ?��&��[|k�A�� =��m�G�l�יm��8��{��vt"�xY�����p�#�`�����]Ҿ~���&m_������'-���5Q�����k�y��D�Ӻ$��ْ�/��+���h��X8-",(��ʭ�w%D�3Ӓ����ş*�'� �YXXd�3su����؊���y�E}�&!"2����҉Y�L�t���J����qsq5�p����J�ʬ�"��n#���Cx��e�����<����a�3�-4Cy�%&����ݘ�un���a�&���������E��P�ʺ���y_�2uiok��kx��M��5;��e���#�d��O�8�9�h.��ք�-�t��}ɛ��p�	' �UwO1�C����ʓ�`��47t]�<֕�����t����ɍ��D�1�K��(��A�ֶ���r���S�v��,?lS���έ�TXqw���+q�2��O���a.�hY�GVG���?~�hbd���S�c��(���.�X�gr���V_[{���f�����}Ȍ�r7�w�<��Cq�9��~�ךW�G�s���R,y��������ɥ����򨙾P���z	*�u�7�Қ��^���!��D�{�
z�z@Wc�Ax����H��S��أX,������8�R �,q��e�vO�\5w���^M�����_�� =�t��yyCy��ػw��**(�F�E�m�/cR������G�3�M1m��Eb�'k��A��R��º�����.\W��A����is]Q�%���`��ߤÇOt������VB�����ә��E�y��]�F�<=�tfa,���
������]�l~�C]���S���KA?䑫Ȁ��{�
7,2��$�x�?_ X��Ȍ$"&v��6��s-��~���eu-�d��{i'q�'���H5g�dR���U�Hhl�ML$����	��sh,1!!��@��[��b͢ʟ�U؆/(��=��v�d���/��~�ՠщ�b���[�j̡�o`��xo9R'�\.j�"?�72F �7�����E����=��l�f�ð�`�����IiCg���� |�;�QW���̏_<y�=�ۚ��WY�M':8܇poD睂����ʣ�S7�rB�bhQ�u�d��dd������¹[9M�)50j�0\>H �P�X�vU����f&*&�g8ȏ������ ���=���V񷢸�� ���G��!��spp��Po�Di�7E���� �����VWA�G�t�a�d��"��-���0�����_�Ze��W�-��'���S)G��G@���#�QB^g�xb���B"�
����ڻ����}�{�I�pr���Vu�y��+�tn�K�rQH<�X�?����/K��Jx�6a�+�+��@	tc�#_m��:9P���.ox��τߪ�}�$;;;?�۹F��a�pQI�;�6��7/v�z�d�b��=[s����z�����0�Z!�����)�G���%��Î�a�ɵ-]��Z�ih�Yk���
j98���2lcf� ���2!�Y�M�H0�VZ�E�奤��y���A���}��8����v��Cs�q�DU4�r�=�*���n�?_ER+���iL��?U��oۘ���f_�{QR���b�����w�r������[U�7�c�Q���sgd�l����΅~��%��~d�/(�}NG�RSS�QY[OȏwU[�����y[��}y�,���-n�� ��j�WQQ���,FGղ��-%922*���E���I�dIJ�aؾ6��\l��aH������|>�yE��g&�����A6�� g�(�`���i�u�u=�������!/����W���R�\����՟X5ʢ��Tj�,/�l���q�U s�'�C�yY������!*�D�#���mHH��6����^�[�=�p��N���@S�G�,�?�A��C�!�����6k�JVN�se��(
(��)��^���wE�2��B����>1�����0=���7W
��_��!��>>>�3���:��GO_�u򕃌`�||�p��l���1�c=9�۹]�������錿ԋ��'p�ih�*[�UUU���T��J*!�
>��x�e��kI*0�ԟ������Ioo��v���\��5%�����8�c�j
���K3�U�o(<z�H��0W/  �<~xkO�J��0�,,�����h��4��3Ԕ���zv\-�f]C���.bf����f�em-�����%����򖖖��h\{?���g1̸苃�<�s��u𝹹�i�����dip'B��UVc#Sr�@�h-�T��+h��� N�0~�L]t�h|8*�n������E�)h�rg���q�����W��������?���8 ��ݵ��)�:��x�k�Ve��C
`�M��3���G�=�c�o,�����Ur�)��@/N��ɗ{�W�������U�+!*ڢ�4Ր�`��|/��	n����[��/]�J�4����+:���xz�k�q2��J�1O�*_⭓��/F�}����-l�#�@feXQ�Z~م��r�������;�S��wO���CPAw�)�srr����6�gg�*����;�;��&���W���J���u�G�M�4���/���1���_�ѯ��3t6�nTV�W���<�k�����e�{�%��i)����-�j����_vDW�<�^h�����������K�'�7�7Q��>ZU�S�l5�� ��RuM�3Cz�>�`O4
}��xM���>0>E�����o���Ρ���X�̑?�Oǂ)���L�GZ03�P��1S5h���,-�\]G�p����:��͛li�jz�~��D�g��3��_�1T߳|����#�8��g'lbC�j�����յ�i���@���|��n;^XLjff�_���k0C����Fq��tu -)%o�����$6�E�(8/��g}��v�#�;
G�Uo����̋4�u����O���ݤ��)����*��	쟪��5�d�)�_�^Oo�S�	��كhȵ�ښr\����I�����s��**�La�_)))���X��<<�@���wl		gՋ�z�<F1g�yq���Oȶ���w�! �X׈���ǹ��z��+��?J|d;V���d���~�#�c�+�����m�K�C����%��{(��L֮	���j�g[���/��D_��>B����*�A*L�z{;ШM�K�G��YYy��r�Q��:je	�ijŌ��r����q����a�regF�����1E��z`jl��Tr�������p�7����Q�0V�����U�UY�9���פ^�Dz�N�ҲZ�F��W�l�i��fEH��P��v��^W}XSdN�0fE��^�M}G:b��y��_�'�1m8"����Ā)�ǄN�e*,�;�n����@UQlv�&���݂�W�P�n��0�o�%)��G�d��_DV̾[XP���v &&��2�9�v�z�u�)'�d0��m��v`���)5���V�԰X�p�[K��Rc_�E*~������ʡ��%���M�,�$��T�}Ђ�>>4�Q[?�:r!�t�]������w��6��xWS���sf���	'U���ł@��A��ׯ_�(tt.�=�|77��Œo�_m����)�j��t��K7G�~���\�l���K��V�	���ۍhD��֚(�5�\���Խ�c��c�����[^��<N�,���AiOc,�JNI�|��TaqwKR@Ψ!�� �=(�cʹ����T8N),,4FY@�!n>�j�"!��V|�M�f���P�6���Vd�@mʉ�{��Q�������[?%\<���׊T\�Dj�$ǜ���PaX�{>�\O4��VQNF����䤿�G�`�#�ϟ?����˒�֣&�dd�!h#��r6��ZZ(�}$l.y���:i�֍��o�vp��QQ�u�wI"\��5��>�l%q�r�w����n�L��Z���L�G��Þ��)p2��6�����A�w��^A$��oj
����50�<�
Y^6G���W���9Dd���rW�o�,h�������c�/.���{����I���g��1��Fk6�����
��:`�np�߬�i�DmǩwZ�s*�a�A.��틎�N��2j���Q*�~y[���X�8S��T�$ȑp��R�2/i��lDZ�W�&�Y��s�G��A6N�ҡ/�h���75��{ק����
��5�5TT`?%������}���a�W���"�MXDĤJ���l�f�n�	F������j�U��3Yi֩gZ3ۚ�-��[�	����_������Dɰ�c��"��,؞�� VuM<���ඳ�ϚkJ�}XEW�*,+�񱶶��{�۸���c��������&��ů�|�
�LLG&w��GM�g�6�;�y�p�D��QVF�c�|�ڇ}
"*��iU�0��i*��$ee���x�	]�1�ޞ������^���(U��I{9 �GDɵ{�g���vmo��?|ͭ�M�sꊷ3���N�^)�GE5N����S_����c 4)�k�������M5�$���+�b�IϤ-��gH|!9%e��AK�\���r#G�4�90��RF�6��:�#s-����-�m�>��V{fA�о���8��(U��}w��fI)���0�[x�s���E�/_ű:rX���᝝�.v�H��^r"��y~��ɰ���������[>Z�q������	U���|�|�����?�]��SP֗�����*�!�J/d:�׭Z<7R+�����Nӭ[����ik#�����;W^��{!P�j�����߿,��x���D��k����������ꩧ�-[-R<!~X���͹�A�N=�=����W��%#}]|�\3��zN��O����N����a-��g���/�ߠxxYoA��>��Ņl�mc٘��aE�<�D[;��S23����M�S�Z7��h���}�wI��@^|�(�>��z�E��KXx{�UI�
�è)��n"I�����ݏ'�Ţ��5D�Ҹ��3@̇�w[�-WFN<Ol,�����]<|a7?�I2U�&����&�ĩ322(.Ex��*VBp���*�u�g"�GY.�q��7���	�L9����:,,�WzW�є"z0�]�DbF��f�g�w�Z���~M���p�gD�JKq���Q@pp��QE��^;y��:�~*͝��vˏY0����҇��ez7Pb��T�g��'�m��7\�C�b�Ɨ�!8�!lo���u+m��Z�s^E����ߐT�Þ�`��|W_k.��>��\I�Gt��EG�g�)%ԏ���>���7��o�����'eT(�wm�����ZY�����A���_	0)��%�&;;R22���Q!L�ڄ��o�̓!Dm0eu�t������(8�D�`>���
2!	h(^U��[�+�3��FS�#��p=�}�[�o�ў�s�g!A��4�H� �s:�+`*:��2��$�7Ե��� ��@G���Җ11���U��B6t�����{|r��P��F��x�d�o��K�IH�Խ�#8?���2X~Xf>�2E�7h��<�]g%==+�����I���R����J%H���u-؋����&Jj�<港e�J�X�jq�6����61�b,�cn���|p7v���8�_+��t����v.i��.~!�a�<6�j��;㖳d���[(jl�����鏩��b��l�����B%ڥ��!吷�&;r�ލ+&���,~�<�X�!��6y����b3���n��ؤ�ސ�߰v53Z ��^�o�t��ْ��wgZ0�.��gv���3�[o��i
����{\j��#�F�w(c�C~��eT쐐��C%xZ�f�mAu>���j�Cnߨ�v��P
q�b�WW���>�k��W�R��������>/�#�7̙q��U���{ji�/^\ �~�����_���9�B�'�??xu��̼L�K-i�a���V���Ts��aģ�~��Wt �8����H��/� �NXI��*z�K�4���}o_7�bUw�㢢��h\�#j�~X=.�ZҢ�ݖ���ݰ���(v}�*3/�������/	"��E0'��6�c�X�����c'���5?���Sd	s���Yj>��e~�،b��A��4f�"����9.�ᐮ�vX�
r�WI�|��<c��='Q�ѐ6f�<���=��3���X�_䕃�N�ӡ�:lmVC'K�3N�L4�-�L&,,,��;:�/DB��=n���S��n���KHM������@FZ�ϛ]���J,<n6���Xr`榸�l�%ѥ���4�����X��c��7�r�Aq�#¥"F�E�Y�DLշ9�����F~`��z:hSU	u7
�QSsbRׯp��yG'@݊���vtT�ͨ�_���;���&�Uq�nOr&	����g+��R9Zs+������d�m�D�7U�$�*)+�����Ω}e "]p�]x{�{��6�����kk'�|^�TVJzbk�W��_����5�79Q�*3��(h��A�˫��9랗��m;Y/޵]�fҙ�>{Ȕ��l��z��e�ZZ��焁����V׎��DR��Ƌ�ˁ�nY99nq�O�06]˓7���Q�,H�M�*�E8�Z�@����77G�����[[kj�T���s���Ԑ�Z/�B�em������s��C1��Z��S#��n�e_�H/��%��1�t)ZFL:�O4���}��X�zŐ�<(�P���[*��%�\[���Q
��#��@HG��=�YJ2i�������5��+%%�5�TLM^G�����G�fW>�T�#��zxof�a��I������G�\�h
�h��&�ж},]Z�Υ�q?	��B�+ .�Cڨ���0&(7>�J�P��VI���� ���z���=��6������y���p&_=�C�@�pE~�J�M����Н������Z\�c�j[>nn����&GgkR�����}���2R'�2# "B��� �&6>��������l�4)[79�x��NEwx���7կ_/w��C̔�	���U���~W[EV��ϙ3���Tcn}w�%%�Yb������be��Q/�́؉�%Xj)�;���y�G�M�>0��||�������Ю����4\\\AoR9H?���?�������aq���9���ZI���*K��F��ҕ����כ	T�q��!�	!m����FFF?���n����褰*�J�5ũq��I�(z`��K������9Þ�9����s9܌����:::�pv1�ǔ��]h3p(ڣ�����T_K�<eB���/��e���R-�P=��9;+�7SO��]9�r�)<�J,
$��p~�Vc�F^^��3�3���?/Un/�E��?r�Ƭo��FPu��8�h�-�JA�����ndz:��IX:_=T����\R3:�Cf66iKK�����>	�P��T]� ��߀&F�GAڸ�E�Oa����a7́�k�
?��w��be �El��	��s��?m�JA��uXq�%A%�ma�I$~xCJW75��J�r��$7ҝ�D�N�4�N�I���X��qp���~�+v������aLF ƫ1^�Q���KsE�I1�I��j����$f.�Æ��q�TZZ*���"-��ȋ�����)-ljd�j8����d}�r�w9cۓ�(dx�u�q����D�{����,>`U�A�� � #�6�WZ��˗/ߪ����� � ��[��Th�khHFA��M/��MF8p���}�����P
�d�%�������-�\p���Wt	�n���_]����{s�#��;UQ�a�j쳵L�Ճٜ��qKJJ(<ѝ����[CM�߾]�?�
���
� k9/�����$$Į������׉����y#�����]`�e�)z4AoRM�5"]7�)	Y�K�7^;v-��}II�&H���	��Ļ�*v��k������%<�Ӎ���;� �1䊆��eA�+q|_H�5t��_ث��t��w�f��ݭ�~�}{��G8���ެ,
䩐����%AɎONr�6ra�负��B@Q������-9�H�+))���q�����K<�W�|f\D�ۣ:��D��x�_�A�9nw��^Y�=�&~w�&������m�j�[��a�(+"��9x�4����4٤�n[-ǵм��^��#/5`YRR�xyyi(������G�����J��� ���g��qQhkE*'��l+�>OeǨ��>}���n�)}ҵk�
~&�]\t���b�b���Ė�;ԏ���׮	X��O�9��+Ϡ�������&�ąVB��O��LL����A�<��p(?�X�s���Qy����7Dd�H�?�B'�wX& Ņ)#��c�VS=��ֶq��Gy^��抝�r 
S�����hM��vq�*�a��;�vBB¸O���ڱό9�ů	��L��sp|�H���	���2�50P76�3��w�����VV'O���@u8��PE�m�ػ�Ra�u�Ŋ�()-���JT���iEcc�?�� �@fǻۋ�6�W+�g^�����jj����W���i��6��Q,�M)��zm��V��r�b�AX{����Ʃ������ܔFLlR^3���_�0����/J2�לQU��a��wz&���G�w�����>�5�_�0�!��y�d�Đ����O����G(��~���YfC�0�s5���YY����Y[��ф���'iy<��U�л���_A~�n��H�>cJ\�C��1�Jv(O�g��,{ێ)�ˋ�?9N�wa�Zڷd8xi�ȀAh|�j��,!�"�Oumm7ww��m�l�Oj������<ϖ�9��o�w�yT6��b����U�È��f��p�yU�����y�G"gT�Rs�N=i3�-3sv�Y��
�3ss��k���nG�=�͞���#ќ0//@�䡸�YKa>���}���r�X,���_��݊�g��r!��_�41Y�A��Օ����_���y�Z�ݭ߽��9"Vl+82�1M"�X�!-8���}�_��׵����������\g9;8Hl�,xWu>�ts�oi�G����aI��KxuĆVX;���u�3;�Y���ڞ�g`�pT�-8Z�G�vD�.S$h���f�m @b�b���3��[����m���Uf� _X��f3Bg`��7Wj��~_	\|�z��~�̓@�;Ȯ�˨�����5����Å�i����Znp��*��\!6�'���H'��u0CW� �O�9(�ku����4�&&1�,{�N/��(͢o��b�UB�%�=�R��|�l���_�w�~_�����$�p0�z�e�E���Ϋ�Q� �#Qh62�%�4ՔVz"��8r鯮ȡ�z��O@<���z����>ɯ������"�"%��TTH����tSs�����w%+j�ql�y�Edb?������r��ZS�_⮟����Գ@�޴�[P,����-?qj�q��A��m��yc�b.���Ӿ_�Q<�a�Ů��V��))����.��>��lW�[^�Cr~��D�7@T,��}����`��WsI2��F5�#�C��$�ŋ�X6�*=7�|�Y0V*.��hw^^_�O�וj�0t%98��5�\��9��-O�:�NY{�����F�6θ1�866�a�nFMWW`%���Tg�$�D�[�f�5�4{��+C	�����R-�	?����z���%�{����`:I�='����I�L�T�����:ۜms[#`CCC=��*��� �>�2RQ���S^�WX��k� X�q
x��ظ�cf�/��k(3ƻUџ�(��Tzɢ�ݱ�e<�z� �z��O��-j+%�.�v���c�T�k�:|�<�(^Տܿ��0���"����p���^0�c��?8|X��Ҿ��͘�=Q8����^� n[�X��>(�,ָb��4�������<�����]W���&
�e��VV/q�YM梀�1i0�]K��/M8�,�D�869��7�E�(��z����G�T����k\���|���j��\{�wH!�w�� f3៿�����ŅB�cbHP)��q?��/�ѥ�ݔ�����xW���w���@ʓ.ȳ(j|�ۓY��'���ߎ��ntS�bR;�9��*Ɋuw��hIM��Yx��lnzu�g<^MR�z&y�pu��ߗ�'�L����򳼽(����[��UZ]��r�6*�v�G�c��K�e��a<�&��U��9���Oƒ�0�T�������s����n��h,��(� �a;M����(>��}�^#� ��Gσƙ�pQ`��׭��؜~��ڼ�	plu��YQ�;��࿪)S��Y�⒐�(%{���8ZY�9���>�ݙ*���M�H06?>����m;����h2�7stՅ��O������~��v����K��Ʀ�7�ܺ�,��bN����4��dD�\8����<fUǹ&�l[1���8a����,!� ��Gj9F��Ue��6ic��dr��s;N����l{X������%��2���	����&���vD�E<]z��0�u�ں�ұX޻�
��|�LW��Y��S�R!Q�t��a,��Ǉ3��5t|��}ǒX�"�p�{(#�EȊ$@9e�C�H�z±��^��Sz.~m>�#!�˨��Y�Й-���m6x��a"�Q�r�Bh��wb�����U�ߵ��B�Ѕ^὆�q@���U��{����Ӵ� 	�u�����4��§��Z��?=c���I�}�?�1��=..��������^�P�@|v�z�{|*���dΕ�D����߸��ɭq466�
��S���T�l��ip=��Cs�`c��Q��1 )�B�Ʃ*9�d����3-��M��9�T���My�CC�.�]�c��ia����}P�o�j�zqݷ�n5>��o�9������R�B�B�t����		����B��蜱�)�����lX�<��� ����H5f�V_�w:`�5r��G9%%���{-u�`��Ǆ<��­6x�wWp��5�k6_#^o+��KF������`��Vo����g ]C�q�����1�<�� ZORP�m&��j?�*��ݎ|�5D�Շ0���`���ŁN:'f�05��f����M*�������SXD��]A܈�����_!KĚdzIo��KA���R�~.j���фX�t$OF��\fG����@�-�u�I�p������||�W��@lc������t.���-��B�j���$�LL�^��-K��S욃%c�B�Q��
��U/��jI��]F����Gˁ�+� �;�R���Wı�+J�=	�EdqҸ�şU%��a�M����{7�sX2Rjk)�3�(ۮ�jSg�%,����~u-_��ЃA˗��}��}y�e���(�<����#�pY��e�s��M��N�mM��"���ܣ�d{�!���w�������H�'r���YD-��҇��;��NMSs���1یp��l��ݧ�Ka�,��N�4�R?��^ј�0���jP�����.Z�Ș�iլ��)��vþ��t�~?�|W��g �|��1-
9y���1�<�b�b9��v��O�f�MQ(_���m<�J�W�зriQj��O��Ed��rtA�8��v��z.�H�}�����C�K�������O�6/Xx0s0O^/�NLX��SB��a�K0*�������o��G��=��[�������b�?Y*p�s�r��mG������+�v���w�Ɲ+���$�f�ۑf����M ����>[|�A�B���RAÝ������v�V3�[��<nC�Nu)��m�rYi���c�:!�&乼`����W�+���C���y*p�A#-m>1ȶ����U��}0�+	�u3ː�d�����@ގ�sI�i�1������������+��^��f��}G����ZZ����P�K��wTBn`�MA�Gݝ�Z��]�����q
��ɓ��Hv����c���l�b_ڬ��:�����|n�嵯5bC�D�W�%�x�M����*p]I'u��g�**y�a/�����Z�����0��In�ž��t$ddմy�OQCV�5�P�Oֺ�t�ŋ�<w{�gl����5�,��&��@ )�
4�k�����{r���H cSE&_|k3pG�89+It#�{upYQQ_�gG����e�Le�h�i�c#��eF�D��K6L�ȣ?�Һ�~�[<��~-`"1l5b�~P�&�mkU�hg�g�S �2SSOq��$8n�2�v��x�⿬��`\�щ�$3A�t���3�	-
�a$��׹�������[9�<Z_�(����:X��[@�_�馕�}ɽԸ�5��Er�t>�ut�p��NNN>21�8纒��T}�F�)C��C��\�0��Q�%���Z�� H�W-L4ekeJ��2P&7�EH�4�#����a����>��ɬ��*�U�&�)�����8�
���{$mQQR�tozJ��9�"*�kI^U{�:�aB!�a�p/D�r+�=3���Ǖ����3�^����,�>���$`�M��b����+���T+__n>K��� �*a"�H���gAK��c�1�9X��雒�@8�Vuҗ��m�hjk���&d�ƈG����&ߊ���^��HF�ފo0kKR�W�޽��8����IM��WWD�EQt�?�������%��l�͍_�qkFK�<QOO�^�{��x�wKxn�#�/eIi'�y��ϱyN͌���B���	�j�ͥ�������*M�^-��N�|�rk�@�Әm���UK[��W����Ι���a������[� %��4�c��H�*�J�vU�5���hw7�,ȡ����ܜ|����U����罎(<�!ф�^{Ur	t�چ�o��)� �£�K�����mkD~���i���x�ﶷ�f��'��fM�������LJ^g��ࠢ�j[�\\�vjJ�9��w+��V�WU�D�Pӆo����������{��I3��f-��+�w&��L�IH���xYՕ1�?�|3�5��G�s!6��}Վ���0v��q��ꚭ�8����l�q��n�ZR���Ũ�<��I&܍�_vm��R�]5)T���*��ۜ���<h��s��{{\��G7��4�ex5���C��93j�m��/�����)��9��T&��ʐ�M��e����{)�As�]�Z!az�VRb>Um	��2�<��O+��2�G�������5�y`���u�%�U�$E�䜜��U�(j��$�ɐ4�K����K폂��`t��l�w�R�
\��x���i���J�#c��s�@W��!W�֓Ehy\��F�8(�6,�E2�Wrf�C��c���y#�)l��&/؋[ZD���>�Ge�^M[��b��r�E%(�R��Dc� ��]���b�K~x����S��� *�	�$Q�㱢R�s�p[{����R�ŋ�%$��.}zf���A��sGsN���Y�E��& ff�2�(���rߵ�f����y�n��?�߅��/��5�NqI��g�'��o� {{{���2�3�T*�^�y���%8���hZ��5�V�l�RQ�#�Gm`� k}�N����{h�j�׫y�\��5z�Q;泐'a��-�yT�TUፏ����ͼ=�:^#���
����*g�g)�S�oon
� ��l��`��M_�����
"Hwww�,��%��!����]��-�J#���{��}r]�Ù繟;�������]�wJp{��!~0�{a6`�0���m���q�H;s����x��6�_r�Md�ah�8FGE)����qTU�(.�wYm�����k\�ap۸]���9�{�+&�7f���5�h����i����,)�ۋ^k��R����i���NX$g����	�!��m�^��c�1��}dw~�zdOV��RHH�U�I��88�MM�)m�T} ��>ݼ��s~�>=�mњ���_׈���"��:�S���	�� �Ư�߳�����:�/�c���$���U�Yq���!�Җ)d����%4l7[e���u������@��ڑC&NwC�]LLLK����hn��7��B8cbv혙�k�{
������v��V�xQ�9	P�>�R;�?8`A�E�	�hv�'��(�5nw5j>��HK&�(2�[Ո�bLZ�l}m�MC�KR�(�� 3�b?���l o�Y�BS��K�7�����nN�U\�= �ӿ=��K�2�#?���:[,JkcuތP��f�tj�m���.�yz�!e;ꙃ�K}����j�zt������%�Z������N\\(�g0���.��h�8ت8(I�����C�6���0�3��b�y��J5�"�2{�
M4�("9rOScdd��s��n6�w���V
�)���%D�Y����kd�>`�Y����s�*U�2<�#��B��@�d$q��^�i��ʥ�����h��E�	�Vm�N>���@�%,,J�-�@���D�j���|�0{�>C�O"��gd�y�O�\	��;�������e4N9��21q�v��G����-{C��/m��������Q.��Y`u�x�Ӵ�(��o�h&���cc��|�3��Zg�ߋ��̤W����Fk3�
�|ii�𝽎��Q�[X 0F{��	-/���֩jڐ��6f�b�n76y0癫'����-YQ�����8�1�%���0���t�)0�ɾ�0R��חd�f��F��c�5�����]��/���C�fs~PI����?w�w�(Oۙ�ꡩ�}}�ł�� ������ɤb�H?'D�|��(�Sn��*3��q��Yc�#2*/|��Ѭ�tAj!��#�2��ɰ�_F��D��;�)�u�RQE_os*0�:jf�%��%]9��p��۷px<�3�����&C����ݡ�'����L���/���[���wx�G�]lN.��j&s`q"�|�l��h�5�-�^��,��t.f�K��֝�N��.f�`��<zzz���Pqqx>�������r���s��M�Ge�Mj�����v�� |yݧ�_i�6�ڐ����[��e6�L'*��b�~��9$N�ع�0Ѐ��Wf�
���U|�n���`�P�o�-
�R��x�Ƚl᷊V��z�G��g�
��G�Hn}/n�V���5N)�s���|D����׷&�{e���T��% :�������D�`����L���)HSJ��&��4-ߘ$Qo��>N�Ih�Po༶_k�~��ۃ�~2X${8,_������,�a{rv(��?bAu���a��.�~[��(V-�����RR��^�ݥ 9��QE�=�H�8m�CЏ�=�g�?�΄w�#455�(i��3Оɧ2���\o�;�e��K�)�ZS�h���(}����9f`�����0���b�e��v��L~ssj5}kF!�N�;�]��a$�Of�r�T�ukE�8j���TI�������>��N��y���
ו}��V�fW0���e��/O��9~���������(КU�Sk�Xg�H]f�d� �?�k����7�g`=�f$��Ņh�R<_o��m4=ž�c���>���do�\�3Q�+W§]�����Z�h1�SX@K�ꁛz��\�`�!={���>e�. -������5�����p��c��b&�s; �aaa{]Pă�Pg��o_�i�G�_\�z���Ej<� �a�.�<}p�A���ѵ��;�5ѭo��b��^V�'��!N�) �1�,��U�z/;��4��7
o����{��s�؝��ۯ�*�w/���E���c'M��w����m{�킞�&5���Kq��Y/�ئf��J�֜�c��N��m*o֘�[f��BRRZ'���A�z���G�j]�v�ج�B�o�ߒ�>��pqŷ|�geRi�{#]��|���tٖCB�rLŋ�'U�W(�x�5�~�x@��3`^�����@�Fܺ�s9��Ѐq'�3�\jcMEp���׆��S�`�t:S���P4��Q�?;B�3�@ǡ��� b�x�DRD�����]�����Bؤ����m����5�=�n*��3�g3QIUdU㑒�Pf�λ�n0����F�_R�Zme{�dz����Q��J����!MD(ۑ���D <��� H��&�=��_���zEȴL���嬍��5�����h᪠����$�:�#��Q�Ph�������C���{@�U+̓pD2�^����v̝���V����Su$�/냜�sT��8u�~�8�:�L�L�[,Qr�	5��8rL�ʁ�R~K4�fZ�;��Vٺ?�����w*���&k�ח��*��b��'�,�e��i;�bBaK�л�Ku=��I���S�lI�<l��k�TD�%2fO8�+�-y��Xە����G���,4.f��ei,C�v������H��v�5j
_�e��x��Ec��100x��z�	>w~��WDh�5	N�7�i���#��lrZ�����B�FVG�ߥ�lpqp'W~�E�0S�1�wZ�lcpA�'\|>=,��������h|��膻����뚃�j�)!8̿�6���Z��
*��'��7���L�>�߁=�?9��]F/�i��k_])���1�qk[[
�L�v�"������9>�<�݇^���i�������l��$�UID�րO&�;��b��B=�MMM����D��0v����e���c��h�'����:�3��5z�h]���U�:�V��&k�p�,����*+��<+qs/���#A㛰�C�w�uŏh�k>��H�x��?���r�quu����;�<�t�:P������%��7WC&q+s��VC*���3��k+�PUi�)��9���v�����"�ƃ�݆�i���2�f����~u$�m�\̺�;?��~K����µ�y؏�:p��H����QuO������j<|z��L��_���륍�6��R���r����D�!v=滠��ۯe�g�2F|�h��̾y��))&���RY""�^��HQ(ss�M�#vr�泇����FU�������p�<Y�AVG����g�a�Z���\�$��,�F�E�%�;�o�6:���o��SXU�����~��Q�?�p�����O��?B��D��7���-�*�x��M6{�����a�����a�������*����N�E^�;�>d��p2a�F}j[/c�&���<::*���>2�@����P1�+�ˢ4�q�d_밂�"��R�3��pV�E`.�&):�
����b�w�������8�`�H�/�����)���Qs.���G:�J��
;��4���B6��i����0	*Bv����r��۴�M��K����--�+l�-x�Y���
 b]�-���7���t0��=�n����>���PAa�3j�EN�h���?��tN����s����{�����u9yy�M8L75�Cob�x��BMw9���/�G��1p�K�b�2#�>>VS��ǭ	���r���SRz36�}h�7��v8�+��A����|�t�ds=�Ã䳾�H⟡���������l��Ќ.k�6TTD�[q��<j��,[9t�u$�CC�3q��Y����8��v�)��P�˰��OY�4ޱ�v��VVʍI��i���tǢ_3���Q�u�^2M7�Dyxx�_bnFM����ң>��}��vkz�|�
 ,�-͔�ZQmou��oUIS���E�?}_.C�t�7D$��˲��W�dw�ӭ� ���S [�mr)Nz�^	�gV;���U��}�sl����(�zA��� o�Po�P�k�A��������Xe��S岍����Y�0k�qdˎ�c���1� Z���5ǡ�k��u�x�#nE;��aC�~�(&|�K#-m*�#�_���r�����WvS9� �	eJ�M����E�)�MMb����s����H.�;s#����y$^q�@�9�
r7��ꍘp(7�t]q�v9wS�4��mث��Tw���%\eT�5��%��o>�?��.s�-rPC3�F[Vzѐ�˄7��kb�\Q����ؘ}�ԛ-g<�B���"�^\��Cso�|�4(b ^ݰ���jT����"4��Ν�&��g�+h�D�%�"pD�<�L��]S2ҹT�H����H�7�vy��*�H�㤊�]9oP�`�5ȍR�����Ҩ>f�.3�3���6� I�^Tқ-C�e:�<�(pz ��{Q�8g�ۈ�h���uPa�r=�9`YX�7����g�xW��:��R�eB���=����j+�z�HN��\~��>���L� 䰸��s����9��0���M�P��`B�r�ʶai0	Y��W)�#*#��D���Iʓ�<�W�9�5Ct�'��;k����;;����vhx�pm�@LV�C���<���
��blP~�}Ž����{l,��0���Չnm�V?�ƪ��R�zZ��!�T4�Va��j6��E����g���_ODNv{�t�S����zQ�g,�.�!A��U��e��5j�+F�Mޚ@����8��\���	1 �u��:��|�S��ad�wۏN&C�*^�4�b,��@�v�ȝi�ڌ"e�ͅ/���ȱ1��%���l�n��0k/;Ftd�5��%①�=��-��|�jȽ����j厃�z	��x�����
�e��\����Tfn��US�:A:J�(��:~��D 7�N��-���2ω��T�N��D8]O"	10Q�b��~{�EK��(W2�!���U�����_�%g����P�~_����w8o�FM��ޕk�������9�y�*K�n/�����<�6|���_��ϯ	�	��-� �~�p[
y�5�;%��Q�*CRx�g��?���	.}?�`�6��Oo���̺1b�J�x9�6N�	[��lTYn�5�-k�� F��_�+���@8�k_���p��n�Ø����KM!͡���K��⚦%�H���K�4|�.Y��,ML�;�jQ��2*�d�e[�L41�hj�`l�.1,'���4zl�ÿ�i�sP�!��6?o���p���5z����1n�4B��j��۫!@o
Mk<r��Y��6�陘��=�5/�mX��w\l�I��EeJ��픘J9��[�m�DP��O�-�����ts���핟i�(Ù$I8-v�l���{5T&�P
��"]v������9n�^�F)&���?+�G��?X]!�>��Vi���k�̢�B�edD>ή2$ ��$��-K��1�j����{#g�Kj���ʅ��LRS�7m�x~�c� �IՓ�6N&�sp�(B�(T��>��Rn?L���xG����65��7��bO��Bg�	�m~"n)b��|%�DDȸ�܁�,9՟G6��׶����	2`%���m-^�F�qn	�����'q�l��~�lE����!�.Y�2���pYn壩y�����x�䚈��	3I[ق�?(�)C�+��6�
Kc�U������oz���Դ~����x�4a�sŊ��E���0K>"�ҩE�:!�T�� ��T�{j>�z������M�{�_��	��ȠG0�AP22"�cs.h�s
�<1Td�Cl�#?6��+�1y�[ݓ�~��}���1�y��UOf]���W����>���W�G,k�C�Լ��.)<�s�B?X��<�e�H�4 ���FF����� O���X�0v���b�8�]�M�/UW�����o�j�7^}�K۪�\ZQ�{Kh�p����Uu��'�2�mzkL]G�Ӹ��m�D��d ��*�䏗^��S�����&`��Y�����i���<9,�>0����F)�]����mSI��k��m����m�L���dcg���@O�P(k@��� ���;W&��ݡO�9��ECz���Y���F��A^�k���z�U0J�?����6NvQ������M�b7�@L��+.�3����m�ђtҸ�㺦$<�SEtf�FpDU6�v�l*���e��-.����,�J�dPy,�h�Թ��k_N\�=&k�3�W9�χ���W�Bh�CWސ����3)����S�FoCKQ0�ǙgG��Ŧ���KJ��v�f�544�<�&�@�s{���NΦa��ww���1@tYc�	��yK�W�8]M��]� �tFlB]_x�A�[ʄ��m��px7�<��#��ɱ�X!n�Q%j���e���,b���dz�sA��ؗ1��|Rr��������O���1w��Pm�>n
�@�P�;"Ƣ��K�O�n%bۙ�?��\;s� �=��w�4���cat~�v�0X��C9�~�*�cN��ۢ�����b?��F�ֆ[s��z�X\ۧj �@уѢ�ބ��ޮ�o<����������=zbTpK̵�gϙc|\bK���(�W4]�ܥ%�NȪ��.t��&h/|�����q�\���%�}�.K{�۩)�����̪H���)��ǀ��]7r;m�t'jw��\f�u�`27�u�#��_"�&W��p�.�);���P~;Wm���U=HM7�l��GLl�Hђ�����v�n?'r�U�X��6��V��}9�Fkc����j�.ښ�+{Δ�w/�}$�;�����]x�����OK��]<6�
���8Aniw�m��0���8�f3��L���N���Sj��]b��Pl�6��g�L[z��u>��n���!=eXM�x
}���ଢ�Xe{k������z��&�D���c&]�^����f����n]������@���U��c����$�*�H��7�.n�,}�ē`�Ɣ}'��� �'M��9��= b1c��ym��K�*�ۓ	kgU�໥V�j[H�
v��+4�X����Z6)&�י�B1���)�m�7�y��Ŧ�e���_�=�j��v��P��y��UȽʹ?����3��*'[�IJ�]=^ǚ<E�U���Ԉ��=Fߔ�K���\������4���o�?��U�݈�[�E\��0�_�`��jEۘ����:�M0���"���n�@�)3�y4�����]�{M��^Eg]]]�馔��>��"�8D���۷k����_c����W>���ר���p����l������Հ(��ґ�k�%�O��(�"g���tt�
�%�}�y���>���\sv����X���*�@WĹ\�\{�Kɩ�bR��*(�rwoUcMO@鴦E�:���޷c���n��d�0��W��To[�-��V�kO�m��a_F���ϰ���Z���?,#��-�� ���8�̗=_6�ٱ}���t��;���+GGl*�N%�u�\r�A���Q����ݩyyN�t��Jδ"�
$�C�W�|�1IP�׽=����-�3�_�Ҵ���]Δ�d��4!�?�$V^iRʎsK�U�sy�hS�������mQ��)??��ɜ�G�V�̬��Z����}�,
SU�!�4�t�7�\j8D'ֵ�������iZà�S�
4(���onX���X���L��{�c��׷_Z�cG����&�'SDt���oM)��TA�1�&��B�����I?N��ޚ+���N\K!RF{M�:bviP�~��b��"�W����&��Ɓ�*׾�+S�簊0!����]hh���9A>�%5��zFh�Ju�ࠣ��3H��&%޹:��(.މ9��9�((qlĦM���2V��H���週�?�]��]5��x�R����o>a����5�]u|�uZLI��A����b`�{�&x�9�zjc�MW��J�F969I��ʹƔ^����Q.�t��I���I�W��	��p(M���T�� Z���m�4S0R�M6�U��y��;4#b�T�v�g,}���?�ih�m���!�-�����m����4��v7Ŵ(���8k0hy�z�z��U�<��fl�r�N����m1D kH��4��{)����v%��\r,һj-��4��l�>����]6dG�3��&�G�ݛ%P�N%�t��)}����"@e�O�o���ܭaΰ܀:E�E4ꅻ!�����<�S+���N����d.�^����W�a��C!f-�q�Pߒ��ʑ�i������D���������Ke(6n�:u-"H��� -M٠�#.Ȍ�߃�n��"�y�w��rX�����$}�QlNV�ӯ)�&��b�9lĹ��͓�ѡ��>�nJ����Jk�%�>`�|����#�k�����0�^�7�4Gc���n�f��ף ��>n�����
r{�P�R�n���1_}{=y���l`G�&�\�4�l�e��*��	�H!pړ�3	���4f��x'<�;���m��X�S>��։(U���l(\b�7�05������.�p]�����x\�Zz�&j*�j��a�ɑE�|Ä��#e���{f^�E�YUC�׏�xq�Q.��s&Bo�����hÈ��=`��gff� x<�9�r�E&3ͣ'Q׳�X���RF�~�b�??`��8�F&��>�[���-��;o�
Z�c�m��m��m#D%itW�s�C��7�O��P0���ѓ��M�5j�8H$������(**�g���'���S���I� �#�Ine�r�/�fZb�t7<M�TUE�Q�I�1竩�[����:��XhS���YE��O����9'�4'��+bAW�~�*��T
��Sn�i�5ay�(�]�6��}��0�����hx�4��.����L�X��� �^�[�拐޽��:�����ϟ�2>*q�%��zz�b��4�ѡ�$���ܝL��S �y�,��W��N�w���ƯA����)B�>B$6��K_sI)L�ٽ��6�G���*�ga�3hQG��s�֑�.�����	�?���ҕ���}��*Q�|u�N�+��FT�B�'rt��%���b�A�ovp4.�w���6-5���V"�^���+���y\,���N��O�<*8�ǻ�'�WA�������'z���n��}R[�f�Q
~4mcG ༰��XG�U٬,/�#Ϝ(���?�`4���1/N>V���!���)����k ϳ����F��-ボ�=VH?�ѻ0CP�MS�M5���rN���<\y����\?��9j�ޅnO@�k?�2h5�RR�R��+D� �<#c�i�x�_�a�}�
��=��:;����Ι�N�r����}A�;3ӗ;���x�A%$�)��T~�'#p�`1��!��4�����H�+�m;�@EK��0��z��!-�N��E�^��~�m���eiCF�ǵA��5ǧ8���%�/���U�g�XrK����SЕ��~�����9�^��~Kv�!ں�Y똘� +N_J��`����& P[G׵8�8��+��!�/�g����.�����c��x��^;�\�.�M=�&��U��j��6�I��w��]��3>�;GG%�i".rB��?��y�?���8����������B�^�䮜���}ݩo�S"�-aD�.���xiD�u#��}�t%fj��E�w6Ǥ��vC�e�����>%S	��Q-�}��� 4���=̦�&��#E�GOo!ff���%��yd}$$�d�a�	��WSS+>�����z$��Mz۳C�Q�[��6
��>t<��r���:zT�=
~~|]]����K��#�*=�����z�^����~�,3g�5���љ��������#'-a�ϰ=4g͚�1�f���JO�RT'�uu�nmQQ�;9=mfb�l�eT|j
?ˌ�-��Zg�,��5�MѰb����������Ŷ�\���'�z(�B�=��U�\'^��a�G'4L��CJJ��h��%��4V��)#�o͕�����r��_��{|���R�j�y�M��,��=�@}���Q�_�K�آR��6sg��A~كD�*��{m�٠�_�ib�����w�PD������_�Uڵ�pp�����_o�p���;~JW��� V3̎���*���:�NLJ��q��r�=�ӿZA��?H[O�VJ`��}l�[B"T-�Q����������̬���q�-�"u`�y}}�	i�����4jH�E��9G�<�6���
�������L���D�D�ĕ��闚���m�-�y��^ȑ}��������ǹ-y6��;��}�U}������=�q�TT�����Z�1�3�=ηo�W���***��8�*�:�{݂e��,��V�19��.�����{^�̲\ke%���9���K�Z�R...%=�htrjȑ�$w}��R��sOɖ��>�cJ_������D���!�bN;Q�!���2;$|DfY�^�볻�yˊ��Q���@���}5#�����B�R�༥%ƣ��y+�dZqDī��",h~��r0�&����@ꮻ���\E�9++kؚ#/e	6�@e�g<'�;(����L^S�h�g:5��I��"�z���c�����ׯ_'$&�J��:��K�)*Q,�	/�8��K���}ww�<�[G_�c����t�<�Oٹ7�HoG���p�6�ϴ��C�K�����==y8884�/|�����<�Ҿ"��%1.|�J���HO�Wq�OB⋫�˹�S=�35-�R4����ƒ������~l�1��auu�������~�Ϥ�z�6$^��ƙPF!/%��!P<RR^�􊷲�(��� O�'�ir�O<B��|��枭�����!k��`�II2�������ZXA
r>=���1����۱ �!�fM�
޺�Kǘ��/U}yxBU�̡<C��^%�r����;l��������III�n�(����t?�E�)
���k�q	��?$��1G�(@OT�;LQC�M\^^�y��MEM�cp�sL=�J7��R����`����4;�g6f�?��ЗO<�SR*R��������/�����@u��t`��1u����.҄��%z�q[f���[W��Q����6����z�Ij�˃�Mr��q���?�a6�SD�F"Hj��2��Kv�����r��os����=����Ҳ2���ǝ$�E��HQ'�4��rzF����gWyG�S^E�Q�N#'����?V���M��І�*At���_O���z��$��HffS��|�r7xH�ʫ��0���ޫ[��WA�7,w��4�=h��jV/u��Z_͏��B��<;���זz�p!�"B��m*::�P)FJ<d�i�(��p$�Et��d\㓐��)�--+So�:���~��ax�)�5���v���,����^���V�=<Mӳ�8�	w,�����e�4�[V�HAw?���#HG������g}+)9R��.ATֈ��NН�[�i+ ��V�����mRҀ?&{�!�8H!$��qH��k+�FSW��c/�DC�(�/��Q��<�J���] ȭX�p�Xp�in�*�R���;����԰d��)L�*9n�'�#��'?�*� �Y<����,��I6���U%ϦÈ(&T�>+MX[ė@�9���Y��WNjx�t��}� �o��Q�&V���]��]((��C����ݾ�#�W�<C���_̀�.�>��BY���m�@F/��Jx��VsXT䬨������^���eŨeG�6{G�f�c�
iUmma���[�Zs�5o!zz����鉉wF�����
[������ש991���+K� �)jzec����,�1�W��N�o�+|�<@�֑�dL��&^^��)��tY<H�7�{{���3��\�9�!!!���8 HI7�)g�J����U�����`����V������:3�6�(�xqF�K��3�TUQ1FQ��6Q��迻��??���	}����VN67C,��r��A^��/|^�S�+ ����6<;3cz�Lk��5���B�"Ґ{HG���a���������ZV��×dz���rf԰����X���a�'�k�KKK��~6�{�"�����Pt��p{��X��㸊w��a;�b���4��XT� ��ZΠ�����V0�����xƢ���}CR�����`�x�U�5{�T�����n�6�I�ݢT��Zfvv5�������S-�1N�z<����0�������Y5�k��S����
�����w<;1{�w�o0�---7o<.L%iM ��2t.���ބ���x��� ��d�MTTUɣC���Cj����YY���S���XR9ق�Kj�lG��Y�M�kfE
_�R�q�QЪ<`m;����a�eͲ�ﳷ��LL�Fl}PPPM_t���}�`@W��*�����"�	��ַ�>P��/ U��B�aԀ�M��䤉���1���8���	6��a�,u�����aO��J+N6����D�<J�ڿ.[����ԁ/>�V�עƾ��?�8�� ֕X �"����y�����i ��x���l�RU- ����%�;95OV��J�?��>\�h�gVVT��Pw�m���|�̠~+GϥX���ߟ��=�ǁ��j�yr�@d�6�z�F��ّaRu^�,,R0�Mώ���t����zG��������H�+cy%��?�����P\V�lE�N���X�vEEMflYzR �E�O�tX��"i�����12r�W�`�<����V�O��]Jq�p?VW3ihi1,�=�l�R�|ka0�����f.nQy�Hp�����\��/����GB�麱�<�����@@Iep�glY�{ ���xs��mڸ��L؟(����S��Kv#e�D+���+q��wy������[�,@�,���b+���<x �ZKFN����f~�)~��R���J���ү�H+Ů��W�e�v�xui����1��.Խ��w�׷C�*��K�6�4���`����C�/� �&ef,d���,K��_���LN���;J߽Xx/�d���'�¸��s4�B�)ρI�g���J��g��(>RH�o�./�u.0Ov\�~pA�ζ������HC��/� �޼C+���q���ݥ&&&V�R�}dv�e����Fމ3�ы|�Ʉ�����-C�
�A�$�_D�[��Ha�>���,����IK��K��ɗ> ���8��xK�+���W�Z��p�		ś%��"�Me-��L燤���h��p�|��LA�8nN�ț���}����+���6&]|�8q}@�᱄� �H�~�Z���3 �_?l�G��'���q�VF�r#���fO`�F9+9�
�z��-�Ŭ����S��1J:�jcVvvv��;	���8�N��o�����Z�R�)��Sۛ(ǹ����apЎ-<*j�Y�]�o���Ʌ�+'JM���Ͼ�<g=E0�SQ��cł� �A����众<�k��R+���	����6�o��x���#	d�����s`�S=�Z��&&�{������X��a��	��׿�g����V1 ����O�z��[�����F�و�5섺�Ȃ��"X��m�b�bq�ƹ�P���������13��%Ď�L�-Y�.>Ś���6)��C��9GDD,5�i'D,����s�gga��NE�Z7J>��"����=W��t8�I��U�2���C�[)�Y�j���̆cev�`'Oâ:~�6��j`��MMHK���RPv6�Y��%�J���2j�^\�TN�˗�����o\������ �e�ms�䝕��	a��ƅ��1ܹ���w�ܜ��J3�e�xpԜl�����>�B�X��J��M�MH�37߭ �/������,�Z�%��<��lB7��K%%�Ž}k}�?)�f��FD�8y�O��77��8$�Z��({IC��^�D�H��^��>����˗/%,o��j����4��@ꤚbX�ٕ�ݜ^�Ե��F�O�.r%7�|�9��x��ͪx����ذ0��b�#�w��eHH�84�����~�BCff��/��9E��0%G��6�aa�#CDv�b�P�{Do���p�ss�Yoyv�A	!��\]/��:ҋ�G��ⱥ{HA�̩t�EC|gn>l?Q��� �XFN�^���0��&CI�TNT���E�N�xH������Z[5# 4j��V���w��Fp������q�V$��b�FF�W�pQ�������Re��˺׻���ߑL?� ��0����Ob�R �6;�T��Q���������(:R����Ng����.:Zd%wW �PMOeƣ��3G�_T��"ԸdX#lzt�q_��57{f%_��kÞ��(u�Z������t�P��˥�_wITտ��B^
QQљKǰ���~T��,+�4�H���Z=e�ީ���dsw[FKOO33��VۏT�Th�v(��Z5_��yk�[YIߏg�vjkk[�YV��*��v����+�}_�B?~����Y���[q�=%�0�C�п���IL,4HS�?��WV��v�ڶ9�����,-�٭��=�g��o��}��XL��� �������b��w/ O�$�u�4����6�����G(�I�RQ9{�fg'�8dϭ�/&�\W���>�N��#��5;���8B#`nn������L��Q�m��0ݗe�|@�������|�
���&̞���"�z�m&DA���^u�0О���cF>���V�goP��}����a������҂�@�Z��������F]r����%�;JM��=h5���`���in.a? φ'��M����	F�5o����|��*Z��К�2i\LX���NRh���|��o1))IԽc�>��0K��2�ּ����%�
z�-hA|C�T�1�&&������u qJi/t���_\�\��>�O�:�3�����
�m��[ ��*�?8\��#�q�1��k%=�3�D�"Ki�`�e.;��AXX0LݖTRz�y��E�,�!eOs]�s5 xm����g���h�����Դ��w�XS��2�2i���v�)�ZD��W�ejY�v;P�aȚ��D�������S'����
P	;īr!)1����a*�Y�3�|}���� m}I��vg��0X}m8��bv{�62:�Z���s۳㩾�{=[`�)^���R����l�{_�p}�������ӧv���F��J��#ww�W}�?�(j��'�F�m����k��N�q�왷��nὂ��ͯ��9�j�7oLML�pkEJ71�i�3��񮳜��1߿��i��l5���q}�~��+��0���1��ه���㨜���6��?�5]7�|�p����((A����1!���~��x.�
���\����Lq�����Bzp9a����D�w=�n�L̡��LpSp��o���C�Y����3�966F�7����laa����	�z�j;Hx�a�\]ծ��zZgz�<<<"ݔ
����׍�[�n����\t2�`�T���:�+ڸ��歞C>��W��Yf-�G�e�����&).�{@�ru0�x{HG����zwS����!=�d!P�O��k����ߪ��K�g�7�V �� �G4f!�*,���#)���jYE���!�ñ�5|#a��{ߔwx�IA��&���<Ѐ`I{FGVSW@<���Z�V^�YC_�3��]ǌL�-�9�dL�w�dw��mP����*nn�5OB��8>8��/; s$;��O�o|���6�!ǚy��w����9�������������
{�§7��/�ol8Ay�1�� =�-��u�|s�]|PF��n F�	X��S׶��'\��c&�/�
�9�
�E�M�8�ӷ�����EL����~�aO%�t�������ҧ?��q��'��� �]㦼sԙL�%�g�"��J�(�ư���CX duu�D�fx-0�):��:��y��T��l��#Q<�������j� A~���C!������(("_�rr�99~e�嵂J�����w����!A�V�� �a�	�����Y���B�O���J���2ܜ��P���C<I�b1�{OQ�Sx���F� '&D^N�C�Z��g{+M��%�N0�:::2=�^)aO�o\�̇d�U���į�.Bj�1�v�k����_���U���l�HS��KU������"`�$I߳���2��h����X����v ����b�˯�b�"..�q���&��r-��WWW�ޝ\"j�=��z��lP�[�l���]x�8�;���8~��QD�p���/����@���
pp<�٨�r��F�<�x�l��~��XSSS^�f�Ź "�W��N�>#%!!/y<�$S������ü�H�?�T�cb����@��q��~;�:�=�ӁW��2U\�ķ^��El�ۛ��� #z�-��ls����l����U�K���]1��v{�oE�������E!������0;���j�3sL֧j�7 ����������� ��t�T���q���I����CIq6 �w�:|#��Ͽ��Q��4lie��vŐ�/�i��f,��;�����muuu<||1�fe32YYQ�nOG�hS�JY�S�D�}	���g�WQQ�c�:n������SԁlC)�ǡ}�r ��������by�����t�U��ƃ�?KKx4��	���j��LL��J��������}����!����t(�   � �?iiA:�����n8��y���k���s�>�]{���u��Yw��c�y3'O�K�]+)���&��M�uS-�g�xE�{��n����a<b���2g˗�c07?O�U^Qa�fxǣ�Y�8����F_�A'�}��ְ(e�W�s8�b���׺�4qW'�S����8g�p���h|A	#�폾��CLN���}dt:&�!5�?���E�6'��?H^N���I�(����o�Ů��O��������q	��M������MC0I5��Yd�yb�
���r�vJ-9e�>F�	����pvO|E�!? H����eAr\��[mں,�X���������M���V �1iE(��*ɥgmU� �}��K�W0z������@)��p��B8�����n�Re��[/A9��g(n�);�;��'g��p���Ri�����ڎ���G�Z$��(51Y����^#����&4�H:�"�t&uȨE�����׽5w�Va' ����i�C��F�9��3P.��tt<���RQQ5����hڭZ'����;�wV��a�$M��|�:0���=`�ye���	����%D�oC���1c?5CZ����F����S�X�:�����1iI?~0Y��������;L�Aߩ<=�i��,��	�)V`L"��gn��vw��U44�9�o�Ian� �p�,���/,L�:W�	oUUU�r')5�H�/=c��j�f9�g��Bp0!a��O�*0��*�d0A �-/C{��!�?l澴�8A$"@��ɭ�'##�u�E�����ôؿ��M$-����W��swq���jw'�y���2qnjK33��R4"�T���W�^5��h���S������kq��ݢ�d�+v=T��_X��e��q��G*�+nd��(f5���3���~(77N����obB�D��oo�Ű3�ǌ��(r��a�E�����z�&���r�.�O@�+�48Y�9�S�>�S/.�`�5����������w���h�a��{��P�&:Pmq:�]�PS�Tد�����=���,�=�O�.#u���k麪v�4C�mݯ?�g������),,9+�N�Q�6:6V�2��&��GW�V2���)F�t���l~�"��-P��GFj�H)�牗5)����Bӄ�����^��plx8���c�H����rM��~�s`2�,j�l�w�9���g�@�i���~蛝͢!`lO8��.%F����P�u�^vc�Y�T�ggg�,��*c*�ٌ��"��X.B�
TD���
(SZ�X
m�"I=����%{�:,a���11o�÷�Z���o�4DDP�h�$''�z�(�H<��QqY���8o&��K<@S�N$�����n5j^�TRB������^�U@�F�%c?n�<c��e``���Nܑ�2��]ݔ+B���je;=}����l�����]I��(�bb��hvW7j��A�������`�����D|���)8s^ ��AY�Ԃ�#t��g�>&.F'����ØrC�ߋ��x�����`s���LJ��|����� �ה�ǃ>�;1\]]�JʍZ������P2�����G	er���|�QC*��I��L�F������ٷ�\�طo߆��`-�����v�ٸ����u���e�|[��kc��3�e#��vu0����F��@ws�ji}]tqa!��'e�I�-�
*��@�}��uj!�B�@���S�����@��uv���zt'Vy�Q�o�� ���s4����K�hWW�6�5�CDW�7��Z�]�P��_W�_�gd���C1H{��U~�����;|||]��>aN�����ۃX��DL��eq�f�H{2�i`������z%�X���ۄ�c�c������,��� �׿׵z��f��XH���62*���뛭ܪm���l�V��Ņ\(�z��3L��|���E�%����=�o�y��9͚�< ��H+��R�q�����NU��<��V�i����������Vg6P��1z�oV�Y�ە��;H�]S��p�WOW����>���M�::�#��l<<��U��j^7Ťu�p�	b��I��}n�Ui��>h"�
s���!��Va��IH���R����$;�n.|:>�@�c��.&f��(�ud#@f���dea�����R7Kv�F��RssT�-��7UL�B���v�z�]���9�<���	�B�׽���*�h@_5�����`�y�=*1QT,ՎO�@��/U�c��I'���8����/��sǓ�|�YE����w��5Z�׈�M�դ��ԣ�4s �nxP3�xS7pz<C|W>C�CVK*�/�(�F+��)�9;P�j��Z.h�Ĥ1T��uwY{q���x�]ה"�������������j����!�Ӹ�z��S���=�ؔ!�bRNM�)�{�!��8w�^T��^��]K�ح��e���R��׊���$��Q\�7�8 'Ν�zbk���i�yR#��y�Bg�����Ɔ�.����J3l����r>��r�C���[���M��Re�L�����"���կ��ܱJ?^���D^�����=%b�ؐ���(��k����Y�>�����Q�VJV�	��R[{{�A�*iu�C����["��.�W��>nN=k��j�٘!�C�I�u>�P�L�߳3��{�9�>����(e2�������r2%�'�7��ۭ`�|�oA�������Zß=9��P�st�I�O I0�i��F�.`X���p��Zl$�&a��pOF���>�!Ad���	��~�j,����X��=1;Қo�
FJPY�a�qE�����A����5tt���� �m�)��<6�£��K��$��5T�����u!�\]E?_#s�]���;�Ce��F
��a����/�V��,mlT'�R2��VD~g*�|�����1�;�ɼ3)bb�F���x_�Wo�d|'1,1�fbc�cٸ����-;[�RW<�Ou���ӓ2|��\�Gn/�N���YD0�B�b	�'�������Նģ����r?S�YilqGhVt4�e�'�s 77�T-@�����C��^wT� ˆr��᳀��eee@cW-N36�E��xj����g(z��98���q���$���4ip�Ŕ�<��'Q�X�z���}H����e��3�6�*JrH���ˆ��.��&�Ť�'���y��jcy�	��������-&5��4�; �)}�h7�#r�>I߾�o4�i���V�;;��1g��>��B�/�;�F�Y���3(��UU��h���@Ǣbc�kk ���&)��i ��Iy+46�,rVLMM���ҽ��F��:�">������H_�;��R�V5�[��y�|����C���^�����f���)=K�	�`h(���~�,�n�3?�|��V�n�*��+���q�y�8a�dw�=�k*5n�.BT�2��zǲ�y-���?]����(+����G'S��욂 Vぺ0����l����nnBUǰ�L����s��܏A���EE�+J�xxWO���B�����6s?Ш<�fU����d��K��ǎP�߼�BĢ^��D�m�vj�ZUUՖ�v�m�m�F����
����<���R�o͏��87G��� ����߀Y�z
�߾�64\A��`cg��l\���֭�@?��ȁ35��,���tJdI��+X���:������/��j���]]3�E������y=󸽽��S�~�'�}3�5��I[���單.�'OPb�iRŤ��͛=ߣ�̱����>���K�deg@��g``�,9Tfe����5sß?���n8s���>���éCJ|�1��w��3M�J�*��ܖq��U.]�BBC��,���o��X��:�geA��/5�(#&��[�Mᅕ������c�7�5��ŵ�4-.,<��^�������j�L�qq.G��LLX ��:�4���Ra���@��2y��;�[=���Tn|_w�:�G�ln��"�Y	%00P�֖ ?*:Z5BZ��ʧO�>FD@�g@r�����id��[Κ���^�AhG��Pl��i�J�������	�_��NJZ�:�an�.t�4�rGg�v��i�; ���*��R��荟]Q�ƻ�^Y�}�5�B;���qF�-�QW���SP���P\�v���IĶ��QQQ�--�`R@"Xe��A����2���hA|󙤤�uM�~õLR����%6�ӧwmmR/_���
���u��	����LU�\kGǜ�ӏ
ɏD�N6�'��ٯ�I�6�{�YRsz=��=몄BqQ57w��� �pۣ{�VHѕ�6~� ���37�t����Wn�@�N�����&���}��U�:���ٳ��{�SŃ��E{ y���+������2����{A�����C7�1H�BH!���x�~�(�1�`�5�a �C��w��לh.Ug�����2ʷ[��o�^��PƯ-���+�t�, $��b���1��NB�i�0&M�� Z�]wz*�)SQ)�Z�!���!��VQ�墾Kg�KX8$�L�D�Ǩ�s�W���QY��lh
��j�N��	���x��
�&���N��7�Y7ղ�*ԝ���3k�D���}��JJstf�������&:1��bTA�5��fffu;���\��@����JIU�gO��f$x��Z}X|�q����������EL��˭6wwvB�̴^B�d����9��3倂QQQ��iH�*����b!�ŻQ-7֋}���1���f
�?�C�RRR"

��
:e�z@�����\����aq��fMH�������6z6|���4w�E	�� P(�t]'ss�6?!�Ia�_~�.�}Ν�E�������LUU-�eT���S�w<x��-R~�0�$_���r�A��ו�w���l��Ֆ����Q�j�K3U�y�2�;O������&qps�@�(f�d��Ykt/�'��'�{";������O<%"�P�nh�aR�&�\�"m�xp�E�#nnQ�ʇ�@�nܸ�4c�7;d���Rx��E%6opO�5���U�耂奬?\I��'&��� ��*����Ţ>��,@3��J4�voS�|���p��M���W�\D�i�/��=Y1�e�q��g|��gZZT>|����7�s��$?��Wh�_�Y�Ģ���!���b�����+�YqQ�lҗtI�Ĩ��%[���=���rrs3�W�^7�φ{�QR,o�7��=U|��m����.W����Ҷ�R�ni%HA�A����%�S�=�6߬2��[}MM�{��v[/����v�P�g��X� .�}}�ł�3���@i���H<L��ʯ���]Q��e�0��!�e&H1���4[�����HߖOP�M@��U��rƖ�����f�w~NDj}xav��k^^c�Wbұ��AC�,7�rj��LݥI*Z? � �erJJ=Ո�������bc�G�|�����$��!k�&'@)�x�kX�]�l��'a�|���"r@G-=K����?	���|@�P��SL��n`"�i�����ʩ�LB���EMLLD�7h��3�*Ɉ��#񻌡׻��wBi�K�o��%̉3�n�W�QL�Ŋ&&1�yŪ����"���^�92�ٛ40����m��XM���&'u���_N��}�};�ss=�G@2��`��d���#{r������p0d�a�q�VS�lZR�ˮ����uj\�uӗ����n����̳���o"��!��V��ں����nȸo|�_G(Y�Ggc�RF5� �m�<ruz����5�O5'_�����_��#�3���g�	��EJO��^4m��7��tx�0��%6��=� r�AF��`/�vmrt�L�'X��hZ^�������ׯ�'L��J�a��B{��ٰ��<���h+�?|���5�a��#l*�}�y����bddd��$�
3���3cq����S�xdb�"k&C��]+�I3�A�xY�9���J_�m�cwZs�y0?L��y3��*(�]�@�2����񕓚���]��Q\u���ritx�W���/�PPP�a1(*����?�G�OǏK��ދ?��b�o �uo��C����GtrI��	��rS:������'Т+iG�>>��,�NN���57�P`��l��0'����׷��DI9����
�L�zzC;M���&1�2�}���'*)ٰ|��GBB���\�#�k4b��T.Degg奓��[�͟��$HHIE�ݞH���<��I.���#��VS�T��!��Vf��3���)����\�CV\u!�ݕ8ew�T��_f�Q{��\�$��G.��,�Y�%��E��8�O�~Q757��4g�14���#�轜ݏn�aa�#:�f�s��/~�PcԬֆ���fb��[e@��`y[u�t�'���PP�;;W��@�-��J��f���T�J��-��=}\���M�A`I+��uN�Y�?�r��������2.G]�����Y���4hYJ����X`^��ލ�	-�:�Ց�:�W��f�Z��0�ŘZw _l+Z���������l�\H�j���ɐ�	��Ɏ%<4�O��X��n8k�����'����(w�h�)�eCb�<��1i�f�A�����ēݞ���X�k�4��,�rϞ���Q�����V@�.o��.�镞DRh����M=�\���ٹwp0]�b��(�u�][��^��Z4v�"% ���yC���«�"���菷��ee|���C�*���P��el
T� ���9أ�:��IS�����cR��$qx��|�o߾&��=��:���t]�?�:8�&��������j�ᚗ5>{�#��t����R|�y��%Ar�K|��9u_�:�C!Y���ҧ{�����,�V���R�,YG�_�U�4��1P������ɟ;&mz(O����������J�&^c�xNM�Z�����en��q}mhNpGQ��o�)��U���Z�߸Y���X{VJ
�ĳ�R�;2l둾�3r}k�B�s�m��@G'�B�	ӻ:�H1��B�k&$H�K,�+6�+ŵ�+��-�
?����}s��� ���P�@�9��8x||}x
���R�Wvy6]ݳ��	�I��?:Ip�n�vt�D�k��[�2.�!P&���3��7[}k�.Ql�#Тs� %)	Z�C�p~~��T1�Fv�"�J/���M��?��A�jdi���NA
�C
���7��٢Kx�<i)b 6x��'_�Y+=�����������=ݕ�	oRғa�Gv���[w�\������M���@Gyҗb�v�P�3��>�Ht�,�O�|6w�Ǘr��ꛦ&	B�^b
� �����	�f�L__����t[�aruiC�@�$̤Dw山��w��~Ml��2����l_��߸�\�A>~���qs3n�ۅ+"���\gb�������Z�8]��F�"��ȿ˴���H�P*���{����r �{*T
�ŷ�@��Av��C��s�WX��\��4�����V(�+��G� ��f�_�
l�&(��T�o��zom;;�-b�]�핏��w&z�
��xTY��M��BX�}}i�Ύ���{֖@��KC�ˁ��	�,����k�
�� ��g;x�ڂ)lllx��~�������Î�||;���>�\��P_ߟC"�c�[^��k�
����____Z]U�Vz�H�b���w �?������"0����yC+��MXH�+�̤��!&�`�:99t;��$TIFFF�%*�]0H��`}+�S��PR�*'������]1�W�������28���	.N���FH���?�B}ӿ�w*K�ov$��k�ϫP���h<�ng���	�:(�1܃>�������a���k*�����AC[T4��MYYY�^Aˇ��[�M�:
x�I��*����X�S��2�ז��� X�(`���?$��u8�b��c�nZ��Տ ����wm<d��qSx�o\]]yl��rӉ�Τe;R��.;��v�������!�P�솭�;o)�	�*6�p���k\y���Gl��B���n�=攩�M��)�
���	�BQ���Rx���Z�����`��d�A��g��Sy�V��.�6��$j<���qc��$CC�T�d�脄&p�ܝwO\N��ZHI�/�@	�	.����԰��Mj���9�0u$�s��X(I�u���yI(���/�e��
��ϽֺyMKCs=R��_�4�R��M�����˚��xnvv�o��Y�7��&@�y��UWA�"�a+
怆�DTj��g ����� ÐEυ���y��������踸��z6n�t5|�N$��Q��6��汹$WSv9��e���C�PGm}o��L��%���3E;�hC������E���t K��ɴ���d5tn�`��N[8�u����kѠ���Qۈ��iH������Vl��yz�DW���+0��*I_ڠe��rr�-��x�3�gؙ�N}S@[� �<x�F�gt4 $�-���� �K�|po�x@��ҜC��V��9�˩�g�����x%��,�bQMQ�rgk�O�c���M ���A��__���M	z����@���~����z�b�"�#=��
2�r3������x��=!^����]����x����B^s(��(�]��S��-���fFF�`e�*B�_����n�|?r!tC�_����<:;;�����c��Y/��8D��jgX�h�q1h�O����%�絹���d
.Ǡl|&V����_J�1�O�n!��/�yCԂ���3빧�!�����2h*�'��$�����22�rœ0St	S���]q��!?�y�'�r�xI��Xڃ��R9�ե;���������A�(��v]� �R���N.��5,���Ə��\y��=G��CNN/��m���m�,�?����,,��K����.�M�h�f��;0��.��.zE5��c��V�;��6k���rwT)��+t� i��D���9���C�J�V�^����r�ة�	vO���d]�m^ ߳'NiG�D �??w�;r�#t��򔊌�HB~24�@&G�SQPhl�s6��������v�� E�k���c~.�o+����ZA	��u9��X�2Q��H��QnR^�W0����ѭ�g䲍s�^�~r}�^N��`
QK����+B��4��w�o_&��V�}�
��2��6��e%c���ۛ���������f�����9d�w� =����|������?��l�:_�|��龘KǓ��0�u��r���TZ�X&2\�ӛ���РJHA������:� *�NC�<�q� ����[iiiVK=ԁ[:�cX�"<�ǜPu�L��:��ώN.�#0�ƀ�6���)Eu�0���}�D @
/ꃣ�&4�K(�[𘾏v�����sn�a�����4k�����~�#�tBw�g�[K�cG��7OI�i�o����-pL���\��E�^2�F(���Dϵ�'.�!w�Mڦ�$�S򠢸���NSǽ�
	��O��f�kxק��k<��C�� 9Mi�F(�Y�|z3�TF�vUm�&�V,9Aj�*�;bbe &�{Q��>�aX�#w�J�G����?�QX������>�.�RM��,�#�6:&����=�4ş��I�Y5���ZS�8{X������ܦP�����b��3ܙc�Ȧ��?�9��������Afᕢ=\�P �u��h�s�HM����^u���"���V��l��V3��	��N���¬��n]����_�5�%�R�Z�a���?�f5ю��6���=�q%EXr�o���t{`XII��9G$�F������iǅ�q:�9'vDZ/-�V�9�բ�Y7!..B�2����H�nW;����`�0�l�>����sna����fU��Oo�����]���ezV֐��i����>]�[�����>�y��a�S��'999���������֨�D,�@���'$$g[��gff��km�JSh5]ςJy���BCC�����@i�^s�8�&�j6�$��v�\�vN N������D�ܢw>��x�����\i�Sig�/���Jb��M�_��Q�|�5�U�6�s�<��o��, �ӤLMM�y��,:�
n��Y6�����!�jx�Y4O�W�vK��=��3|'����.9?�}q� �M
�c��kc(Q��N��N�?lͱY���H��d��H��W�#�]z'�X�wd	ܔC[Q{��5��tC�oA۠���y�
j%y�[ Iӥg�\�6A�>r��#Z@���a�s�q�=p�څhy}=�ӧOF���;o���edd��U�K� ����GN��?B�Q� �9�w6[Ӱ�ۋ�up�s$��\�.}�W��s�L#_eMwZ��+X�g��[c'���W�vJ���{��!�*��E����L��U&ݛ����Kc�q�Mh���f���\�=��aee%��!��e��#������;S����]Яx~`4DD�7������������a&��\8Q��2b��[NѤ��~���Ғ��� �lV=E�I����������g�����GKSFF�f�����j�0%ep������&�`Tk�����݄�?l��������G�A�j��Qe�Z�6S��u\H	���:�a^�#�g��=���f���Lak��艉	�nkЂB �����n�:/-�F���:�H����ٍO}C�!z��YQ@֑kCy�22����p[�ͭ��P
�L8b9����=�����:��dk�`k;ֲ)_}�+MrQ�#)i��w�9ׂ����/Η6���C;�"��n��y���<��D�(��;ÙZO4ދ�ٕ�N�Y�^��E�r������o�F<��h�]���M���d��ZeZ���Q�Ҳ���(R�N&!��i�� ��u���l��̢{mng����Z]�8�|||����6���/ZZ�����m�]@������GO,�P?�()!������x�w:g�-,�A�>Th�ȬY�Ӎ���fP���w������,� ^��`����s]�]}7-��?]y���.��8Nۣ���陘���J���t�ct���321�TT�/F;������F��o� N��u5I[VQ�v�9�?ڈn/���Zp�U�&Gӑ���f%��۷{cg��|7���.�9"��[S�6`l*��$@Oj���}��x�������T��<K��[�!��-/����돊�+�W�������B4ߙ�w`�#1�=���]]]*����J�UU���uy�����N��n��<�5S`8[48�6Z"و��$�?9I5??��r�=T��Sw�sJ��8�ܠDY�}c	��N���^ǹ ֔/�B�է�꯭�k��*�de=�2!��d����rS3�����k�7^���w��sr��C�8���3�%'w��'���ޅ���V1PB�����������f�l|[��̉ʟ-�
]�`�e?iŭ*O&��5i��d+��C1�hOO�o߾�È34�gGnrO6h����K�]�蔕�ޮ�ݲ��O�y�,�0�0ҍ
*@���̓��0�^s^�ֻq㆘�>��沎�[�[K������
l�������*ÿ��\�?,t��;;;���5B#�,Zw�OU����+���t%�!a��X٥go��8�� �b�d���*�N����V������3=I����W߾}���Ls|rb����Ǐ�u���¢�n{��j�~#��5�s��ۆruD;H�k����S|����!D�5D��Rb�/)�ޤ4k���n��XX,��h���.�m5�|�_�����Z������r�f*����)�[�Ԋ���mf�2��ϟQ�L_%�݋�Ͳb��8�='��)m���lh�}3Pda5�Seg���U��/_��"����2�|\d�~
J��JJ��~١���}f<s��USR��p�;��3�5���s�<��j��q�eT��%&�������߁۳O��U�ϴ�\ܒ�ŨU2{bi��xP�sz8�\�l�p#����,���X%OW<!���������\�T�z�F�ϥ�8[u�"����r��h����0� z,��A��!g�TJ�t�S/�V��B�H��I��7���X^���2S4y�U�#�It;���e�-,,r�f&e�l�ك� �����Ykkjr<ͩЭ;�q�f��4�w�Tn<�Bŏ��/�j�>III�d(�ٯ�D�;X$���t%
S������N���+�N�R�%�R�m*�EV��⧄�w�H�b8���TASQQ�����|��maP䒂��;4�3���b�W߫�55yA	w��B����i�<�&X	;oӛ��5���T��lsJ^�
��֝��=`�A&fc��5�a�2B���L��L��L���9�c�e6��(�� ���B�W�*x���AN���aTD���###Kqs�Ngg[-DZM+mm2�� ���%K9��X�g�����}���oo��`O ߾� bN�p?9/��"ۚ��id�*j�$���D��3IԹb�@Qť��E����3���;��j����ʟ1��8�T8n������� ��Ī��M��0nְ�n����I���Z�3�3�"��2�n�y���'�U��5N�&|"���k��ђr[Ff��mg�g��2cڰ��	,"����Ї��,��U�g��%@fr^�5��ϸbX6�|��]	�K���-!$@���3�g�ZL�7�j��4HyW�44�K�26�[�o��}�Du�JW�B����ӫvvy�yl�B�*��Ku-������$�5]�;ڞwJ�=^^^��YZ^��][��p�۩i��:ԏ�D�fc��@E�{�Q֞�,))��Y�w��u�W�E���s�aa}�4���Dj�� ]i�E|���m�f�.p��B~\pӒ����(`������oYYA��4�cA۾�\5�_pd�\$�2�ݯ��r)ss�* � ��5i{$+��Q��n���Xj������'���:X%�N�22L�QɟS֨Z��8r�?��pC�/��O���&���o«W��t�D���k�Q� �1H�ٸZB�c)�[��7�M<T�aI	�߃
�f󁁭u,��Ț��V�lgg� E�b`�����u�0��)�<��'W��aB�Hg,��=;;����A��S��z��y�?�&|Hw�:�Z�8j�gc���P�'L���x\�N0���2�J��ap(a�o�l��MfFX�
9+(w@��/X����r|Oulh<ާq;��b��@�7Fk���2$�i�:��+`vTʬ�3�j�:�Ú�����[ff�.4�Dʂ�%��@�)�yp�r�����&�r�����0y�/{�sHV�WJ<y�$�.�D�����Ø�E}nmo��t@�y��A���ZDQq(w���$K,:˨͜`x/v��j�

�5��HM�+3s� ����xX�ME��,|���B�#���+[=zgmjJ;N�����7�쾵�)ȸ��偸�i��A 
9��_��)!�Am'�!σ�����ք������9�Vw�b�3;�W/%�[�a#�À������8�L��G^r�9��������jjtA��k+��k~��ۜ�_�7z^����8�:�;7J�:�_�A=`JIJ��u�����z�<	(:���F\�r����F#+p�8�q)�8�3	���.�;3G��/��AC(�:��T�.����i�o��h��n�1���z�W����A�]8<po�ꄩ���.~�XZBڋ�[7%u�XJ��b����!��jf�w���ɸ*yCNcA-|�1N�Li�O�kȏ�p�ZwH.�Fߖ���6b\ �t�\b���`�^�����P�L��I L�KL�F�r��^V�^ D�u������)����M��N�����C���L߻����ť)��CU��j7ɐD�;�3J6*tĹ���M��������u,��X\r��{���h�ZU��˝�.��9DF�H��x�<)iH]�ԁ�禍�D�[r�S�'c����b����C$/��e�����,v5�9W��Ny�Sz5�Gbk��9�y�OQ����3T�8���hs8d5g4&�)4����|�	ɏ�%2�nTt?6�h������չ���ʈ����x�����9_�Y6X���b�@���qL��=C2zXdP)��]���yv��o�x�o�7���Fx#��o�7���ƿ7�^�_�~B?R�ӓD^a�����a�	&�`�	&�`�	&����>j���WjL0�L��t���a��[R~����~b����0�L0�L0�L0�L0��oK>CEz(�G�'�����Q�ފ��נ�L0���hes�c-��R�`�	&�`�	&�`�	�?�3mF��}�������rs�n��L0�L0�L0�L0�ӿ1�j�B@<g)Dш�����p���ݻ']��� �o�&�`�	&�`�	&�`�	&�`�	&������R2�+�
L0�L0�L0��I
���X��.�`�	&��W��~AY��^&L0�L0�L0�L0�L0�{���R�wW�(���L0�L���xw����WjL0�L0�L0���1��/(c���{W�`�	&�`�	&�`�	&�`�	&�`����k#yЏ�w�W����ި��
��8��L��Z��v�L0�L0�L0�L0��/O��Kɰ����+L0�L0�L0�L�=��$D�?���&�`��ߙ�)� ��]��<����*7�P��&�`�	&�`�	&�`�	&�`�	&���z)Y�)��w�	&�`�	&������A��\�/�.�`�	&�`�	&�`�����e�W��&�`�	&�`�	&�`�	&�`�	&��=�|)YޝR������_P�>��\�/�.�`�	&�`�	&�`�	&�`�	&���z)���:��w�	&�`�	&�`�	&�`��ߔLʮ.��Z��v�L0��ѝ�{Z���Ç�x��^�e�^�Heܪ`d#&���0p�����i!�NCxO�^H�����>	&�?�Z���痡����ol�yW��W�������������������:�p�R�r��m�C�Csss���`L1��Cs�92p�G�F��g�·C�����\�"z��;76G��I��:8<���o�DGU�^�5T��L#U�	d�L;�!SLc�Q�[��#z��^�<���W���泅���c�Jt�!i�UiW�Mu�T�װ�(Ssu����n:��G�=�"�K�bˡ�ܷ��0{voc�m�k[cpe�zk�N]�ET����躹��iZ�F���VtE���՛���H}�����	Q�ȕ!u}���wln�.L�T�����:�Y&��f�\�A�mw�@����v���)��S26����'{���DI6������$��.$g�ܓk"d!ȉM�(=��⒱��pر�����+R�4��/_����7	�|��c��p���J�w?G��� �C�x�k�V��,e�K���`�����F�cZ���[�o�<L<f³���]�ŗhB�;fQA;˅���%9V�@N�eR�#Q�n��y��;S�r���{�u?t�u���H[\�I�׋T�eRH]�����}D�%��*���g`W�H�xe��\S�[��T��\��֌��l��6�=�Y�7��J5z�bi��a��{d�'<(���>σ��e������ǻ���J�E����3Ol��^[��(E,Y���ʙ��؈�L��
~�(�Ր�d�#
"O�J�T�p�YXZXq����9;��ɸ��F�u-�� �2��=�����D��3QQR�1?�B*)�D[�n6�mQ�^�s�����dC�x����jܾb�~�0�T�ˢCè{8��3������:������l@�����I���~?�j�7�p�{Jt��@gg�JX�Mi^۾���p����?�����9�芔�B��8/�Kx0\'�ݏ�mƨV��w�lV��aw,���w�UT�#��dŕ4����0ܱ�>�2?.�z�t�2;��^WSW���:{�h���J�^qT��0�Gٕ��ObZ����p���!��H:�m;�0=.(��eu�t�`H2��n~��}RV�-��X����]�Z������y?%�M����#���5�B�?%��x:��M��r�����5Q�� S�k7-؁����H���w#ׯ�&e	].�i��*��GM�r�m
qZ���o��I��>�D�߯��ש�S}���}%�._�k��\�Bف@8��q2���/&Y�⨳����M{����
s*%m�]<�E��h�z�z>��x����8�T����h����(.�ѭ+�/κ������fpHm+�msj��y-�I
�_��B�K%�d���a�;��d[���?������^��8��(��H��u֫�5�|��텕~��h�v56FZ�?X�V��ȃ~P&�	�&���|5�X��/>ݽ)�`gWd�yl�[h@���\������Yyb��h�p�aƑ?h377��r�>H9�K��@�A�"F������J��E*D[����6D�9w+��H#g~m�8�<��@6��;88����u!�bu�e��m:�D�*��R�֗�1:ܟ�_��~"�aC���$��ё�����N���0T�t��2y0����38f�)���l��#|>�ko�̗���|{Y�a*��s�l�b�e`@���'Q�Bg��A����S�F�҇wf	F�G�*!"XB.���-��_��徶[�/0��9P�#R#Q��$��-��ow:�۳��9 ��dҡ��Ч�ө�̥7�@�1p�S-!R=�������n�����L?�����zQW�*���HV�����hBv��7�$�u�D��kιv�k�NJ�'����X����ל�]�֊e �ܛ�:��Nϝ*�צ������O���hbwQh>�G}N1�m�����F�;�����5���d�z�]�[�QiQCmL�����V���q~��W�{v�2�e����-"�C��2���k~8���_���a4�(���ф��ؑ;/����st->z���<���k�fW�2������kpegg�w�4�HQ
��n�&���8�ܽ�A辬��N����&/ϴ��N=_c!��m�՟���/���x�&���<���i%Y�nn�s<��w�拇mGG�`�bC������X�޻���Y���G�ÑH�v���L�jv�d�f_�y�b�����'❶���Ú�x��Pݰ{�XR��B^���Z���č.���z����M/8=���tp�D��w�V��	�I�A:X����a�'�`��G~���"m��|?	�0˧�mf�^{�k�Η��$�L�xS��,0����^'Am���o]�M\��������g�C큛O?Tq�QJߺVD̥S��/`.�LU>SUSk�i�2��6�{=a��!�=�%����V�����{OP��y�_�����f��37��(�ڎ^>}���K�V���=�,���篤�������j*�@�RT@�4��;( @:!t���{U��K'�I��"��N@z�.��|�}���p���F`@r���k�5ל;gĕ�6�}៯�)�FA=M�|AM�9����(�77��rL��k?�������BB��t�����)���3NJ��^�7��&n}������\ɽS����d_45G�E�I�pss�]�ٹ��i�'����G�x�G�<�W��_�j]�|)�-fzx�K�8�
�{3�}hP��fl����!�/�sI����O5ǌ��=caA��?W����n�^%���f�"�����*��Bic�$����m�1��w��J���J���h�QǦ�y���w/@\�]/�Ŕ+{�v���D������=��X�s�S{����/	~��m����HJ�0���O�)G�·'S��'ml�'���!�g??�p�p�s��h��0�E@��&ja�m^��J*%����k|�� G5A
�����׹���mm{iISa}��{뒜�܅ВZ����W�e�2�Nl���$b�����;�D���J�6m(
G���V��_��kk�Q9V����㦴�����1ы�������Q�Sy���1�٧?hqKQ߄����I�;�1M�H��P�U���c=19���R� �%A=��}���l�Jː�>HK��[u�sɑ�~LR@O�}�g���ya���qީq>���� �C�OWP*�ْT��
�.�K��9�Mz:A���J� �nO��^d~����c��ӧ�A(���o������n�a�枈&��{g%�r�Z�N	۝�2�����Mӏ6�l�"C_����}�	��:q�[�.���C�G�����/����#������VϷ��2'�d��3%Eg�u��R!��Lԑ�$��͟�'�B��MG���1�� /E��_f�4�x
��4�D=L��Ώ,;8 d�[��Lv�*~��J��yyY�"��v�_3؟/al`�����%()���<*���"J�)y,ݒ}Tk��j��ZX"���u]
$���
M�I�<N�w�c�P��u����'��ʉwMEE�i�n�Fߐ�^������j)��["KP�_������GIќiE]-��b`���k���X�,Goai���򧈀@>�L���12�*�WH�T����Xj��@pۚ����gw��,�ȶ_I�34tvh��w���-z/W�FGG'�<��߇W� ��ﴜ^ijj���O$=c@�ȗ��ir	JI��eNn'v]g{x��}r1�z����|��ϯ:��W��g�SO��΍��_o,T�W�-�j�¸ZY���]���ɩP"�� ��6j��в޸���,f������V~���RRR
�bc1������;Y)�S�PH�[[��}�?"��%z�,�@)M�yv26��'��-0R�Eڣ�Ag�s�i��l_v��7)�P�Hʿ�
8��Y��O�}{T�.�5��}o��鋌� �{O�*s��?�W?X>������]�����z[�!�w�>sh.f���3,��q�=��邟)��^��iE����1ޜ�2A�Oe}�**�$�&�^t�aqDt�����^��-�cخ�޾�U��"�oM�~�zz~�#R���$	������!0=��DP�
UUUU�J��Ard���p��e�Ǟ�Յ����<�)A/MO���SQj%��N�G[�y�.�;zh�II��������+�gҔi�Z�Ҥ���<(Z�w���x��iUwww�e��0A��H�vm�������AK���i�3�D�X�޿��#��v���%g�w>J����DH(�"��@�&r(A��Υ�7h��K'�N}߾b��ڒ��H��� u�
�-��"��X����Z^��'u�����{޾�§ÊqW�s.]��\-9992(I��8$�����'xv�������Ǌ�H"d�n�9�����&_��9ބ�����Fr�b+eD�;�ܽ����6��*�q��q�Bq��'R#��*��y�o�\f���P�w_g��bL�!i�to{�)�ĳ�������њh��Cvno�u難?G�HW����2�V�cl,��4!��	�Ǐ5{b#\S��4Jpp�$�o�A�r�'W�R7�D`Y(廮������~L��VPT�Z�K˅  L����
�"������ɉ��<T���mɂu�֦�f�d�+3�1T�W��:qO��f��O�L1�esW�����e����BB�[�_���b��PT��/Sc�=��)��桫��f�~�%"b�`�����R�_Q�ȆZ�d�I[��ޞ��E.���h��u9:̷�Н�W9H���~��/!T���jJz:�����III+G� �*o�)_Kk��H���x'��;��猋>[~/�ˠ�����V��ֻ}�I�R���(=�~�n:
d��Q{�OΌb�i0��"���QV�znn�A����&(m�.F���c	3k룙��V?��io+���D�xb�`N��Td:�}�;#�%�c~{��OWޚ.o��9pN�a�6ri��x&*�Sܾŵ�C"�m������ed��Oc?���������Y,D�&���oף�8������9��.=�F[*����i&�ZU|2_<�!1�������2�x++m�6�f����]�/94��G���|�3�-�"�����r�� u2�ގ�N��������$�͟����:��p3o����ߏ�$p��wt�֓��t���%bҎ��ےP�����*(�C���*�b����8!)T@�ER����gIK���rkS)H�����������������+W�bּZ3G��z+1R���L�G�ͩ�Ϫ/]]�3�ܙ�����^�Wti),N��#F�b�X�̗���~7T�ADDDu� �gl,��?A.�;4\��;��C���������� �_�?�:C_Sϰ�#��2���| C��ڥ�����'��f �{,�BN~Ql�L��q�'�r�K�1zsz����%>ޘ�?���#x�
UdT�ې�j��I+:p+���:4Y�<�dw���(�?D�����o��ʈ��2fa�}
	�Lj�~��-�&[��?�Y�uJ���H�`{w��/�գM^��A�S��7��TLO�>=$�J�prRgg�|���ēxS�<(�`��9��c?�rH�͛��	�נWX�ĄE~\�2��}��]�=��~�|��2�r{�A$��5�JT��+�劃����r���((Vy�^Cq����u�S�Q���m�y���x����=h�	��>t�����[yI�y�/ehE�0���|�%�{��m�3��&�$�����?�J�Θ#ۖx}F/�Q7�e��ߧ�A�e�~��쭬�
���k�η��?�xL���vcs��EPg��ܗFT��¢㋁ ��A�At����PӺ�g��GOAs��Տ3�\ќ���I�5��95_wí$�`�0p�]�WE5����Z��ǯ�ə[=���㋿�Uy�����bR>T�z���۷oR�ºxq7�h�/Nw�@�(,(7���T����>?���	|MP�W���`&�g���o�����K�r�0���]y<c,Ż���^J����`�Tޏ0�>�8�C���mt]����F2��sM�[?�zBDB�%q;ȭ����(�����Q1|�ř�)#*�-s,ՠ���"���VJ�܁�~���ѝ��E��oO=�Y<��+*�#&���ƴ�N�yW��˦�{ �O"x�� ��3j�O)	���X�=�8�7�q��V�`���첀]tKi(2ƞl�Z'�x)�aަđ��s�Eu1I�J7�j�;<����:Z0��,��}%u����i�H�x�3�h.��z\@h�2Uq���r�C���Vzʰ��~�D!�znAAA�M2R�"ά���]E�V��$bY�6���ⲞVs�fIQ�=��?@b(���W`��L �+�����K,������[��v�J�������_��l������N��a(�}���R�4N��}-�݊�T\:v��녬1+a_���nF�q��z����  ��_����(a�/��.k_d����h�k/��QW@2�"ӟm7cr[�˫��Ʀ��r.F���������\!��j�V6/�"�X���Pv��D��,ȳxk{����J�D�&X��/|y��|2�Ȗv���05��o��}�<���󷶶8"8�~/;�7��N�|�^⾽�����:c=�ަ�ʄ䯸��OL���qDr]�������l�0����2�� �PI��K!z7�W2�h�N�j*ԞJ��k?~�h��%e����.T[�P<E�g׽���PN.X?���K�4��ԍ����hO@�6ƺ1���A���e�Q��\D���(����-���{1�N���s\���1��x�"+~$��y�5��Qc�B���pku��[D�����Z{'>�_~-}��ׯ�o��30�ӭX�}b�rM+P�fp�����M'���C���F���Ǟ��Jp���Wn�I5ڥ��\��D� �Nlm�j���\WP�v[�' �f�7L�b�ș�	wՁ�	#U�<9�C[5��S55u%O���l�W����F��l^�������rH�%511���	��5�ڣZ�)�:�y_fxh��f�D����&7���EW�,#0�������������7���ób��1����sJ����4�4�#��X��a�����o��QR96��kXgeM�N�H�J�x�)��xeϹ����o�qa�-� ���@�w.���������dѝ��U��s]�5}Q5ͬ�5�]�!��f�W�M�������Hy��t~������u������q3O�����fj�,F�e5����-���
��Sab"�>����q|����S�i�+;%ϸ�5+� �����l��?<�x�q�;ہf>��p3��mGp�q���6���R�#�����T��@MebT�<������{|�+k)fdם ����x�'6z�%u6��j��` �J%K�\W�k���F �&�k���9��E\?�=ʞ!�=ư��|g�X���^��|�i`T����%g�miɬ`7*�,F5]���ǘ����0�z/  �OShmm�e.��*��y�)5&%��;+��PM!ѿum Cɇ"�����{�6�c�������v҅�\|d|`
k;;�"	u��C��u	
L#�xXޗ���zu.� 6���I91��)qޞ��(#�`�[���l�9�,��"�5d����3oO���-NuqqyI����ʪK��pau�a�ꮧ��A�t�+�Rp�ոs�Kc���i�Vg?��B�&@6������X���`�HM�;?�k���k[b��;iƋ�9�3'�o�7Dr�S:rǫ��/c��~}����P����)0��/,\��j�|Y���j]�#*,^1#=c�8�"��aK,w� ���1����c >F���<�~hn� 9N��P`bJ�}��(�tf��&��1��ƭ��O�9�
�=�����ӁB��ճ�e0|[����C�v�$��vy(9�L�
G����\A�����b^�>t6��c%�&5f�9�;5y|rNNN"2~�-�\�!�\oqc�ݬ���:Cj;VŽ�O���Ĕ����0�C'>d�勼��É����!h���7�B�����X�g��|��r|f&u��5-�@K����퉘���x�u�jd�M��muI�Zl)����L�ߩ�)4��"_��ͷaz�~������p�&\���W3��������%%mK�ޕpO��@�������>W.�x�hm0Csl���]�u�?�o����{/_�lX��hx�����ˢ:��u����ُD9�o^�&��l6O�ˋ�-���%ip�C�3���ߔ2�+~��V65� ���8+���������)f���PE�� �;2���wgg?��+F*�^��gQKK����R�]C2��8� O��4ɥ���H
�s
���]�J�?[H[6hJM�v��_��(��/N|r�P��	�du����(�V�~͟��p(��Û(+��z��\��I�N�[Cl�[`7�� _�{�,�t&Ԅx�'�n~�6�Y) ��w1(��^�׳��[�f�X���E#�CW)|��eD��^�(MTDQ��U��Ѝ�E�˅���r,i���������rO��APP0b_������/��ɩe'7�7����wz��6彐6��i�b�����ꗺ�u��A�}~L�(�lC[F,u��Ս�ί���P�I�H�(�y�B��oG�s.����sM!~X���1h
�_1�<�aI�"�]���E�٘�����Qu�
��.G��F�ΰ;
���C�@5�J�x"& �X��O�8����!Z��L1��ff4�+>;Y��)�%W�4�c��/-��'CC����m���2�� `�/��U�Wn��8"�H�C?6<�t<����|vy}xy��d����r@�,P��Dh��3<̅\�0y���f������X]�|���H��Z?�"���lݪ�h�R�6/U4�$�'�1����i_X�f���	��E�׋pcu�ľ�����b�Y��:ށ� �(��~݉\���\�;��fll,�a��Suee����1i봬ɴ�kEf6�K�G�+}%�x��X��eeh%k�	{`�k�qc C�nH[���$��Dc������-q��z�T1�p!��գ�C����]�m"�^���`��L��"��}/��58׬jZ��8�Q��|�7?:2w�T^V�mq����!�XCu�t� Շ9?ɬ9�������-�B�>_-@ƃ*`I���Ӭ~~3���
MLLD��
�{*��k��s}6. ��s(?�;o"-�����L#h&�dt�/���ȇʾ���CjF�@K(��xUW��V�x+��OZ4G��\:B����Th(?�5u(2�������C����0<L�!�/N$<�&���U�q)2!���t��lq��,_BZ�oOQ��E�E��b����*�HL:� S�������A�4����Y�����4�q ungo䢚�9�xސ� ��̅Ȍ,8�*?E���F(�Λ��	�єNX���W����2���&GFF*Z}��3[�L�7�&�ߌ�����ٛ�'|���� 8��e��ȡ����B�2�����3T!5�7 �6��{{�'��W�˱��b��� ]@�r��|�_�lK]�b��eh��+*[O�� ��ۋD"5���M�������Mu"�Pqs�8��X*�1L�
ɯ��-p.����k�`c�T�j�+�ū6z��Ewc��2�_����l��w��"��I�w{}��^j�~��$�DR�vq�A4a��jv���|��d��L������#�I��9GFD����ro���3A���y�(^֒��kf�f��>~��=3�Q���Gw�ݛK]�[o�=��C��?n��J�o��~��Oo�a������V\?5���o���MU�A��q�-O��9[��*}S�05�U�������� �K��0*h�9g��1����p5��3�+�CuT�g�7Y:E����0gьC�fdq��{i��}Њ�ɽ�|~2m����L�¿ �Olk��� e��K�?V���6l����n�8�hp1��ũ~����Js�p�oB���C�Xe���X���F���钳SOMO?��Q��j��<(p�ݰ����`#�J��`������A�X��x�@���Ƈ�w��v�xݎ���޲M��<BO��{Z^�� �\��p$ZQܠ󆅅�&+�Fw
����3���`]����m(���2R�8૮u|?M��͎��q�4HR`��"{ii)�����|�G���I�Ώ�-��71�8��JV_SS��e? @��*\ �q���I�$V`Qu'��|2$��)��%\ƚ�б�yx�J3���!�]�o��c�{� � �%�DA�E.n��&��O���������9s����e?���	`{��$"��ܵ��A+�'�0��Q`x?}��/ �x04b��+.?Y�"e��a�ga	����kr��JY�f07`歭-gIVV��j���T따�����Ե��F�r"�|���,�ٽ}�T+|��>PSR��)wHG�hA��NS2����S��KJ�n�g�U!#˖׻
�x�Tq(ݻw�&#��A���S��6� $�i��>�qcY�7�;8Xz���|�2��� �P�$��i�]�o�Xı*#+��z�{��6�����ֶ����]�ّ��C	����v�ټ�>=�/�O{��uyՄ���ڎ7NSy���߹,"�!�jWDNN����|�@�,)N�U3	]��X�	iǠl�:'''+]tqKˍ�����w_�e���Q~�Y7'�d0�Ήa����q���-h������O"4]/�7��l�����AGҺg�������I����¼�=���[����Y�2�,			k8\$'v7�syxl,A\���*�xh`�H5������p��\�b�
���A�����Ʀ����"))T`����y=�jR���nt󋁯,�6oz��OQj�im�##�~z���"�W����Y(��$��-��B������s��51��VP����L���F	����(d^���<`-Z=o�k���k-��_\I�jn?cv�o�����㣭���1w8=l����6X1���N��+yR�L��Y�U0���0e`C~e�X���FW}��z|g��ѣG���$!'���j����¢���W!6I99�n����By@[��@y��k�����������h�W�Y����]���9�LS���������e�attt�Y�������6�G�t�]���Z.�����:�붏7GEݶ�������;9�0-�W5�J]�1���,�ߑ�����Q֡��"�b{{;�O(:���)^��ia�z���N8&̢
����f����+��ZZZ
k��J����>=�X�/�X�@X���^lC���I�M�2�����:P�<S��^���5�,ѕ��0�꼍��]}�8_��g�!�ƶM���WKK������uz_iF:Ǐ��ȴ��ȇ�� H$9�A￺�MD 	�m��<%�ͩ�#�vj4Z�W"M���7��fqrz�|������������C�J�\����q!~_�\l��Ӓ�+ԭ�0-��㣣�%�/?�����2ǮXz��E�%}������������/Q���~ͳ�U��\PG@�����k�� �g�$�����#'��e�>���bTT�^֡�/���,���ff����%�o�:��LC�{�R��-�n`�M�N��n�n��[�233�,�U�+:p_�&�3_��&�j�ٹ��2P���c���O���[A���(Qy�"8,	�*; 3j�֦�2�՛��#	m�c.��q��kM,.��u�,-U���E�>�a����������\�RD�4��7�?�P/*�{L�[�`�(����u���E��.+`��9�����s�O6.��V|�<߲A��iw&l��9��{ɭCS��:�	�g��ߤ���4���~Fmcn.�س%�8	�I�g��kBL0a��%ۭץ4�ov�� �NO�k���J�nc32J\�=82.ʼ�C/��{Wؙo}p{-�u��q+����_�T���y����'���Ffo���]�����c#q����z��?`�/*T����,�f�^��b]�2��B�1l񗁖[�����W�����[J�VX�2�*a�Hcn��5X� K��zh����*[s{O)i;UZJ��O��=*:��~��	AE�?&t�pA�5U�L�^Ħ�F�OW~gn�pr$��SU��oo_~6���l�{}��L�%y`��G`��T��Һ�����A
�[���"##���E�
:+E-��b̠��탍qU����MlZ��늰0��9���A��՗���S��Ƨ��::^'�a:���qbr���zw[��|&���I��5![�@�/�F����񱝭#4mL��KD+�i' U	�i�5;��~-rX��<1(���0���:i����i�>���9�,ɜ�>�x���Y&�~�|���i�S�%,+���m8r���(x&�o��v+���5ətc&}㝌�f8��0���D�#�T�H��**R;�NR9���V|&J��|?���+]۟%����K3���tbr2:�***hA�Wz̄�_WS�����J�����'B���V�r}R����L�U[�+��\�{�2bzxǫ��K��-+��ݭm6����-�詟MStUZ��,EJ\F����b�׽�9#vUMP~F?��d��fK���b�pZ���Sq��$�_i *�Я%/Ot
���\��ܒ��g}64��OF[A1�)0�~�������i�=$�3_�J
�+��_�Dn-e���вS�%僮�w����J]���ףǆ-^��8X"����.*FM߷{u�G9eeo �Cz�Cڑ0��w~|�����k����}Q�8`�Fss�7���P8f�&���:�ۦ8ݺi[P�چ��Om�6��C�X��P�ɓ��ڸQ�6��#��ݬ���7n.l��ܔ�䂷��GOe�p�:��Oe~���{@���K~n��g����\�b�����J��B��jBOJ%�&f�<8\��z*}���>�}����G��~���YԘd��r�k✜k��6�Ǜ~�NN�����~N�~�$s	q���s��,T�C�	N����='n�ſL;���D��r���+G �<-�a����?*��k�=�}$-'��#��E>������V�Y���G����lnC����J���ܵ�4�����=���������%��4�;C��&D����_Ƽ=TF�p|�e� q�岹��r�Y�g�r��|��_R7�0GUS|G~�4�A�\1�kīqm����j��^C���A�����>���G��(���İ8�+"��.'so����������j\�UUW��,=h$Cg>��f��Ը����X�r���x��v|���|$�2�qZ%qqXbXR�%���k� �m$�'n�F����}�n����n�>m��QQ���M�[�﹣�"��Kj���l�2Cͳ��Z�Q����*,���r�7��>�?ꛠy�+1�/ F��C����^�aeG�Ѽf��r�ZB���Q�m��i�;f0�ظ��\�+���Lq�OykAp�$<K�@	�1�NU:�qgW<��Zߟnwh�%ŉi���H� '����>4��i�X*�
~������}�/�,G��$�VZ�e1:7]�p9c��V���o�ϩ����m�]�:QR/+ܛG�d�=��Wjnn8���gf�����Ȃ�ֱ��oʜ۪Y|���%>��j��� F�le��)��z11���x��l�!���5��_+���PZn$�|�0	l-M��zlw��b/w��L��xN���~��� ��[��R�H<c/9��X�!���"��??s��g��	a�pj�K�C|�,5u�2�0k�V�ӄ�cGU�9Ut���j��m�� ����;����Q.��ц�7V��W�r7�\� �D�P�8ifTUM�J8�Ԡ�hu3'�|�]dо����34�w���kɖ��\o��b0���]m���p���C˓z
�G�������f<�^"	�]��$���k|��k���A��_g�H�ޗ��b�d�Pd���6̿8rr�M�0�U%�ڐ#���`\���ܢ�]�qVX������*�6y��	I5�����5P�E���<A�q\���R��*���,ۺaB0���q;�}wm� 2#JY���NS?��+���k4 }r�s�*����h�8��Tw�)�Yz�%h�3(i绦nW���Mc+j,o!/�CƤ�K �R��<9������'s�k���1M��DG"L�h]\�QX�_����3G�Z�[�s��=���F'$�� +�:U��EG��m��`���+^����v�KH���|�����  ߔS˰N!�t�1�������u����v�_��xii�w_EM
.3N���U�b� �	>�wl�	99���yz�o��Lz�iT��EM�@�t&�}��a8��Uj��Y#��%
I�\��E�ٿ���,3�;��(0���}t��Eoks�ypi�) �T����⽃�F"�Y�Byaa�c���F�n�>�}r��ip�+k����J%s.�Qɮ��]_8 �<���z��v�$/��7�u��
%ٵ��ʌ��ן!���9����
��TqGcYT=�m�i�k��?d�X�>49��f�����݉qڙ��|k������2����0zn%n�VK�4���i���2B�qI��M�ID�0+M�&�T�X�������X��jv������܅����^�����:���y�����AgU�߇��W4!0<�e��V��K�5Wll��Aϭ��"Vu2:�Χfp �)����yjZ�B��c����T2$b�茕$XkݽxaW��("*& �Qm�u7���[��;>��X3׷��.Tg���,_yzN7���uV��C��H��[��t�I��R!�����ީ?�������>��O��pq�g�#�NSYX�	o,Ui��Q��y7�B�$j�_4lr�~c���9{�~��]�%�+�6����*$�:9�<�Z��3O���ڳ��E�>a�v�����;�xtMV��D�-��$A3u��u�'\�3kc�B�������9s�tTݺ/�f̗���4�X]����le�P
$��ou�;�z����U�W�w?�(�RG"��[��П�QONl�}�򪧙��jzz( `_fx*�I�<y�ԗ����e���b1�q���lj����t�R��Cf��)����aLl>�qV��A�[s�Ĝ�;z@r?��KJf��)��#��%�h?����X	j���b��U�+��W-ς��ɸ9�猐�0��U6�Yt�Yt�֣�"&:�����g�&�@��Y�4sWHl� �A`���d2WL��,Ϫ%v�F0&&��$#!��i�ɕ�==�q
EL^�"u��ۆP��0�-	�t@�u.b3���n�<lv��P��PO�
�ҡ�cyI�\��peeD����|:ҫ� �ˬ����j^�,���4�h�cc�km1zI�R"/e�εxq'p���{�]k< DL��ȱ$�fcw���b��
����o�4�����K!g���ʫ?c�%���DM �J�5c��@�vI�sA�*�?C�O/��v�-��cd@��񿎮;>�/q���?�0��/��CJ�?�[��
������"A��9�7�7���C�ߐ�7���C�ܺ���0�i=�w'��� ���������;�G��?E�7�e�L��?PK   �<�XT��"  T$  /   images/53cc934f-9b11-4097-8823-694d19808ece.png�V�W���;i�鎥YBD��n�k��NA���f���e�%�}��W�/oΙs��=sg�|�Q�@U\j\��jJ���

�(6�U����������u�N���7���]�yz[�[�x{{��9;xXZ�Z��dB��QP���+)��d�g�|��=|�͋�PT�f9+`4�P�ЋQ�[(o�>_�T�1��tj:촶�[���)���t�������O�Y���������r*����ן��j��Z��v����	����}a�JJ�,�����|~݉�ػ��qek��#��M$찮�����!�=����:���L���f\I-��i�=(����g��[I���Q'F~��6��;�c66R�M��~G<�2��}F�D%��~���ڴ6h��;�"~�f3�K�M�	����n�i�{�Ź��1�3G�A�m�b�S���L��F@̩`m���ԓhsxC�[�*���ja�b��+�" m"0��Q�M��O�x��_�f�㣹��nU�0���<���@��D���;�l�����3B�JK�P:�\=�>�{���R}<�^\�a�iiݶD�<䲡����WRl�Fյ�t�ɕ���*�7�R�b�<c�iN��L?�L�|=,u�|X���K<���5/�*�}k�S�)rߗv6�펽�E�P�kJ�v�_���h�e0o��%�H�"�ŭ��,�v���˶�z������kB��&{�+.8|6)u.^��~�rv��8p��y.(��7�z�\(�S�-z��?��T-�0Q&N<�/ٙ���i7-q�!�����{���I�Ot�2-�MLKYՈ�Ln�SI��m�ڱODsO\��3eZ$9xzeU��)㚗�,��M�pN�.$:[Z|='���3���)�����fb�ѩ���Ԣ5Wd��1�4P5�b"��Bg�!��D��A��$��'�fS�Wn?���[�+�=�����<��&?���\,���-�%&h`�W���#��9����ڄFd��>�)�ק��ݽ2��+{�a�����w����ӺS2����h��-w�̾zG� �d+���#c=�G�~�Wؾe�P�+n�����f��G=���Q��F�V�0�n>���DP#�Q.����ųN�^5i������Qc��-kA��"�����4J	Ĳ�[���k
d�I'��%W�k�k����@��b�)��H/L��rxg�CFd�S�����uEt�HEx�3D1�pU{��z]*+ޏ�Ցe����*�u%�9��	!_2)����RhY�n?��q��	46��W�Zv��T�+����i	�)5�pc�C��\ѐ8mZ#� r7{�M7������K�7繥8�I�c��n� ��:z�(f��6,tDODw����r���{��%���m����W1\��-�4k��*�"�قg�6��hp���Z0A4c�]�
E�ʩ>�8l�y�nT��S.?	���8חT_z}7
�Zs9������F�|&��焺�~�	��x�\�;���KI;Qj���Z��x�coSTM����m���H��mʂ�U֊�wn�l��]���^�"�Q��p�L��i1�*�{EX�pr�df΋u���erG�Z�k� ���A�ջ���}�pf��`���������=�h��_����	C�W<�ķ\1Nz�K�'3��U~T�0��%������u�ڀ��Oo������*���V�6O��ɂ��k3J�8�'��W	�5O�}'��^������g�$�����}���C���v�8�S	��?6����;"��C�Vn�Ba�����H��1҄�-j��%ö1���2m�D�9zˡ3�"Z1'9���-	
���v/g�J�q��`QK}hִ=�{� ��fTM���*_�0?b)�Ω�wMkO@&�ut�mf*t���늾0��d���|r6>m�AI�s6��'�-��8�����+Y��������0��a1��"�(-�͋��5����S����9 fOb5��� @����w>O?��`�~�2�0S�ؒ��1��`(L�'��K���t��?�*�K�,�ᕪDbF>�Z�F��`�y�;�A��y�tj�XXja�\l�)�b�=/�P�J��2V��56�Vk?����} �Շ�G�X��T���\��W̯k�;����ԌL^�0��ŏʥ��r��/0�Ai��@^�0���{�WM���[U\���h� s��'n<ͻ)�\Ǒ��t�b��i�H���Zf�"�9I�Q"O.�,ɗ�6���f��t�ĩUm	j߱i^���~��ïs;��������u�)�ф�]]�m��͓�4�/Ikf#�b����b��F�wk,U��D|}��>���ĔIX4�w�4���ENQ>��ShJ�MGGڸ���.��|kI� 8��0�r����qH%h�A�h)��[���)�9����F��@Ey^��k�z���^��}�_A؇!�I�i�RI�\d�(�+�#ʏk|7��V����������<P���bfG��Oĥ���L�����{<�k���^�UG|���U�y�9�����O��Ah��k���q��7�K��ܹ^�Yps��m�3x�k����#ʹ���~'���/1�yb���Mfv��9Y�����镰B�3���5�=Y|�X��C*�+�}��A/�|�\͈�%���L��n�K���~�8�A���ƨN�D�V�Ģ>�чv&�ÿ��`mjg0���?k��=,�~[_1����	:U>U�p9s^j��wa:����� �~��1��+)c.pq�Jt|lto��:�m�;�R>�hx�\�1�;��,b�y���(�*_����q�P�ﵕ^�W@��V�E���SM������5L;��ި�Y�=�ò�3�-��AwZ���L�v��A����m�D�ͳ��V�5�LV����2�\�$�{߁$�P��7���l�"��o��a� ��gfA`7L�p��K��� 6-'�7����I���)>u�����`�]��]�U�>��s�`�#02�@�;$OB��>ɩ���:]Q�t?S��<�E��N�a�UŤ��!�Ŏ����=s�I��y2e�?F�� �_�*��L��=,����;�A|C{� ��m��|^u��a�ӹ*sg��Fʼ��08�ہ�Rd<�} ����,�Ԋ�~���A`×=��ˁ闑o��2��Ϧ	�R3~r������1��{�9}�>�P����f���^	�,O��bg�ꎫL�%�X�e�k�Z0�+�xX<����7������͢�c��ĵ� �9�s"R�^BOXpWf� >�I˖����!d����O��Mr ���Н�F�&������F�D��l!�|���*t���;wZ:w��;$�e/Σ�R.D��Fl��:��st��r^M���3�q�i*C�3e��z�w6�v��,��K��g�M�
��'��]����d�j=�do!��\B�oGԴTM�߮��V��F��,�?���q̠4A��z�ƀ]֜x]���gLFFG߷��W�6�;ʪ�&�ãA�`�A7(�s{�9����f�8�uP��t�7�|��,�ĵȃH�<����w�u4�M�������\�_�i���!C�X|uyr��59�"����Q]5~���'�c;��4#�
t���o���"�4�Ee:�/t�S�|�IJ���4�G�gᵕ����1�\�ч��o�5��%�t�ة�3����'�{�
��o�˦��x�0F��|Һ��S@DQ<�^�P&����tih0�T,�����L��s�wbl,�0��Y��Z@��S��M����&I)V+\���#M�/əϮ�ɪ��6���9W��]�Hy��tnC����U�Q		L�o1G�7�,!]�Z.��$T�GO*$BLP� �$��:z��}���c�98���S8T�1,�v
$ �kn�Yh��AF���$4�͘;�;�Z��#�mUznH�^G�}�����ʀ�����[믔�G���Y��P9�|�ڙ_�m���>e:K�r��I�t����`m��a�z���>9U�~��!�W�mv˶KN��q����L� �J��:�����o�!���[���x��\�UCS�5]B^a-�p�B�ԗ���m�h��'�.�h����Q�0L�ƕI�Z��Tr���h0���ϛ�$e���7/VH��8]�
ڻ:����v�Vo}J^��/�B?�	����Y�G������L�st$�P[m�q��
y{�RYR�Njz�������K��L95n`5�sD��&���Ŏф~�ʸ���ߺ9ǻ#�b����q>.d�c�X�("�P-ç	�d�L�~B�8Gz�cή|;�ƅ�����.^��u�)m�̉9�8�k���p�^��X~z�R~z�$�_J5B�}�� bH�O7�$��~�b#�Ӱ�$>w�$�KR�|.w��=8pr�`8rX�D*@B��m�ON ���u�ܞuNb�!|��aHȑ��co@�į�+�_5�0?y��S�M���NLi��?l&k���,"�~S�u��x�2�H�C6702��J)l��]|��qO|��F��Y�@�pZ�N���|�yN�b`��>Waa��/g���0M5��	��^~k�%s�2�znf�T$�_��Tj_'�?�Y�������o5�FQ�b���C�7e��$�����~���08zǘ<'���� ׍�c?Yj�����? �4p~�>�`�>YӶG�w�$aaU�%挀&��uN��f	e�ݱ�E�Ԫ/"�߸w�B�X�̫����TX�)���4�<U`;0��=BX,�Ix�:+�s���p�%��)���Z��$����
��g�k��E�b���5��x��D�^���a�+�v�˩ax��,�&�����{J0��)U��[�R|,��I�F�.}���&�^ ���̀�\C��^�vʀ�5�R�����r��%�hU�{Z�@wpx�4��I����6&�v�p���9�K[���P'�Xm�.#kQǌ��1b������MJ,|U��O60T����F�B�g��	���H���xYPOk�p:rlE�ϕJʸ�����u������v'V�˛���r+O5�ƣ�m;��1}�$���?��Ӯ�����@s�} ̜n+�ǫ�#�]5L�g|v�©5���	E"��n��1�
��ӵ,�_����-ת��������K{g$�fI��K��e��<9�Ksa�ã��=����n�u=��|�߂I;�π�C@y���l��ʊ����N	0�t�F3�����������>d���o1������p)����|��WU�	o�f3��$xoE(�?z;�(y�#���]M�s�M������8�(��Hx���/��� �:��Y޽T���bc�c�_Rі�a��<�bad�f���9����A#5��d2�pd�Q��w�cO�_�iM���F�O�w���)R��07�b�����V�R�~�`�P&eH��r�!����*����2�?��0���l�{l5m7ȭ��V��'�ʪ��-�����s�����M���]�D�T5������V����4���;]%^�P�(��f�l��@l��e��O��ʅ�λs�����!=�Gb�i���_�0�!`.c�^rkHx�V�_��O,�qs�{u,����ጶ'3��~�{�AJ���������.+���v�������v�Z��	xKϡ�O��!@XiV��\���b��]0�BM;$���?]d��"��%�&*��Oa��f8"
#t�_�Et�#rԴ�Pp@} ���/C�㋚��fV@�.�v�':)ZXfU����MTu����2�^lm8R��o�V�ݑ�K@�i��h�5�W����[����Vp��<����䆸[���(�2�	�ר��}b�ƛ¶�cƙZ	���ڹܔ�&'^�p���L�ΖoM��p�`��6K��$�:�0J�cC^�:�6��QѷG�W��!�W�yr|ߛ��ۧE���Z�7^㘲ޝFr��S�S��.��7)�3+`�o��j�p��^�g��5�w���Ex*$�s��4?"��_��	��A���J���������ۊ،�CD����f�F6:>S	���d����#`�p�����J�2�i-ʝ�G�a�Qr����C�f7�Ol�zY+��
�}M'iN�$���P�k�:/�?l��Zq��}n� 81D�a��v��Nr����4sU���=��|�_��1����5��rcsݍ�h�1*�*l +����V�߼f�'��mLƮ��D�и�2���K0���LP5G-`�}��&�����5M'�0Wԫ��+��dm�_�GT�F㬖��OE�	��������Xel�OiDX-��妙�1��b��B!�{j��-�:��]�rƤ�Fǅ�_��/r$xتы3�9��4��'��I�8�[L�	�C��6;�#322 �H�6���������/���A�h�C9�gMI���p�F���KX�����],7R'�I�M�����;��H6��+�L��G��A����(m��+������5�)�����������h�D�˽w�G�7�n�,V�+�ktR��,����OҭD��g������}�H�lA��pf<ʂ-~X��-�^CQ����wsSn��	>����!9��"�&��h���܎���{��^����Bid���R>�EG��Ex�K�E�{��$�O��GZ��"0Wq�p}�����g�Rk!9��7h�Zߠs���ǅт�_(�}�	\��*::;:>�!dm]\TM�Ա�^<����w���<�&�Jv�ȴ��\au�:�6�ⴑ�֘�BJ�9���`��b���x�}��sۊ��A~��ĳT���9���)첊9�9��w��� ���Y#At56�d��VW<9�*�h@�B��NFQ�Zr�C��ܶ �G�`�.V�7�� �뜧���F���R����Cq�~��z~������,�>"�D;k�teW^�q|; 17�)�|��t?���P�M��EbZ��2�n=���K{��c�ƛl�<�,��FXԭ��� ���Z{��&����˲��T�;�vg7�(~�IrǛn|ߨv�|�bDC��yf��c*G�r�]���?����Kc���jcN�eM�[~�����t�pq`�Iv�]�f�����N�U�\��ЀN�.�n���6�9�5�Y�f��<*�H�@�B��T�q7�5]�/󂖏�V B�F�h�2!|d�m��G�O۰'�ޗ��GM*� HInP{Eeg �K��)��µ���XP����{��ʬ��-���/��B�E�ӛ2�F����._��+Zu;�'[ŝT_��=��g�mjQ�%#�f�e5�������Z��ˠ|�^pO������1.�7�]�#�ѿ7��~=y�[e�i�m(�p�ﵧ�w� /P��<s,$Iָ4�!�����rW�u:�P�y�_�G�=R�u�gs���$G�[����)Sn�3��%�"B_�8�� !OzWj��.�ﺞ�����ipxĚ�u��\�;�z��w�,q "7 �������(PCKnP�� �0m�Qɚn#�뭒	�#��V����g&^�Q��C�q���T}y�	��qA�LMK�~}�|�C��Ua�Ύy�jQh��?�{�)�,�ucn�I$������}��i=6p���^���:�����px'�N*"�'�Ic� �J���d�e�ʮ�����be�Y�l̞�E���Ix9�r�/r}sfm�s���3募��|v]��6P&}.au�d���X��s�j]�R����W�"���j���u���.��%�D�`��S5��>��l�D��'s����H�0�'D���;N����IpX�ʳ��1�&'�����S��.��F�pk�O��]m_N�̖.vJF�=�2��f�ga۶�f�=p)�o���W���n=��$�/����UF>�<ސ	���΁��boY!w�D�\L��輽�hqN�m�x�^w���$Mo��ִވ��|�/F[�5�%��Mww���5G��ko�cBp�KP`�|}4S=�jcU�|��"�xn�����Fz����Zh���V��&�n_�DD`��*JQ86�E�u<��0U5�>�}���tMBn�`�����L�����jQi�����P�)ؑ^��Ǯ7�.�|ܝUF��?�=6;}K�<��;�^��F*,�?�c}Kʏq�~SƝ�b/�/0(o7���ز�t4s����5Y�_)�4��'?h�P��e(N �,zp�R�j�@�?=	���$�v��vya5*o�G�M`{%���`(Ԕ��/�#yJd��5������fL��e��8�/���Ӑ�{ys��y5T㜦�#���$����rC��C���Mս� Rl�7���qd��y�O��Dk���q���=��(:-��SE��x��2��\��}����7�F�r��Y��m�4�{�I�W�!���	ggKA���=Ef k���5%5�� q�6㺁f Z@���%w���[TVZ�c$
�Hn��Z��x�T�V4�PK   �<�X��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   �<�XH�:9�\ u� /   images/5bcf48fd-3e7c-4271-817e-97f3eb0e00be.pngT{XT[�7����t���tw������]�tw�R�1tw� 1t7Cw}{�����y��G8s��k�������(-��N������A�,�4�ݑ���O,q�Q�_wm�}��>������X�)�"!�5#�Cn5��?$�V���4�sж�Grpp�3�0��նҧ��1L��!!=C��^P�1i{��N~��d7�A��W���	?�<�<�qziX>}|\b���#DC�(셟�����@\d�z��/3��v�?i��KD�"y?�@�
a��^0O�O���q�{v���/�[E�'+�UH�j[��Q�r�d��~�>t�ɺ�s`t]�,m	Ѕ����G�y�S��O���KG��J��!:j.�:JSg�ы>��P�<q����f�6��`9�|FM{3DpM�N�G!���|HT٬0'{����X��}���Y���ꗑ�C&(�^_��������]��O�4��3}j��'pQ�N^�=�Hz��'�`�E1��Eo��/�s����$Ovt��������-��/ɻ�^��A�P4~[ѯ}�`
����U�,�M�Z��A_Z�3Id[�]��M"�z�q�t�X����,B�y��s���䵆���N���ƺ���f���Rv�1�54aW?���ȁ�u����,����m��ej�ԎNs谰N�Ƭ6y7!=�[��oXk�(�Mw���۞�Tź74]7={6�.��s�<�J���8!�u:�Gɀ눴���߳&�0�����Ⓞ�%�/P�a�HRR�����!�f��ޛ����	MVZ�R�����a�A�M�#�]s[gJʑR��Dj���[�6��&�y,��n�e��p�$�Z�Oe���}3T>$<�W���XW}dH�FMk����Ɣ���%�}(��pȉ��u�&R�ߌpg>�Ki��%��_+y�4�
�FB����>v�psȩk$4J¤*�"��4m���MX ���UIj@��c��SO6����d��GS<��l��2�-�/>�כ>���Y�%�t|Rz�-� �p3iA�I������D�z=q�bn�T*��uY�t���I���=>u����Kص�`�v���LK�	���7m
Z/�綟����t�8����4����Pq��<����Eb��5�`4�I( ���_�~Yk���sSAQ�l�zb{b�����L9R-Z���9Y���q�8tyf����O�9�S	�%bR��̿������H���u�޽'��ﵴ����ppr.,.~)*�G��Ш���������D�������]^֋����|��F�K��|$�p0�nc��J������*�$�S�L�2������g@Qą���.��'.W���HF��Ϗ��˻��W�4L���Յ4q�������?�r��@*�4V��chݵ��~��O!;���	��L`5��H����.m���U����ł���V�趶�t�}�̆���T2)˿s��5�-��]>fTH	��qb���9���>��$g���<88gH�K��܂�X-N�wο~����D2S<�0�����Ô)����)��&��ɨ7�f,�b��}\����l@ݷ���I���f.>�%e<]����sQjܼўo�~��k٩�/��B��8������Й,3vtv�ۼ6�_��N���c�xxx�����5d޿��������7��#t�pD��zo^�u���n�G3(��]�-E	�7�lll���zz/T�A�}�ߜ�V;�K��Y�z���x��K>����r��ˏ�qd�ѯ/2��eC�'�R�|��N��9KA����]���C-d��xL�x�����hk{{���Ooo��D���ш��dy��TE�˩�yՕm������I�m� .IЦ9����PU*-���q����_�����Mu��/P�,���+Ҕ���+y�,�v��}�	�ڲ)���h�h���ݿ�xuue4��B�����MY]]�=�xkPd���VmӾ�����(�q�S�U��wh鋫�"`3�٢�d,��m�b�M�Kv5
T�{��a%�h�n�O�D&%'�󺰁A����ۈ���k�������.Ov6f��s:\U�1y|^�P�;�s�D�~`)��}L�����FG�G�(x(+P�'O�UZ̬àT35��ﾡ��-Qnt畈��_�N�u�{��Qe�D���'�zpxX�S1U�z^*��J��XY1�r٥)im�p<<<��*���fS���1%z�O�S��!/�I�] ��=\�mu���u. @�l�ܔY�	�&Am�$��ۤ���������@23w�X�h����@�q]���7jH&��G��4�o�/�����)5$������_ %k���j�ŀJ��:���6��$9 ���X�>�ȿ3U9�>��|qu0U<�N��;D,�1AH���9Ϗ�r�/Ҩ�̡��:Yii�.�6Z��o1
��򔔔���.u�&�f�T����≄�Ik�?�O�g���w|�rs�k�7�\f>�0�H*��Η�nip�k�興�7��|�_�Ǩ{/�˞���0�>�kf$��"�WV�oo���~���t�LoS�+)�E��0�4�-b���ˎ��xٸ��9�V���z&�Z+���Ue�[�H�8�����B��`}�ٗP���z��RѶ��.����^��d6s��WRLu�����b:N�����R(���'>>�F�"��٠�b���7h���v�׶���؏���^�=��hH���+ 3�����H��1���_x�__�^�B!ָ\ۙݫ��_"����M^�/��&���5��%qF�b��ED�@H\jD��s����LZy�!Wœ���o/�n%�s�x�V,��:�_��sn�P�A�|q�p8�F]�=,�	�`�L���c�(���/{�M> '�+, �	�n166v�9_�L`��#��(�z�ăH����w$�V?�KܡU)Ӛ�s"��j�ԑ�9��`2��:��_ZR�|����?1�{�z����'���GZ6Cj 	02�J�`3�(��3�x ۆ3%���a���Xq��j�t2����8��h���8`5���œv2 {������P�H���W~O555��Ԑ�NO;GG������+KmC�w&���SL$n���ou���i�9n_q��w�<�2��N�&�����f�G&%a
XXЍi����on��I߸u�Q�����z%���L�J(�ItH�a"i�˨X�Z�b�u#���J4xΧ�~Ӣz��U(����[�d��@|���0Y�u������@�|��������0}�BA"9�aC!��D����aj�z�����O��c�5��(m�E���Yj>�AI�NR��IӢ��)9Y���5�
p�������X�PF���o?�^����'�Jl�F��j�.�@e��Հv!�0W/I��u���:4��Ld�W:ZQ�	�M&�Mq))ʿ�}�;7腂�a5�ԟ��!�g��X��3rrrh�uf"�auQ1� 4ݏ����A���9�_@�ߖ�Ek$.�vW��o�FXLLG�7���?�(1qq&��ԃ�S*�2����J�<����@27!�;���'w���d��Za#�ݑ�{��\r��q�x�3�H�r��ݽ�I�7Uan6SM�q28���������ρ��~5�����0ˇ�ﳆ�:
"�O!�ā,3h��^�^K���z�ku;�Q�a�G����o�\�z�T�Bӯ��rp*��ͧ� ���ݑT݃���	�4x��cx�ED��Uʌ�m]�)`�� �[}�D{��qXB����:%j�J+�	��VY�κ���r�SPxc��Pa1�S�^����­࿿��]*����O��+g||}}a%*u����!+m�8���Ā%|DL��ȿ����.��V�S�.��c����3s搨���҉2�~�A����ONNN�j�MA� ���}���O���r��9�ӆ�, #}�>�t��R@Z� ����;��q5ސd�i�J�Ѐ:@�w��0qG���db�X_7r>�R�?佴�C 5u���3�� Bf�}~2e��9/��V��f�RqST�ǔavxrb�=QD�>�~=��\iA
*��7�x��������?���CB��<0}�����>2.����ݚ;h ��J'�,%�	�?B�qc1ɠy{��������۫{}qL�R��9O�z�����(6���w3,��J/��oX�~#;5ƿ�!c��r�rc$;�x���/��D����o[��,�%_�=�Qe������W�� ��Y���|�c�>�lhh8R
�����M$ྰ�DS��(jYZY��Po��|�i�OV�N�&�����P���2����s��2��8<Z���{?U�߂I�6y"���?lO���u9�[��1i��(|Ĭ߃+Ǽ����\@�T��NW��x&}��i��7[�
�S"�Y4ݎ�"����, ����^PG���Q�Ĵ�$M��>O��R}��Ӆ<J���q���}d	[4`8����g"�g<>�ݒ���5h��{��.Nw)By�9::����F��s<_��%a{C�+�ӂPO��}"`� 	ģe�����t$�8�S����§����2�fc�},�L�F�?�O|� BFȶ�<��-�e�!�	S�#��h^-�������)����,a7���<Beɤ U������]���	{~iIf��U�kDQ�M�����JȈ�=�Qw�X۠�*�٥D&0r��5���4�5Q�N�uU �IWK�@�d�u�׬��t�h9[�D}\@�3��y��D>�t��� H��`��\�o������� �P�s^����7���x�`�����P�-�]�x����Z[�1�pT�Κ��͋[C}��e�h

l��
LL� �?�8�m*�6fZ���䍚������3�u=H�釩�/����˗/��k^4�e"L�	J,�B�gjʅ�B��":�IH���]���P@�Az2خJ�ѩ�����^+�m�Ka��� ;;�=r�㙱�)�_�4�emo��?��Z��餷��G�hM�X�C��S��}I�{h�JEKXV&ypH�=������3칐���z�'DBH�UDђQ,ФH��2�4�����p���v������j���&&��t<�q�ջ8�矋NϨ�<Y�+���r��z��`^T+������B���I��9�-o�CM������E��=�tj�5�*�V �@�O���k��N��M��{�" i���"�8�kxJ��@3�@���Eɼ��ϟj�p�s:�J�ZՕ��6:�m(�-����M�i�wP\1�yo�������i�32� �T�7	���]�_l�}��Uu<v�>|X�7L�H�,Mi����v�L�c��F&F��Ƨ��b�ߔ�7��<Q���F�/�8k`d�(*"�4������K뇊ѳ�/o� FFڀ�l9�;ď�px����}\Vk
,
�	.�1�R`� A��6d�"4��p�|�B����΃�^B^�2�_��`p�гCO�w;�������?$}� ~J�(����Y%G��/���򏩨:w��
�<��p�C�Dw�5,�:V�N1W�H!T:�?�Jt���u|��������Q���e�Ar��Pt.g%`�RG�Ύ�vm�6\yG�PM�BsGE���-�=9�ZS������T���b=�n�ר�v!�U����j���2���,w�#*����>�ټ7��V��?�d
O�F�s<�����`r��*m�߲��|>�8�����
���Cd6�dy����0[T�B4�#W�~l��]\�{��2<^:Uj~����:\.�(,��6�)�����B�{Z[� ����؝����;�H��lX
D���&�@� z/������K�Sn�] ����Cw�O����U��	,���>ڿ�pjk���m_��î\�yа�W��3�T/�M-ZX�g�.}�ޗ�] ���322Rw�<�uk���}��fx��9�b�?�񰣽��n�P�Ċ��'B�����&Z6�f{߹�o�+)�j��r��|s�9������e?��q�E��������j7U���Zj�%r�@�~%���������P^�^Wm��Ӈz/>)}hs4O�k́�]\�T���n�iYm�H��}K�`���<z�V��x�Dl$����Z��!��\@��r� ybiiY���d(�ռ Pn������� �<���n��uZ̿�L[[d��VA�}rY��:Ŭ۩z�F�I,�ZR��Ǣ��&C�ϛo ��,5q�ſ�nX|CS�S�����SW�Ʃ�Tu9�^h��/��/A�;�0�А;9��ZFU�\�69B�pvg�\���Dcrtt;�U-�mlJ���hX~*C
���l��ULL{#�r۳A޾�S��@Lh���J��� %�x�.P�U�r��ttt��)���/��ZR�%���CHI�[�a�p�����͑�>��*��rt���(7�ZI�2?�(4{�4��nkOչ,L���K7���B�D�Hp�����E�����w_2 ��և�i�jo��|.)���|}�u@J���oݏ8��|d$�ġm���n�ި���~
���F��R:Z�@�SR��PQN�+�P�"�F>`�~�t����� f?�~��$^�^n�D���,ƈn>�&h6UѿM�G�"����tY[[�Lqm�,��Z�o��+WJs�1)3V�{l�wr�P��n�]oM5q�����؞� l�����;�o��f�JU
�O�ꎆ%�צŽ�󛴴R�9�3�X���L�|�4H=j����>[_;3�a��h�� [�E;�l������9�� j�7Wŗ���W/�����uk"��Ru�����ʟ��Z_1��<�߃h$�7e�x{�yE	�B����Rk���xQ*x���}ݎ m`�|Ǝ�%�L�ѩ�{�̫�sqC��:
�0��䲥8�
e|��J���9w��1o?C[Gv5��5����h=[��Mf�8�ӯ���������X{���K����r$���<
U��ޛO5+++�ۦl��bW�K�555��d�[�a圻�a�eȤ�pڴ�g��}�~�JD��0�����g\�E�g%�L?���f&�L�h˛�A����`��(��	Y #i���G�3��Q|��NS���2ᩖ�E�0X<B���_ڵL[�>��r�cY���CLzq}fT@����2�G�j��œ;Vވ�5�`�S����v`1���F����HRtclXT�)�)��R�j��CHD��x�X9�.���G#��3�]|7g�����|�A��9|:˿�<��K,�FY��i�7�ް��1��LG7P֐I�[S�2��uW�Q�Uj���f�+&��%d�P��h�[� 𮺽���hi��F*@����r����j���s���g3OP7pT�sG���@|b�������R�6.�uu,�3�22K�]x�,'ˣ�LNv�R��e="!1���X-�$[��1�UDIa�=��o��d��z��/�����:�0�֗̍���d��������tD(������g�]�;(�T�)w����S"6���Z8b�D�Hc&̹1:6�s�W�9 &SGsn%�fG�%�"VO
�_c���pK��-KӮ����`���O
�̆���]��7�q�B��ˋ��S����&U5����o����7�
�u��E}au��"^�6�)����3O��J<�A&����&�<j}��{��,,,�Y1?��:�l�Ӕ@5]x�ݎ��o��"�';S�O	�%k)�����F�B�yC����UX��]�ޢ*�_����MT,]����� 4�RianT����Ͻ[��4���{�]|/ﰷ��sߐ����R�AH"�����63���; FCτ��Ҝ�<�dNL�.'�M�Nj�Ob �M��vl�*���u�P���3�j����J�౳�� ������z}�9T�oS:����� w�wֿ�"��d�m�����p��������5b-�CK�F���4+��5�>����g Ps��(Mл������+_��)���=�6���|�(���%T�}����q���*b���vg�5q�L�h!d���EGM���|��nEZV�ܴPe<�ܶk�DQ�[�Z-�O�������ҥhE��f�N�6����>�W"A�ame�sZH�*��ې%s�f|��Y��Ҏ`� ����w��%uu�7V]aR1����~}A�5UcO[Y����[�6��*&�u�͓T�
&x#ie�`:���l��z�k�A�Sf��✐�ZjP����v�P�jk
�h��bH�����+X�,����J�tľ�w~��YhK|c�8p�u
.�׼�G��A>`�| ���IBvf�H|M�p@7CY�$��tv[�3��pgQ��۞�n��S�r������Z�x&TMMM�����־���4��8��>�n}q}���ݖ��R�0o:H$���7nXPɤ�@�QUX�$n]^<�c?	� =(g���j��-яRX�V��zJ����6L�>�AR���0���jj��l�p�����]���Zڶ���@�h.��&>���)�W�kl_�\c��
Y�ث��wx�h��;G�w��6	x;������B�Z��T�-"��{����+b�i�(K}�M~�l>�󐹾8�*��������n��6��H����';��k�헣s���{s��=�C����
�_��(!ad��;��W��<Ez��-�[� S2Ay�a��Z��Cvg���F1�� �̮�E�7 �K&XM�&(f6�f���;�0ac��H���C:QRc��6#3� ;88����W1G�ѓ*����f�/lN���Yo +lA#��#r��᠞�J!���/��v���w��������G_�YXT��l�lPQ�"�v���Qr������0����QI'1�gE���"w?�c�F� �W��3 1˽9V`��?=����t�y�@g���������9^R��7��
gڧ��Վ�����G
p��ɉ0fg}/*j����Մ��������Y�=j�G����!�`bvDc��$���K��e��\�θ��l ڥCS�����'Qv�у�Mͭ��LLJ��9:J�@;��.�6��Ɲ��R�3��<V� u��-��õ����3���"X ��+)�i����4�_�*Zb��}�;r�}̡��t�����J�Jtƍ`���x�?D��|Vj�_�r��"�e� K��x��s��k8��P�N�ɨHE�GD
  F�@�ON^_�\	�ë�hS�:v�b�{{G�+
��PzRtD&'�.q�r8ȟ�^�÷j��f�"�DcbĤ�]ex�q�k��}f�h�:hK�oB��3[�@�gt���fe-5��d��70���O�*�<.���)KA��I���f�x�liU�� �,�������322dG����6�3�qO[f�c7=&��M7�5�,�.��Dt'u����8�Yy4N�+��>ފw�h?��Ksd�����g5�蓦���C�3�Ԝ+[@�wh�B�Fpvv6�Ӷ	�M�����_���� w��חX���-F��^x��}��ıUr�-��[2��X`P�'�+k{�����Z�	u�jǇ���T���嬢�jr�މ����G�����}�9�($�	����5\�S�b���^h�.,t�y%o̤cL�ы(힙�f�ݒ{��ξ�`D�b�`%�D7��]&#�,�=j�D$%%K<�2�ω��'- �ED������V��u�P�t9��sD��Z�cxzt���{��A��j��=d���*lEF�H��$M׽PGt�Vz�!;D@ 1/�tyzz&�a�:t�*{�5ed"��U�ke��(��0/�|�%̙�b��T/$l�pIӀ%�Ҝ|*0yD�0�p�-���W��J���@gk�ì?�3��ݻwU�����w���L| �����w�'''bw,��?��7w�����*̱r=J�f�n���&����u��������,/=�h7m/����w���(��pu>n=I��ۙ���#`b��0�}ʟv��+��ߤ��U\�I��ё��dy���d��@=&GS+❫ �]�2�3��c���eh=_JYc�c�R[N���JKr��=��i[l8�"�1W���V�b����f,�lq�#�Pw]���>A)�o�ӣ��q����A\w1����A9���L�P�M�Ԣ��N��v��>J^�Ttx�gg�l�]��Ӻ]aa�^PP ��.I9*��j�iZ�И"�?���2�All^�R�s� ��Δ �(W�~V_���������A�"��;I��д���~C�Z
���/_0��L�h�<���L�u����=��KL� �V�~]���:,� �1L��,XR�$ 0 j���иFJ�ԅJ�H�����M?��8�hY(띐V� %��PH��W�����u�O,�=]�j��ؘq�[�%JΚ1�1���;�����q� ���*q���g/'R�۟��sf?�aL.����^������a�R(�����6� ��bQf	***�{M�d������WT�<�A���4$����:X�a=8Y�w�k,�ፖ����,��,�����-�����G�8����
���I�m�XU�w�9O�K�����4��]݁�~V��G��K�"����m��_hNU|FIq��su�g*'��0'��|�-0�oc��$H�o�O��A��%��gK���I%C�X;����/�GK�g��@4τ��خb&s�/}n�P�T	"�&O���J���6WeI��]{`�Sn:�T�� �C�4�>}z��e��8]�)a>e1!��,F���T�j·�ے�d�g'S��nN���~!!�-�0�k��[<]~�O����;T*(6;��)��U)3mmiQ�� ���@�fjS��?9<��$0�M���& �a�G _ v&�M�8C���#���w��l��0�!SW��\�,Po-j������DSC���B���Z:�JüP��B�9m��!�����{1��yN��f�u���S�LdV���\�qqJ[�3jNW,�����/�K\vWi�$��5��&f�� �����0�� ��П��g�������&k;�gk�D�D7��l�\�W�s�.��
5U��7e�M�B��ڧ*��z�p}lV��g�Ȭ����%���hf1�(��=¤���lN�⑇��R����'-�!t4�M��<�T�,E�6W��7ܶ��µ͊���l����D�f���Ek!;b2��u���?>��
����,B���?l�������Z��]C�>�S����z�}%�~S��$���5���ꈭ�,�D���b�l��@�������
p
�j5�����G={�fR���Y��|G(a�L@N��>w���G���Fs>�Oّ�����^oK�n<��z�M�61�)k3c�f4&����t�W��6p�>,SEj��6+�]�ʾ̅�e�~Ng��	}!�,J=C,��O`��v(L?�T�2�j�wq���}L׷�IӢ_�؉[j��J�~�>{W�w�M&	�)4>ut�'�Ux3�L(J��Zi�3]@�a�,]4��:$*X��f;�骧�p*��;�ބ���i�NR>�*���Xz������Dʵ���x���fQdnт��r�����Oe(f�"���3�N�<Dֆhd�.-Z$Q&GZR2C��a[g'�F���;'#�i3�6#BB���%K@v6ᅦ#YX �[��+�� k�J���J�붲��2���9��]���,�9��?�������--�LY}��­��hI�u	�S�l"�ELn��8��8L�yu�B�gS(6�j>�E�6���ݝ�#�q�6�8�����,�[Xk�N�(�rq�u���:9m6�ӳ������L�z�A-�Kzz�R'l�������p�&O��U���9[{{�W�|r?�����̙�~9���?�Z }Cq5,%2R�������)u��k18���3�j+p,%80p	<�u����5�'���~�wINHs.� ��nU$����wU��Bmפ�	��>��`�a{ U��A<+��^��&��'G�SPQSq�����S���w�,�������UWqpss*��+��`��������љ������ht8zkǑOI.������^�d�T:]s�`���C�B�f�	��RS�r�ޟ�;U/-."�h�s����
`|�S"֟8�s���y�[�T �P�S��h�Xh��XXX���tV����p��rss;�(P�*R�+��[b;(b�Ȱ+R;<cg%�U,�/4Z{����4���.'���.O���;6��!��)h���,Sȯ���l�����5^�@�c�&1]2j�Iq���KK#����9b�ھhY�'G�:^��L�ny�2#�?)d���};'.Ǯ�v1�AV~M}�prdg��J��V�yf0Ԁ�v�B�٠a�'y����֛����8�Hٷ5$���@��j�(�T( ���oG���n=n��.#��7s��=^2SsSqr�؈(��O'ե����p�\_�b�A>�n�_ٵ�QܢR��0����u���z��Q��d������`��7��P?<��O��^���[�\����q���b �$�lS"n�	��VքQ��p��"�W�3q2|�_���n$�h�^���
@��Q��S�jɊ��	�,��B��']Z��x!9��v�'GF�j9�X�瞠Cj<vTC�__	�~V�p�{�baAt�0_l��/��m(�3s��82�V�1�%x���{�
����<���ƫ	x�{�����P��Gc'�z3]b���)��#��eu����)Ns'r�ƫ����|�'g:;��>�i�e����k�>}���q&^��e��B$��x��ʵ��s:�a)G���%�U���ίG�H�^
���z�V �C����R�Q���X����3!o~a�ʩ�D�f�z<DS�W�L��t��_s����]|�����k��ֆ��/צU5\�S�8L�P��F	�����<<<g7����R���Qx�*a��ˑ2�@��@bUU� 5E��!��c0d-�..J-���K6�K��)i?(vt7��b- �2�|��TT�����r�Ƅ�w��]�T�:���VS�{�ۨ�e:N~pr�M�D�$H��c=õ���9���o�4��z}�<O�4��!Ġ?��8���@�[�R��Q7�璷i�S�����hwn.��d��"a�U���ֱ*�Ѳ�M�r,�e��,=�ޖv��r\rN�j���S�$���_a=7;�n<�3CGG4����4Wkbb�L���(Z��=� z��t<�T��V�խlm��*PB�0���Խ̶711	�M����Çj�6ߨ���#�$�:� ��p���&EM7����p�a,��l�UvO���[;i޷{L�9.�'o=�2�2g��kQ�r�&�E���jq�2h�[���?cڿ���4�ʵw�c(?�VL� ����� �\��"��S�ER��c8Jz���p�&���{Lz����EDD��LU����
��5����ޙ�r���[�0DDK��^�_7�����z%7o�k|ˋ�o�����=�`HfF����KuZWﳊ)������~��渿�������<��ꉌ0�DO��@uJ�/69����bᄡ���j���M0�Y4*^��M�5-$M��L)V��~�I�#��;����W��f*�,�z�76O\�w/�w]ꪝ�5i? j���`l��E�H�Qͬ��c|z*��P��[
<<f�����L�$�&���	�zYj����5�R��D/�V���\�(��W�W�.��R��$�ߢ�*,���U8=7\7��N���܀�E�̎
��حۨ�t�K���������e߆ɲ��)!�F^�?[ĉcR@^Y/u ���Q�:���r3�Fn����_�Fl����#K������-�o�?���zyyq�CBb&�N!�DŻƹ��`�ę&��c�X�;��CUN]��N&�����76W�o�Vn��Fq�z?h��(6���k�b�=:\�4F�lim�t�'I�c�FC�� �Y9�[��7FSA)cu:�0%�Ԋͯw���{cb"�n�P0�T�>w�QP~�ړ��������2h����x��Ȗ\4��#+��B2>�l~q��E���A��(Bq/��p���"����w���c S��� =����"D+�d=��a�}������_P1���
�����^\��\���/0�	�c��݀>��v�锌;[y=�3o�@1��t�twpq���h%�Ii�%w���^8�%�����;U/��]͋%��Ƃ�����s���to���mr�j���Bs�1��eO��J⫹m	�<���A��;�Q�P8	ɝ��N5<ӭ��F>�y�47>��sRj;�ؠ_SH��|vv��_}}�]��F�+-f�5V�>{ۆ#���s�/���&�!��uy�;�揳�o�ߎ$%�?$?L�B���\����H�:73��p��֞��2ә�,{RX��>�؈��܋��rp�b���Zs���º�-ࡩ	=��A�a<�\Y^�/�-��v��'�,�u�5
��o8�Z�K'��5=O+<�}��Qr��j�D����6��$ܐ�����5�;#�mVRe��LjE���%}�vضȟj������W�.��xw.��k%�,�����dyo�&�R� <\8~��<U+y��--m0��*��@���\R��i���?/6��=1���Hق1�{z~H%����Z���4<k�	W�jH�l�?�+ṣ0`OX��׋~F�=S����
s��޹�o�����+���i��0����u#"1�EgC�Hy��ڟ�`Q8�U� Nvdp���YN�
ƛUPQj�\�w�+n��c^Y]�b�6�OBF�9�;��`*`�>���q=(�҇{"F*���~���t�k�4\w���q����?yw���x��#�$f�ďm�tX����#YFC�����b�?[�������l�1-�&}�uJN��4���V��j.�f�=�F�N3��f%y�Y��Sl.f���1�)���t���XK�*���]��R�>_�Z"�-�������=t��7$I[��M.�ϘLI�\<ȥ���P�0I��"xz������0E��_�y������q
��c��X�Zg
����V�?0�}�R�y�J��x��a��6����I�p0��@����	�(C����l��_�ύ���/G>_9C���C���zUn>S�Z��,ś�K��X���mF)?=�96v�Nц�b����I��0��wD�����9�K�m ��+;�!u�@G�.+���=b�+�'L�9��lV+P�U�%��:��1֩�W���%����';Pc�#����_Y[�ck8[ E���|��t����"�v��M��[F�px���pM�c� �9���5G�Dl���,�2{)��������Ub�;��@H܎�G��M����7�AU
��C��\e�j66�Cqz��xo�@ ��"�KJJ� �(P���vz��H*�����+���r�/�&L�"�ĖN�.�I��t������'��.))���H:�b``@$%�8!#/�jm�`x�~|�f�ǭ{KKK@���+O+{�Z��'K�ZԠ��`�4�~�c9(/?*�c�P?��
C��`���F�J���z�ҭ�*0a�d����[�{͝oj��x��Ü�A�{x����Ԋ\v?�L+̧N�S�YC蘱ǵ���>l��|DDt���rb���'�~m0U����6i�99(���|�7�
U��.�_�Y0�����{G��p���N	�5���9ʙФ�����^�5�wZ��|��U�h St�m �z�9�`�'�Zը,�:�(xn��ѣ���%�\F�\6�Y���Ӻt�`b�ہ�����n~���8�>��7;��Ꮔ$�7NoC�/1�6�.�n��k�}��#��ӧǂ��~z��z�@w���<�篗_&X�p�W*���ݨ?h�lWKoH�]������ŋv�AR�yvj��E�?��*\���w�Ǌ0�Ϛ� �K沲�M|�L>����)���������;$6:�95uෟU�1�_�@�9� %�Q�x;��+�����E��g�ϟ���]5��<}�
��SB*#Wl��tmZ�xe(,=<޾;�C냽!�s3Yn���n��(��������2��-�1\"3��t,?|-".��)�£���7�<�Ԣ����Rf,z5���|~���P]�v�:�aٙk�&k�%�IڳW�p��'���J5e�)%�k�����Έ��[�ݦ��u��_���������h�IT�f�%Ԕ���` ��Z�[|e�pa����Y|b�S��O>Y��!�.���P�%N�㤥��q�8>/N)6�x�+���6�K�a���c�J"Ҫ���b'����}\Ӄv�����/~�$$��ݬh�����Ԩ�_rq���)��'J����L�]o~�
I�w$l,RɨkD����y���j3S�s,�7�S.�k>Uq�<�r��Già'2rr8���T�����~���A�}\�O�?��J���7W��I�m���ྃ������751y�4�u�B��V�ԕb�+��R�y�>���5�����'����!��l����\���t�iW��$��&��1�/ݴ-u�{s�� !�q:�[���*��qE���.M,�?�<U#B1�r�	'��Ք��H��5�R-��>$mɔ�%(����?��8X��p�{��%�*��s;x���Qc�n�˩R�qnn��r7NEk����)�V9����so�\PP�؃}Gzl��D�Q��N�Er>�ռZ$3�X<d&�W���=��I�J�H~�s�r<�$#�Ž���߱�����震!���]�U��>��
>ϗH����@	ID�vw{�213�wpە7�kb�֑M-.����(�.[=�*�h�3�����5�����T	�'U�9[2z��`ˑ,,@�i�V�*\\��޷����I�d���ة�Z�������yq�2�sۙ�8�t����>�6gBB����/����э�rdl�o@ :�ӧߋ��V^�	�~����3&����'��h:˰��h�(HKI�����Hwwww7"�)��tJ7��-�zf��q]���s?3kf+(|��z��{�W�����P7��ݯ���E�;���Li��?D�c]%)�:A�im��S�7ev��
Ӳ5�G�kM���&�"=N9�-*JKi�ڽ^����477����;"��i�����3��gӝ���?����x,f�|"�W.o{(,,�@��͐����߫��4���W���d
���P�}L��~l����:��z(I�U&V0}~�111�>���>�ڪ
$^�tmmm
**A F�nO�mB{ӡ��0�e$9���O6��srr���vv�������W�������{��q��_OOOİ�<�b�������'�ڑO��ZZ����� ��\�LMMaaqA;�@A����� ����D˫�c=���SG<��˦��Tt+��<�N.��.��Q3߽����[�^QIK.���`�B�M��`���N������c�N8���wO�oZ
P�-��_��;�~�Xb��d|�R�-y���r���1�	���bR�4[�ZYYU���\K��]S(�ʢ &���"ڼ�����֨QX�3�Җ� ���H�U:�h���y�˺�������L�2\��sf��B=(I����/^�\�3�_�ކ���=761!nkK7<2��v]�YSO����6.!�sA%%)�%%o�h�������I�ml������{����£�H&2��3���qԐ�E���@���~�"jKǳ�������5�ǝ>���l3lKXUJ������P4��0t�Ԡ�$z�d{{{��H!���s����R̳���D���ͫy%5=͋k����G�<o���w�q���n+�ɺΎ�H�'6�r�bU{�z�ls��T!��U*��)&�'�=0w�r0ǌ��Xx��@�@7jlZ�%����/.������k���Ixg�z���v��ta����ђ��#]�6=�<���>������|&�o��Wnn..���;���� @�ݿ������6D�{~_Q1��X���P����GOl���`�k����hj������z�dz��#�C+q��9F���:KI�Y�z���O�O6JUM��w��k��r:� ��M���cbd��C��PU���w�`g�_��u_%5=��d,5����5�ۡ�]��|	�&!q���%$zj��i{pd�n>wƣ�Lչ�3.�x"�����#���1f�����\�^l�^��֥I�ܝ�Tp���w�ɟ�c�ոˍ�Ye�=>��dDV�G���:�U:��� �]��}~'� ��s���]�%�\ٸ?*�v�xwW<�fnZ�'��	��/�r�mt�B�:�F�.�~Enpp?5�Tg�w�䯂*�����I,��b^ܪ���GPP�v&r&~ӏ��Pcum-��.!CW��x���@���ps2��v�y�0�쬝�������GQQ��(<D�XA��5�j���F�y��Q3���EEp�����p�Wŀ� XB޶�*�������EL<t���⠧ǋ������&&���,~�-���̼� X��Z��i����!766l�4F���#<͗�{{/�,ku�m	)8ʧ����iP��86��Wo.|��۟̇WgW��DJ���"�հILr{f<�(ݖA����@:	�<����&�f�H��p�ɢ/EY�v�bߣ��Ʒv���w�B6"q�%��O�S,l��N/�~���J��.�A�$D��t��}C��㳕�SUYٗ'��v�ZKK��몬;Q��>0������uv���C!���^鴢SWW�b	TzptTDI	#!11<��=N��Ŏ�������&<�0�RR�E�91�8þt���z9SSJ�׋���aA�ۮ�[^�;����x ��'�vt�9���h�?Y�5�B�����ҿ��,"&���ny]O��'+/I[Cw3}�,��r�k�[a�ޞ�Ƨ��f����ܘ����/ߛ���m�?Ci���R�z���Qo�^��AMM��j{z&���l�e��Qٷ_W��B�eU�%�ґ�$����wq.�� e��k��nr�ߖj�-j��>�P���\�Ϡ^o��`���y5���$ݰI��!ȱ�N\�|�����c�:�(�jy�uVkv,!�g~��iM���!zA''f�z+��b>-�Z"����f�wj�Z�)��.q�������=x����%�1ZZڸ�̨?,x}� l�)���%��\&g��S�����aWW�|�7���Sf�a!ii$�����PRɦ=��}��F��hq��{�����a����Ѹ��Դ�H��g�	�O�
6@U�� Xx������vvfaU�x�}!A����tڹ��|�x*^#�%�����	��D���h�}�¨nγ�+�wm`Z:�nԢr<��Ry�c��;�<X��0�S	��/��9��_ppr2b�0L��+5(C/��ِ/���_��_u$���U�7&��ʕ�\�|ǮF�i��!|pNr�.��U|Z�J����A��.��t	�����>���Y�J��꒒W���c�����D�2�u8]�9��������j�V&��t�	�5===t�7��&k�,P�WHH=�
�m�!5��G�4�j��t���)���}��A�9w�gI@EQ1@��*�����0����:V�������^��7C����/���#�H~~~Qr��\B�����G(��e���o����VS������j�g[x$1�Rz�M�ŉ�V��hyl@���)k�G魳jtisj��o]l�})�g РD��e�z��C�8s7�ԯ{�VM��#C׀�%�^�l�G���x�~U�Nm� `��)��R�q�q���3�y�D��(f��.b���\c>A�oMȅA�3�l���͇OF>�������������_���nhH���c����7��a��#P�R9쉏���N]��D�I${����>��yg�J�rԪ�P޽{��Œ����q �q'��6�vǧ{��T�]����9�U���\VD88�&�#��ģ��Ǎv˟+�8�?���v��1����|�* �5���<4W8�9����q5�/6��>�U����	8��&�Ǌ�򍕾�ܖ�j+_�ś���$�Y�>�z������ɒ��Np�'t�ab$,jW�GU]�/5~�_텞��Y�0�1ZE�Q���⢼���U~R���G�$�h��&?����8��ǆ�]��=���~�0�+�77� �S��Ie�q� 2֍�pP�y
������x���������� hR���{B��yy	�CTljy�����OK"��� %�@�N��)!AA ��c�I�����Z\�>���O��҂�u���k'Vi���i+L�sxѮ�(Š�nQ��g��e��`�G7ggg�GN�]I))8�����%��+B�XW�H8��y[JJ"�=q���>�}�cA�NQ�E���:�d9�F0 l�H/Ws�ǰ<=�����H�U-A����7�g��̬i.o��|�a�̉M{��0� ���vZD��M��_��*|5����.ү���6"���U:��SQ��k�����n���uJ��t�U9���t9����N�`X7;]�\�ueUP\<ww&�%�˽|^����
w^��&^)�:����P�%�	F����F�����v;&H����h�P �:�~D8z�`����N=�NV�ǳ�9`��� Qh�c��5:��KRٷ����g�������iK��zNn��� ̒1t����ԭ?pG�`B�r�D��η��S<�,-i�����Z��	+��Y��������r0�r||�gV������ZـC#m���C����e��`*��Շ��߯��x���=3K�\<ܧ��#�%��3������<s�}���Dc�Sc�f������* 95���:�#�=�0Ĺk�c��W���v�>n%�����69UȤ��)�[��=rs�Ƃp	-��p�����g`"""zcf~نԿ/T��=p&����
��w�Ĝsױ|�f]"ի�o��F�}���=����tC�:=��4���`bՍ���q&�{�ѐʲ����֖H&n(�aK4�����XZ��[�A��-�M����õ�N�B
�����b����f-?�	����F��4s����^W��/���X\$�頀\��q�'�3h�$��*����`��Į��2&>>���r @ #/yxx�q?M� ��BC���-8��9mմ���>���*/,2�Ǿ�)d�o%tMtj	x��[�����5�T��>���yj��U<�6�9.9����.� ����]Eu�-��jѾs����d����2Z,�W��<�t6�����=�� ��"A�Ļ'uEf�sĈ��mN������S���|��}��ыkk�G���>�����ףcb���W�i7�j�~�z��{4�u����������Āy'+���J����t��cu�U�ojq�$1��3��2#��
�o�����`�!��5�c��]��H4����G�1X�ɿde� !E���̡y�����'�(˭?�t�#���f��eUS�J�xA�4O&={.�q{JJ���)��u��@����G�**A`v�Oue/�����>�_�333��*]�4JvI�c�  5&�E^7��*�_��7���d��{B�:K)�����f�TU�ws���it��klk�����u�i`m9���Қ���GA49�������{�N|�ڠV�8����✷X��$�E��Ȓ�����<�1w���`��(���i��Ś�n���ѿ�\Z�}�岾~>F4��#{��l^t�b�R{�"kc�� "���9J4x�u9q�AKk���������-��D�(i��JI��'a�.ܲss�jhzR���bss�CQ�Q����bw�ͥL^�ܵ��Պl�~yQ��CB��ftjcr[�]�0^�ӌahh]8��bhjJ���l4�c������H������&<�U)����"<P3�׫袨����8�^�U�+++���&�ǩ�PN�b�٬g�!abb@�*2�;33Sc��ܧ�����S����H���D�b�n�x���l�_�cUkM�����֖����2�Ke�\8��n-/&}���4~�1��yd�X����x9J>����x�@2jg8���D�%]�TI���9��67�}}{f�F-(�a���N�,��z�}�r�%l��w���*5����-7&++۷��ọ����aj4���w󨹯&յ���K�r�����x�^ׇx�ļ� VD�;�7o�y@�K�$DA�@A�	�>����q�O��������݉B�XOO�"ٌ��Vw�	 ��c��#M�� !�N�E)xOLCC���R�b7l�0]�j�7���1��<n"����g޷y�r�RU�6�RT�HKM5����U���f8�S/�D�d�'��\q��2:�b�t�}�?�]gc���K��.���¼�x�K:6//�8\diE�4���))_X���6�=5w��a�;�	Fn.�bI�iv��ݾ�d���Zɫ�k��6��f�t#��:�И5���i��U_�g���\p� ����1(9�UU�m�[-��	�����h�x%�H���=�8��Re^9jcc�h=��ŋk�3��f�F�yi��;�.����Y���Ұ��*�p�'�^V0�>g}8N1�F��L�"�cl���M��Q��1N�����7F.��R�g��}��� ��f��5�h4���I��@ʊ8�����y%E �Q���X�d�ے�/���d5�ߚ�t�.?�������qa`g��
W�o�����59?���B��P(�s��c�R
��#l/��K��a�7f���[�TT�DLŽ��XtT�O}��Y�c7�u7���%5l&_��@v$_�&FG'���:L��2�zw��>��rb�����:�v��+4�Íe$�X�����ͨ���� �|���Q��O"Q����
���p������!H\�E�.w����y]~���$$�"�!�r��v�.R�db;�'�[LH%�]�sJ��\�k����h�be*�ԟk1�|lX�lD,f�K���H���8���x�C�)?����6��x��v�����/z�O�m#|������DJ%�O�w|����b���EAe%�LU�q�k�X��	��BB����I,o� ��AB��v��'��1��c�����E�9�=��"��o�!  t��īB݃�E�����-�͙������X4`πh�3t���*�";�,y���.�TW�;.��Oױq�>Ř5:0sa��H}u gaa�F�ͤ2��8�t׷^���������5u޽�������_���QGŦ�������$g�5��ӱ��q���}����?c���(=�O��S����f���r��ϟ?���;0�>-o�׏�[5(8<�M��}Űں�o�:x�u��\T"L��f�$��?��pwi�,O�ʪ��A٧�8�$Q����bbb�����G��rMޑ�	mpծ4SǾ�3.���h�p}Q����a�����aA���n�i÷���nCI�/άK�X����2~�7��6��.�#���f����|$��ĳ���@����hJ�Xjv���%��������щ$���Y�gޜ,��[�� ��\.����m�5�7Y
)͖�[��'���>G��lqf��L�kk���@}�,�v[��f��CR��ܪ��޹TS��� XoT��A7¤�y�C�s��`B�Z��k �m�J��ccck49���+��%$���%�i��Ka���C���l�����kSSS��s>��迫����n��FQ�A���	&G:���T�ٝ�P	���9�Ɋ��> ]�����rZj!�F�jTr��kS���J��W�c~�/�/��R<�py(>&G������G�$
]�FQV��)����Y�KȖ�bO�n����g-���Ə���ɥϟ��-�ìm� �����ˬ�{��|�!��ul<���Ɓ߫e�g9�&Mq <����k\\����11��yq+�%�ؾL�;�	�d��B��C �SBR��Ǐ�D�&���ħ����)H����Kt��s�@W3��ZZZDL�Yc�FI�~�K��J{��Y���|��CTD�X,q��0��*�V8���mə�!y�Ri 6�M����L��I▱!)�o�lt�����]h������$٘�gcJKѷ;����uts	~���<�)�>pDp��+3z��b��5��Oʅ5sb��k9_>Vn[[-;%�9u�()b9�"��c~�S��-�����O�`Ĭ%�Z�z�1{(�R���,�7%�5i����NN����Op�A�F��~���ج�OM�yy3=*���	�����E6S�m�C��8)(�NF�����Y|)r)@A`[��DY	j"�mKg�@��,���9�ۡFI	��������!��٧.�f-a���r��Df����qD���\v�j	QSJsg>Xݣ��H�뤤$����3F�QbΦ"0��M�Ŗ���K��*�CFѠ�]�:�g�󚤝��#J���p�D��#�}c;�W�Y�j
�����L�"�%���ڈ�d����=�ܖ�i�ڕ��#���LLL�21��@���RPS#FT�����dz,`�/�Õ��	������Ȗ��,,��G�B	��΁�����0�}��튩�h���NY2�Y(y�GCԫ���G+<�D���4R�A� žXȘ��b�E�3����q[Gɏ�w�d�_�`o��A#����N>�ߩ���JKnv���E�#������N���=w|;Z�^{D��*�V�ؘl޲x�"�I;u)��c�"�me]�hP4�������|2e 912"������P�q;�TF�a?D0TU{�~��x~~��z0}.�y��"WII����Y�����o��'"2_]F&j>�5pk�,fQ���sƳx ��cr��eƍ����\5I~��J�G���9���qi_�mL����8����v�J-��lI�n@�B�h"9�)���`;bQՔ����p��q��bq
������-���7�q��<��	�&]Ŵ�4/L�5���kim<PO��nƓG�*(*ƗT �ҟ]bԊ5
r����?�)����.��o�	�������}�Z��G�/��m����$�T8�`�7�IDr���� ��ï�ُ���H�߾}
|NF���*t+���ِ�"*h���ۻ���kq���7�5Ř��{r;�֜�,>zh�#X7�+�R$K�x�1֟��l�l[� F���j��f`r4��7U��{ܨ]�m�ZL|�$��I���HF�}�?�n��C��e����Ey|z
���Y���4��H���_1�A-;;�sٛ^l�NӁ��������xk*�s`4��"�4���l�E�4�>�g�Ǥ�⪨��` Y��1-�
;���~C����2S����#NU�lid��#�KɄ��́���J����8i`� xƧ�6眄c��2��;�BZYA��yx8���BU�zH��=7�Y�����Fy�}4��T썦�=�F�����g�~n�&�|����@��<�;�O{���I_JYB����EcXKl ���<W��ΪT���8h��RR#��3��ٹ�şk'���l�&c���:��>� f���"�Ӓ&C:��G33�|��C��̦��GGLf��2Y����ٸ�.ԇ��k;;!���k��*H�ȸq����bHMq���N'*��?O�ӔQ�F�:��ϋu%7IHI	�x����H�m�mo+pJk������X�4,���{�B'��w<ݢI|dHEEmv+��+9�Dp&u�Q�8�y�VZ��	ZPJ��Ba?|Ш4P2Gm�
j����c\�l�f3�z�M�����s�ʾ����T��l4����z��N�e�i��5�8�}s�e޾6 �1-��F�
�n�-6��o59��e̋��c`b:��}Ь}AOO���H�%�hl7������'5��R7^�c;;9�d�;AA��yr�����#ůii�%��Rl�CYғ����=�ϲJ�B�vI.�5A�e؈��Y8S�"�HLxbZp����LVI@L}r��y���v�TH����	��X�,>�)Sf�����~�9x��R��;���L�����J�������v�X"�~�hÞ}۷�_[�O��U��m|}}����YP���!��������
x�a^z`����_��h4P�Z��\�-�����L�#		�8g��#Pd�"#���ss��^Ъ+��8����?�=����/�t�X�qqg42$�L�fA�{��t��Ȧ�_�J�缩2Zb�EG��G�{��H.M���7a����B,��Őa|��@(|4.�HO�?�i��m��Rr!��*�ǳ����L����,�>{�_���_XB��#����~//g92ۏ$�y\�A�o�Q�������(��x��3,66ES'99#'e�kR��������g�K��2h�#��ٙ�f�p�A�-6ؒWWU�������%^wAQ��l�6J�"�����K� ����*�}�f��=�Ӗ6�RGl<�ϙ����
r7�؁@����=[��~$9΅�b��r�q����,:N������k��#kv�d��uQ���^�T���bʙ]��������ZZK9_�5��BytkJ�F��o���]E9~�
1%PS��?[k*=��Ȓ�#��A���]��	ʣ�D�R�0	
!��K��5nGZiI開t���a�Z����'+JՒ������PhBB��Aug����q�vsk�H��A/��vo��IV�V����޸�h����IIX�K͘�u�>"�LR�x��&\5�X�6@�ƛ,�,�����.]2����ϑ�ʴfSG�!� �Su��f��K|haY��dnbj
�)��~�I<(�5�f�B:������y�MLf�W������`�k��w�/�­&S̟�V�V7���]���[Հ]���~�[�FRҕ~��+��"ƻ9h���I��������{��bmcs��t�2.# ��t�����)[����zz1�H8��啕���Oo8����}|}��vsX��S3�}�M�����I0����M91c��QNmyIt;��{�����q9OB龲��t[' �����/��j�Y`l�1��R�n�������r��>;�T�D�uF�˚�ʊK�M9_�����#N���š��X�/qe��$�0oYY��cji�j��[{ffT��FGFz@�3ٯ��=C�g�8����i�OSr����xbm������վ���6)''.H���|r���22� I�6��~�SL���v8O:æUg������񵧧'�h /����v�*����D�@II��h*�Sd��XeW�_`�N����+����dZ�ARd08��ui���[�Ϋ������1��d_��l��g��j
���d,@���),���j�~���r��kq���a<LB��4��}��4�{��x�{�nR�AB�éM�o6oS�.̾���� �9+M�����(-9�t3[�;8(QZ�ՠ���-&&��ir�������Z�byy�@�+p6���~��lxı�:Jr��=!(=�W�������۳�I �T):*/������n}wONb76���g�@�~�^�?T?=3u�Vh��焪 ����+*$..Nu��'���y�]].��?�a9[��u��ga'!�jr��ZZ���W���%LKk��?̌����>2��DG���Ì��+��8�[���L$�p;9yX&������������EU}�D��#�P35�޵�w!��anG(/+˃^!��-)z^���%9oO��_�9Yʤef"300��H6|�=���0�C����Lq�����ϼRZ��!� -Ibaa�]-B�[bQ�]M�W1���Uz��ʵ�0БZ.�iNU���	q�������g ��MRR�A� �EjO�.`fv�k�VWITUQH��5�\]���'榧_�E��CW�D��eϟ�sEM�r�.��ͯ�Į�?'L!���q�
��
����S����<6�s��d���)���JP��R��"�F/��_���Lt�TW�`ԣ.{�@M靵��eE�]����IBq�:-�۬v��/�IKK3Y�~�^hC���`�և�����g%���tFFƸ�+P�˓|�m��M�Ύ�n����ga!�=��8h �^�� T�^	���W��2G�!>\5�E�l�[f4'����HKK�J"���' ��d �H�_<����9�bP^�zex�p 
i�� uUe:�U��7�1����"J$���`<�,)2_lX�N��.�8c�ҙ _RQM��Es˫��vϿ��e���G�_v�Py�l���4�)�@����o� �}�g*�<��{e0�K]����x?�j�J��SP��>z��D���!� �o�I�:��-H_���B��d�⹹�9���N,�I#��P�Ԅ	j�ff�`��z�/.��r��KK�����_)��GF"	���L�� 5���� ��d@t����U�������T�ST��{���L��Y��l�_��Yi��}��$�b�,�=�ɉk	�xoO�!] � �.�h"�,��7>�p$��P}Ъ7�����Ri�W�GK_����Si[ί�ˎ�SUQ���Í ����;Չ}S����<<�ٌ��{�ₓ������p�fJ�C��t�Ep��n�,�ʾO��864�H{�o>�� @1L>��$�h~��O��Eb��j ��7�Ǻ��9Ǘ������︃C@@`nwsuen/���:���쎎��X��� "���ED^ �ON�5`�SUU������k��y��k5�������%����"�T��������!��x0K�߅��͛o߿�����G�V8�`��c� @�c�Yr��D�������Vh�D�1����絃�H�΅^���_�n����������������r��h0��#&tyԦ?v/�R<ގ_���4��*�₏.�BerX���cFuoi��Z�%��hã����fJ]�,�>O�|�B��D���2݉�/a�`�~tb��V�@{,���͊
���]�V��G+>g�*J�.���!w�Ġ-��'9t���^���
���1o�K���w��2a�����^���8|waj�a�9?CC�74>%����7�)0W��_���K8�8����!��4��� Xx#@YRO?D'�GFj� �'�/]��Ǜ@}V`�@��L�*���Egz�[�ML��:iz���8��@K���ekԫ��א%՗�'$&B��C�9��0�����Fph(<����0�<*���k�Ц�� 	�t+�g;*F�t[Mjw��	|���#m�*D�"���|�b���Ԕ3j�ha���LCt80��&�!���.��zsB'S�.
{a��ޜ��N��W��u����l^xZ����rS�-W��}�:�.S����sJni�7ox�3s��W��qyd��3�6��ߩ�G��M�n�I�*�_��9��P`%Y�9
E�O�>���ݑ��J�U��~���������y||���g��i�993�y����Mhg����.�T��?�I^{K�,�\�����A�U�@&9�]�~�����Dhq�M�H������o�@/4���<��6+��~	�\QJ'�E`�^\({ 'p;n�"���j�iR.Yr�E����VV����ox�x\Bm����,��
�*5���U����K��pUk�S��L�a�J%%++kA�	������=Y3D�2�~�����F��,�C��]�'�%�����ppw&�i��)�����:=99��*3R֞o1����  LS��[0b�PP��h�q�>�O�m���9FDFBn��`���<r4�������N��2��&�h��j��P��&�N��4�r�����b�Mg��z�o�nZ�Y���\mmm06[^B+ai,�y�#ɧ��A�n!"!a��������B��Pmv������\5���L����zc|���)H���,Q̢�f�N?Y���xz�������wf+�����X��0�KJ'�Z��������D6��l31����,L�z�T:ٖ֙����go;���,2)L{/p�f��w���@#H
�_�խr�z���*" �q��?v������e���)(^@��`������&J�N��VW�$����R(�O�@��I�	\C����J��د�xx��V}o���*X[G@����İ	�*P�7���R,��ǩ�M��EP�Tq�Hu�1DEE_���9D	��1_c\�7�������H{�ITQ6rə/yi�jk�Ȕ.��Ӄc�	�u@��{|d��0n)��a�GK������Y��u��t>��QP�r�3?C@E�Oe��]������j��>E"�� *1o��"������oλr/��{3;Q`P��L>\�;߆֍eF���Zs�.����0���$%�.|��?�6��C�����#(�������Ry�>r��G�<Y�?��ɀN����gR��JRUS� ������;/��+/.Tht�z[su�4��sv~��E�8f��9�G����3[[�1J:xC[�a��Jjj�ƥ���A����}��T� ��7�q�;�]��}��������M"�������Ƿjr�{BE6��0夆�F7sM6K�s�5�����V�$�9�E��R��������f,�����u�v#*���2�r{{�36��B�럩5	�x��v&��o��8�"dP�+�Eq'���*<�p"7��&GFvv�����u�pp@F��|J����d���41##�����ԡ���@")!����v�~��!��^`#�_ ��ӥ�������G�J����B��/6߇��R��$�
��8�� �Ulpa������S�@��I<�nXx,}���}R,Dk��fU�g�_:�F<��|B?���n 3l��,)y`�h ~��Z�cwB>�$##�xB���Y�BBn��!�ue��p�k���
�p�D�###3�ce�����Iȹ����.0�M��:�?{v��nt�zY.nX��VAa��Cgo�l����Ң"8�l�.��ץ.��@��� ��i�����N6�X?mk� )�I陚� `��p�i觥�Elu?��ǜ�ֽ~�62��񂙙٤5v�g�R�k���3`����LM�c��TUg���^�2(|��}F��\YU����V�9���w���o;S��Q҅���O��8�ppX��k�m���r���\P��9�؝�bרc7s��,�(+��i)f�I�1mWYZ�I��^�􎷎�C�E�G|�=-�k"�h��Rmb��Y�*vi6V�Ԕ��r60rNڡt�T���S�g#�-�v��z��ȯ��Kg��F�"����]�+�|�I�:���gY`��*4H�wP��E<o�@���P�y �n�[pk+�X,1
<<<���9��
<H�a�*Ն� �*���<�R��wE�`�}2rrt��?�Y���Gr� bM}��`��c�ڽhڲ�8�f��$7��猆�Ap�n���J�^CQsvI	5��aDs-�H���CZ��(��lu��}\c�Vnꪪ�����qD�Zo���q��AGG�����;g�����N/۝%��YXl.%e+)S���]Ix\�XIYy�=���Sk���F�؜z��-t��`��(US33���| �֏�c���i(Pa��E���V���1�	�c"�oz|A'^"H<��LtZ�Ç����I� $��SG�ƀ�1��T��GXYYada���	��ԗ@�E�R�R���d�ǀ�3���><`Rr��UW�v����W�b���F��[ld�jHjcHKû�:P?9���lrڎ�+�vM�&�R��%&$glx��PK����ef&��2�������5�Fz͟gi��e�n)�_�:�F�h���%��������P�%mR�a�c"��������[��Wt�
Htw*�1��⦦&j��"��o��r�x�� aSY-12�48rb�D��A^�e�����q?���145>�x@e1���� 2�����v8���T��zU/@D���Ĥ�d!
������TT$��'9u,�8��`3þ�+���g�(Rx������La[!�G�d���T�GJkJ�z�����UD^zAQ���(�ۃK)���tMf��䞈�U�o��`u$�����{{�&��'��&ǩ&ME��Ce􊆦�����������mm��]a����4����]��8�'c���C���7T��_�aK�� ���I�������G�a���z U��!��ֳ]%��[�ۭ�)���XW5��2��#�-��;9�.v94��A ���+�[�.���iH	kll�Epגɣ�W<�ܐ5�s�x�RG�Q�rU�Q�S�o�3��^��G�eU1 Suus+e)ۀl���!�춸sK��}�g*+��0,¯ ��W����X�F���X;�WRRs�$�g�Uee�����m�ȧ���ʤ�����Сq��$�v����.`m2y�Q���������{����B�j66l�9����"�!h$1j�ZCL�!�??���|�/?Bo^mC%������������� �[	�1�-111W�IIA������y�e5�ll�>Is=�f�Y!�33d�33r5D�3�m��B����nB��UU}N�5��L��� ׽\�\����PH������g�=��pk\�0a,�<ӄr��|,��8�rS���ÖЕ���6����0����v�!jG��ft��Ly�lR� ��|����yA�f ݒU�UO�eѳyf`c����3�Ʌ	e�h��0P���q�g���� !d444�	%c����JiB��U�qRaI�@/GǏ::=c���3��CLdC�\��D���W�����(���9��J:pgy+�tQ.�EEdn�y�[�$�>�A������˫�j� JI��n~a�m����5-�QAs��4�Z)�R�ZE�Sh�t����z�9߀,�'&j�Z�L}�{��h�$��Ʌ򮰼�,.!�9Rx�*tn14�%�&=
$@u�MQ{{{] �a>�������������11����VV�����Ô��_�|�z �~��	z�"mLJ��Y�[�&(QR�URRZr�d]B��x��0
�83 ,��G��U��G,��SGXɤ�x%$$���9��%&�S�i��|��-5%H$>,�I��*��5	�D	m$��,�-���:�L�M"�R4rKKGVJ��1p#�u����$V]����X� h��`�kl%�HHa�:\��g.,!t����z�����D6�.�tr**8じ>���r�%�S�E���y5����[�#G��B�p���T��FF�;�+ܺ�N/�\�Đҽ��+��aeN��/�4!������I���5��⒦�Y�|�ꊺG�E&���]/��g�f���g_�dXs�G��m0�J�H;L�5c�#��w��jtCy�ht�������VD�h�П?���0887������z*�+-��
��ԆxjIH�<<,%�ŭ�1���2w�*4:ӥ������s���1@��?~�8]{�OAO/��z��U���Rxf&a^M��U�3kBiY���N�@c�C 7�_km���ɛ�:�'�	s����M()�!>:���~ME��*4�w�0o��%4���[=>�M!��y��$����������VNh�%ِ�~jOH��Z��X��V�"spp\-�wa�����Ax���Ǐ=���n���C�H?`�b�88��O`�ƞр.�y���S������������Z��xll�u�	Вp<3V�~ z�����g�>�{�0��f4Ǯ�f%0]#TU����9���ݷz���Z~O[X�^,ļ��l&&ǆ��w���{��9��D�S���@�ftb����\?)� ��g�9�Y�%�+II��333�U�<.���օ67s�������e���?�FFD��W����#��Ņv}��3{a�Dh�,(�H
�����c^Pk�3k�\jJ
���DX�͐r.ڞ��{J��3��hh�-*
955u��a���LBV����������*��o�D@��S@DZ����/H�J)�HK]@���D�[�|����{�T_��=;�3s\A�-�������	Y�2��7����i�u�m&˥S����@p0���i��i��.�b���}|پ�7�S��碀�//g��l�A��t�Uq%qqq-?���_�Ť�I�ʚ���N:��.���,���ꈜy��sZ�p`��(����	��������
%�G# ¬��Z�>}V:FjQ2WTSRz{|+��:�B���.�S���Յ161��B�fC�r�\��3iaeiVZ�`���d5)���]���K����ww�߿��9�\��9M��@�+|O8�U�S�c�D���3P>�3~e�B�h𠀑&މ�ݏ�כ��ԯ��V���¤�8t�w��\�>wY���9��A�$��҉II��+�ӰT�9�F,�5����P{�نP|l��yjƑ<��f�bj%����ϟ���!ԲR����v3Uy���;Y�����ڴ���zi_��p�^s������Ops�|���C������h��uK�n�z�?�x>Q�G���T�N��|��Jk��9'�22� ���Șd�dݣ0��ل�x�W�&�P�\�4N�P���EڔT��~Qņ-ͣ�|�$����lK�4���zT��KN8ͻ(F �,P�ޙ{��lRMO�v�&����������)�_�����5ߢ^�T=A�m�\4��ǃnob4�ay�c�(1ѣ*,s�\L�n�O�۽�΍����U���䊔4�)
-C;�c�P�������9lE��F���QYf��u}�t�N,�?&\�K��^�fG �T�	�[x�Si�������ꦘ�:�B�z���=ŕ��Ieԉ��m�CS��n�°�u�8S�@,]�+<]�$o�=�")"eq__?���P�{���
m�G�{��B���zZ����+kiYU�������}#�RN�0mt��W���%��R�޲nD���) I*���K��״q�[QB����p_�MW�)|3��K
ͫ˓O͒���XK�<�slQ>^^��;y�C���C09��
���Y���/T+Hc&U(_�����*Yz��D�@8���������
e,�Q�]�3Z�/W$�ċ$���dM��j6SA��"[YֻR����sO�莘<��@� �+a��N��5
S��]�&a�궍�dEYVnn��x���	.h�40����W���/��Yi=V��Do�l����ڂ�>�Id��TX��v���
�f�4C�Րݚ����?�����`���V;��7�I�m�y}�=�̱L�����_�����'z?��Sx�3���d���v8C]CA�hK�)�BY�=���7�: n2�^�k+c��B����zaTF��:"���=�Z�A���L�7�߬���[�O��,�f�P&��4��ӕ�M~.ؘ=z3�[�qq��o,O�> ����8�yn��J4]&�'���j������L0�
?���30��E؂�;����A����+���l���v��22h�''%XOʡ�)��&�s����5��*�!"�C��i���'��fo���N@sJ� �ǌv-�f���Lb"(�҉�KR�A����pT꾫%�L�y	��L�ŀ!`PI��y����[D�K��ٹv�]���x.�h��bk�r2�u,U�:2����x���a�L)yy�	XI[�y�=>���m*[.C����\�:����O�>���!�2(���3���s,��vo��а����#K�?��./����g�l̍f�c�{\y0n�ȱ�W��	�<]5��%�8 �5���`."�eE_���N̏_2%!���crL�D YR�99z�m��ʯ{��DB�O:���Z�llү��n���B �f�l4� �9�rs5K%0�y���!�N����
^6�)(M�I.ɽ��-�.?�2{_��X�]3U9ڄ��~ ����|��yҎ)�����G.�����r��|FQѣ����5���h�P5x?^�4�^��S,w�������*�;0�x ���lmRb"l�*��tK/
g�!�+>>Q�2��2<T�����My0���U/Jg�}1��ӓG�/A����,=@@uu���T4+7z]�E��ˋ��.v�Oζ'pH�� �-!L�9�c�	��*��Noΐ�}(����V�֌/O���[2~��#�~C04�ư�.yD�
����Gc��������Jrrr�8��������կ�7���-��Ɍ������D�̪���=y���=N���<aLL^�\�)���� ) 3�/\��U�P��!9��X����������R�(.�,�D�X�P�eOȬ�����,[7����j�@ߛi��〗{�w��n�.��Yw8�j��Lnl���5��瞦��t Mv�e��3owZ�2^�D\��]��9��T����T�N/zBS��Qz,3|���i�J��LPӋ3�?kI!�w��l��̕Nj���2w�@DB?��^붧�`�e�h|��5�Ӓ60A�Y	���$���/���@mK��;S;4�X�is+��'���O�d5����� �h�@��� nj]\]i�jh�^nf3��s���B���[�:����P����������Y�Ε��-��BC����e���D�
'��E�'�E*5�^��#I�O��3��� �dj`n����+�c&Um�����3ZK�P�e����;�����Rbgq�����:�6hK�j�'k�w�{)�������u�A��rQis�x �aY���ɹ0Mp��m�����qo���!���W���3�c���pֶ���Gۊ����9���uk�!�ů0h��2��L�1ڷ������8� ?�&���B�FP4��2t���g�鿅�q̬���������0ٓ���鍻�ل�H�q;ڝX��*qTʎE�|$� a�����QizI��:2F��^M��DOR�9	�O�,^ZT�GU�L�=�g���F�`1��#ps�\��EX�����@���� ��K��,U{˾z���X�b�Y,�;lc�����?�@� �bay���ek2��mll���s��LzciOO��A ��B�����CLR2��ׯ27�24&���[�4P�0T�s�aii	��Q���'����OW����>GA3&������M��<D"(�d������ti�"Z[oF�k�@� 7 �
/T�;��a�ʩ&������R��Ŏ��eD��C#�����!p������-~M�սݝ������7�;�{���3��,āT�VQ�$��o�4��\y���)hi�FFF��x��i>����u.u����T���<�&�2�#��-S��#U
�@��{�A�'���Z�N�6��;f&�󩧿�������R �M ��8K�w���k�°:�b.;;f�����k5�#� W)�� ���.�}�r�sN	Q p"ܱ?�L=KR�w=��,j�r=$C��&� �@�rcQN���w��|5Z�-K�,�c6_aE�����c���ʪU3OИёus{y{���'�movy�{����\���U�~>�U���+B,��$��tA��C$И��ӂ�շuz�N���� A�~w�.,ʲPQ�:����9��dIXoԼ���
..���zz��d�P`����k�QP �_�H�}�ss�jt
�@��8O�N��y?}�1��YW
miNOkutu�G@{�|��Q1ii�U			�-`
��G���N..�[��	ѡ�CCi|��o�x�o���tפ����s�ǀW�Mv��c�z�&бNoS閺�$I������P
=��c �z"B5ŘƲ��23��p4���h�i�`+��m���rl�A08ߑ@��r�aơ�����ˬW�%���n}m�L�K���\���}$ !(6 ��/�y�˂�DIO/����� �mtL�q�f�d��w'..�.P��d�Y��m器���(��RL�k,�+-�W��cAU�)\��;�]Fύ��^:X�\�顺3ҁP��ֽl�p�@W�5I�¶I`�ˎuy��(3mfB[`�JO��r�hE:�Ty<R��6hDs��H5F�V�}i��H�48))��(08:�X]ׄ��Ŧ�S���>	��A���\�$���\�Fv ��5552C�VCa��М��¥S+�7W��3h�(X)
" �m}�����?������H�g�gdi񻉎����Uy|}�q'4Q����t��3oF�dT�����q �1 ��dȑ�{�y���7��HFX.�4���xydJ�CKּ�j+h7���.Glo�*��3J;يtaa���JY�T5�=<~����vr*K����N�=�ij�U���b8ݾZ+=O��p=�1K4�*�n�9P�E�)�����Q�O@@ ���0�Ey�7Q��K-�L�okjj6���^{��������iz�e;�E!�7��`<�����������:BS~��܇6Cy��a������t�)�VQ��\a��k�S'��h��U$�2�db��ޑL�򴎑i�'s"i�'�{y�BC���1�$ʾB���ޜ��h�w�+��������%���B�utl�3 �9���8r�*��
R�=�Y�/ÌB TE���Ⱥ��](�]ڙ۞�7;��S��UJԁX&��p�\�㦷�T�:4���g�T��CW�s����C��;�_��p����kX\��K2��)4��*�P��&&:**R�"pc��w�u����Q�$��pCS�a�V�ommA}�����`�@6^�C�} ��CD����:::��ٙ� 2I<�d��!Ї�?�����}B9<q��"M��k���ԑ!�2�<L��a�_vpAu*9ϭ��{������.���WW�+�o❛�����t�NO"'�V�����~,����?!&�Y�pk{�92_Qc7c�nŘ�Rp8c�a�;]��to�����
	����oT�A���0\��f��3EC��)�x�N�/���2r�̀��f	qX�����d�jL�vޝfϫV���zcr��X�
��q�R���������oX�a�4�m���|��Ó�4O���y��"S������M�$��"jl���ghhdd����|�(��^���U����䊟�����L��E�$� ��ڢ�� x+Zo�tM��Y�Ѻ��effzl��;��@�[�e�KɁݩl%�h�I�����Euw�!���>�	�)hf������öG�l�B�ch�VU6�#���W��z?����w����R�`ڄr/�7Z�.����
�󃥍��Ky�h�6`'�[7���"������F��?��&�Ѯ-6y�����#� ���ʃ��9�VX�Ca ������9��VO/��9�����w�.����-~hhhq}ۢ�9�5��j�ݛ_X8�e���=�r�~|F|���s�
}�TH��sA1�N�'��y����}��T� D�5�f�	1u� �:�F��
@��n(q��?ʌE_wz>�ߛ�q��}޳5�D3}u~�xj0��_�3]�QҖ�i�h�=a�?��Tj(�m��� �Z�2�Ŷ[���j��|�$&��d�WYW��d��6��\RdJf��K�ޜ�������O|cT`g�����7��רE|�Ga{O��i&LM��7��c~���l^i3H�����cά
����ZB�2ct�]�b`1&��JJJX�Ak�I�u1�$�S���h��v9�ަ���,4��v}����~�N&WDJ
� ï���'&������|A8�_��ad5lf.H��L@�>����L��+a����{Dd (�Qwr�Jϟc3!beE���W�<����Y������%����������Z1���#��/@�)�O��f�Ī�!"�����h~~>�V0V.�L�dT��
�8S����=N���m�?�
&0l��4O�A:�Q�Ҫ���g�����qF�g��r�o��9a1�0���(e�#�h��'�ߜw
j&��ރ�H�b��O��A�g�x.?/P��
 q���K5c/HC)Y�l��@���c�� �5b��'��<>;�Jq��7���(삶���7	�;`BB:��:p����w�Fo�M���0E��u0�%�D7	Q�׾jL<!m��n��d��b��pM�+��5A����O��Dށ��|����U������w�AS.�á8O�>���q�������{X��> �h���V��r:K�2PKT[�(�:��ˋB�¯��H�	�l�k����/�P���c��m�y�{�-*�A�����Y]_��8@k}	2s�I"�#"��]�

Uw�--������3��������N���k�S����\�*��R� &Y8P��ll�@?��V1y�ޅ*(Q�2��7�,09d�mi�S��%����>{�p�IZ"�6�ᘄW�񪹢G�'�*��v&`��c��=A8,���Y�4�r$��1�O�HW��:^��wX��~Y����ժ��/7�LÔ3}n�%;�'��R={,{Y����?@�-��Ӿ@�{S"̝�ud�u���ܓ������9y���.h߿i��ե����Z��;�=z��Ԧ;�k����{�=�S1�N�:o���ߨ;�zn��&�"Cu)��Z:t�P�ݰhB�9����4m?��߲�0L0L���p�3�f�����͐���Q�˻�LMª��x��	��!�\mŪ� ��h��� ,Sts�&̜��!�wB*򉊞X:����2Us���3~R�����|4��'���~^�9c'F�M�5)�U͗���McC��4�A߫�w�%�4��HлѲ�ޗޤDG���� �t<�O,>�N�A1݁�u(�|��*,�,�(j�B��[[1��zM��j������;1?���x��^P�&7�6X�n('e���g��vAOo�T���v�B�X�!��G�Ő�\K�
��#;qw6�����`a������0"���YS���w#;]�-�
�bе��=qp-٤��I�y��IG7�߈@9�F��⌰c��g�ZB����xt5=2�����fK l��n>Z��r�͠~]�v�w����E@@G��.W��ݬk�����h�K����׉�(�8x�p���+z ���ޤ�+��I�Y�4,X�E��i��������d�!/��n�`�ㇿ�9r��0��W�E�]�7VX�CCecR5�*���2�hV1K�A�vc�v@Ȏ-7/�ɚ�𑕮 B��Kb����*1��fŲowl��ܛy2�/�9�貇�'�Dxc��$�jf:�������4K��&(w�G��ݻ��.���x�]��n;���֩3�\�>�y���Cb�p����8,�(����6��_��Z��xFGR�F&�9���	A�ܘ�B��S! ZO��hx���� t�������;�ot������:tq{}�؄�� 5�\�X����ץSO�SwFl��7�mYEp��#�����|3��y�܈j���&�Z��4��Nw`m�30g�딈i>���5YU**+KJv�b�`���\��D\��焌�M�`Iվ���8gs����)I,*�C�ٟ�s�r�'��*�����K)q�o.�;�R^������ǅ�1[�ip��g�wZ'+�iە�!|� ���g[�u0E�Z�Ҕ�
�ٷ����2�t'!�utM!]�e2��=>)CC���+��%.�<e����w5n�@7�t�)�����N	T�,(Z�3�~��Cg�ɫ���$0�4����f�o���"�^�ð�X{�C��%Hĸr!"u�9ampJ��;���t/|7��3'�>i����e����jmS�`c�䩳:�jM�ga�#6�t\2pE�����Y�|�Vn��e#�m"E\/���7�d�)�z/�3��o}���f�������E���K����u�H���@���gg��{����!9�4Kos���Z������������N�Y
T.b�?}�2WK�Qm���a�/(s��!%?�U�Y��b�QΜ������@͞)I�;E 2G�v��9�/X����T��,[�*�h�~���mc{.���⢩}'�%��K��\��l� �77W�^��>�������@T���]�����+}��T�R��`�|��C |n�E1VM������)b^�\>�����R�?�ZPF�����U���̀�b���H7�E��U��c�Ht�=8�~qgo���|��4��4}��1�T5&r-]�x��Z��)��YC��b�� �0�)�v3��v��A(`�����i@�O)��o$��S�TW��x�K'�A�H��@�H�JJ�0�Yϗ�4�?�Bϳ�������zM3�J�g*����K��d������&�ߗ���Tv��_EKN~N	�u�	9�T�JJ.�~bߙZ5�~w$���x���D�I	7A�g�ܾ����	q���Q;��a�B�ݕ+�Lx5P
�JX���QdkۖrQd�0}�o���w����R�#u��cq)�#n�t�ze�`( �&�؏�� �U��YJ�7���~o2ߔdY�VS�}��52ب�bp?XI�N���~�O�v��$��0�-;p����%�ܪы_��W	�]8��5T@x��m��{g�m�9.	"|��W��.���˵���Pi=\�@��.i���"d��蓋4��l�|�a0þY�:2�X�Z`��ʢ��l�X������=w������.n\�u�Ȧ;թ��>ܰeh��CYYYM��`��C���iljZ>8`�?ԧ���s�?$��K�1�v���at�	�@��!`��Ѻt�N�K4��&�����-�m���� ��Wԇ�IqW��Kb����\�i`m�KBd59�g�-�)r�犛	k�3ԭ�������]<4�l��z)I�,9��V�וW`�0����2c^?���m�է�|HH� ��m��qV��Q��H[g�C�_������YV���}�ci��@�l���Q@�T��(�h8T�;9='�� Z��p�2�`
�՛�^�$��M���%��x��X)�p��H(�{2��1ni�xM4<���x�T|=���)�Ϲ9��Z�L[񱱱A;�z�R��э�Q�d����8�L���� �FO,\XS~��@�F<�ZDD��_���a�UG�Q+).�<EX��w���2�� %\"�~�?!�zА���ɳ2��rio{F���I��h�pԸ��m�JO���	�M�<����Zh�]�c&3'�z��g������b<_�8$�`1����V�׿�1��2�+��m��\I)(�o�1ҩ�3kW�;�����
�g����r:��3���oͦ���ҙ��33���e���`swR����s��2w�)���ٶ��ҵkk�q�|���
�kb�����4�bK���]�Z~瓯�� O��P]���B�-�B�:,�K��dz��[4�5���)������g������4����������Í!�u�+Uʾ'IFEfa^t�tE���1���;9s:K9U�HF��g
"/�/�a/��=#�o��my��#}���]���pг����K�����+��u�Z����ߜ�aY�m�w��c��=ƑP뺅��~�T��o����T�>����Eg�N��F\~)�5p��*�:(��m+���Ө5�~���#e�i;x�ˮz�Q�?9%D�斌�_j�v��~���J��]
D]�ٙz���ii�$$ϰd�1�yB\�'��ֆ�櫁�����ښ�Y&I��]��@*?'y����b;g���Cd�t���־
7��'xk���3?|�Z�_G+P���Ҕ�wD��ͬ�꺴eX�32�����,��ߊ��7��9��M��5+�i$yՈ���+}	LR����}����$����XY���?��iE��FIL%���%˫�8��(|\����q��6		��m��z���Wn���v�׋�I��`�G�{�G0������]�ϼoB�Js���v�ck����m[{{D5'!��N�'�ú
��U��0� ���W����:��Ņ����(�8���崵�c��V���O��i�dm�k��(�vg���@zu\��.�rY�w�x�4��^�[˛�{�@j�%Ʊ/�����OB#$J�g���Ẹ�вѪ��JM-�U����. ��_�v��!!z�$Onܑ�|d�h���k��K����k��]�?�?`n��=+kF��ZY]�A{
�L�A���6U����ni��t��@�x_/�\mww�˰L�`�|ɘU����3���'�/}e���=�m�/��%���[Ѩ>R]3� ��ή��*������)ѭy	޳��3;��(�}jZZ�Jw�.%�E���`�������R\H��;�$Gߒ	���5O�%� �^q����}�-6�v�t����o�U�3(���"�;����v�D�Tj �W�y��}4^&w�{nM��jv�yZ��1�ۀ���n��Zj}�����e-��f�;�U���\��6�{{�8;}�A�u�;��m������:�or�qKU�5�/�D0�ܽ�(-6�6ʵsUd`k���r{TTT��.���W�����R��A?`��}�-�"ID�� g���L�~�g��ʴ���s��� rB���8�0��.N�!���x�7㱯=��V��	Eš��#ST}���|�������� 9v���j�J>�KN�go�B�mr7�qݿ?2��,���~8��[����53���r1x7	u��R�q�H}��j[��Z���2�?��ہ�n���CY��Վ��V��_�V����%}���VeL��7N�Յ��@�ގ��D݋& ���Lu�����������-�vX��ņ7�?��嘅7ꅙ����P�cb^�~u,�������U�a��Tt�����8T ַ�`n�M������u�����j.:�n�xWP�VC|�mTR���\�����!!�G���Ixa��w�7��p�j���6x3��_J��.�.�VQu��Ì�1�(��<H���������}|�5�R�l9�/fx$ڢ�:�+d^���t�ޒ�������H��}k���O�)6vtڠƳ�Y���rs6���<��R�����k~l�'�����AV�M](��?�Rv%�����r��|,[�6�;ɡRV���؆���1�R����GCC�Z5��ę�Q�ޱ@��ne�$�:Y�(�8���+	�f*�{��Ԣ�"�4@�J�|͒W���)�li��a�d�#��%�+'
�O��A�����0���� W0=ڃ���:����Xg�ݬ"�UਤN��RR(�n{}\��O��l�����\u	X�0����r��������8�̲��5I�v��_f��^�32�ڞ��T�Zh���W}P�|y������M�{�\�9�{-K�h�y��a�SФY�b.�#Ve�����I��4�_����JuJ��:6�����(�m������><v�����˜�������.�����������H"N$�����*���I%������h�v6�ae���d��t�P��>��댨!���������\�e�,��+�`o�bʉn��ԫɟ{[�_�M ���mIj�n�a�;���Q�@�^2��^U�cT��>1EL}c�b3���l�n���ul�����������]ᛂ
 :��'N���ɋw+'/����󇈈5��r����1��)7)�T�����ϻ��0�n..<�{5�_��	�8i�p�>�$�7znt��l߹8ӯ�'����?=/�	m� k�������Ű��h��=]\�s��}g�v:i�y����`g��_����"��*i�-w�qQ�0'?ϔ�)��
{:W�m&�|�Zޗ/��X9�|����HH����Ho|��,��7�%��t����c�+��"�:�������7XM�-�o\M7�7�-C�о���G ��W	�v���d��/� 
�=�w7a�����ڣ��m���93�� sP���W�阘����i�Ƹ�556��]s��m��sV�����N+�����Z�?�b0%��Q�}�h[�ݻ%.. �`�	96s�0�����|X�	He��)�s�D�`����yxx>��h^��Q��5��Y8����k2pe<?_�*����G�6\����x0y���^�2�k����ʞ��Ą�(O��Gzc&���
�ĉ"M���6�׿P��/��3-?���TX~�ݟwQ-��G��G�������Q&6~(e�]I��n9��� ��9"{�:\ޜ M��)e�*.�u�|�\w��gh$%���H���NtYn:�v�]�ڮ�q����O�;�[�_Q�(<��܊oD��(��q<vc'Ӹ���1���w�n��1�l+�Z1��ٍ��(՜ȇ��+�<k����v�gm���֝��'j�u��U�Cg��Y:�`m�l-v��2�nn/���`k4����	~?0`N����+a�Q��
����E��.�����3�cA�W��K���;��}*G�`��5
����<�Ho�O�^�<P���k�Iu�:q�8��{5K�sR��.7�-J:}�(�ⴈ�܅g��,�?FIu_(7Ip��G�������9�m���X�qL�/�v/�P��������'��`��H�x�� )>�bO,�R�T���:J��џ��<߰���Ǘ{�s�7��p�Qq���ڶ}%[��1���$���5Z����.vWk��zEX�r�{���s��^�q�q���ա���yϫX;oF�drE���\��*7]��c5p8x��?~ߢ��y�u�� �����j�� FG^j��0j�1�u{�ww
�ٿq�f;� �^���T�.�(2}{����SN�t�/��bc�&k��z�)��Ŗڮr� �H���;b�o�� u�h#B�(�T��>6�N3a]xa?��#�*�t^� �b��z��nux�]�t�σa�m����҃���Zϊ�{��F}�d����>R���C��Ρ���l�-��:o�{s6e�Hҿk���KI	çddD� <gLL%o��~�ӽ��r��ؤ����55`U�|N��MOk�W�gV���^��Q<*�9��߄��D:�_f**I��|de��5���
��粝�Dũ�֩we���ͨxhG���=G����u _� )~9����Kr6�|���<�+�ZK����En�xN����-a�f˾N�z�������q� Ռj.���}���l�����~�H*�u�=K<��cui�2߾q�dj�����7�P6$U��}�q�UՍ��'�1�/�G""����ī��%��Wg�\7g�\���+3s���	밀i�+>>�U==�Q;ۊ��+�����u9�xa�����n(�q8.m���\�,��,�͊�{�)���8uw/���Z�Z�1��j�������k�ၾi_i戆`X��Ѥ	x�C��=}՛��H��GMCc|����f�{���=�¸������Es���LYڤ����/�����8�ya�D��/�	�$���Y�7󟇦�O�_��Ü{<�߽{_�ki�v�ة��M�o�a�*C�jJ/*��~���W��D����L䵼#y�p��T��<ϻ+L̪�N�[���&�	w��N��_n�+1&�Z� �xi?;N5ŕ/�48T���!�F�k/��Ͳ��f_ 2�zrBq��T|N���,u)�^���2�S5B����v`Li�Imi���1��9S��k�rfx�=�����u��K��(��8��W����ַ�B�i�����窝�Ʌ��m�����;S_y���'Y}�����\�j֍.�������GE�ݬ�.��#��ھ�wXaѹ��Z���]JA�k#�?���ߠ�����H���r{�����/�djq�ǋަ���ٙ*��'��	��ʫV��ey���b3���2��q%/�	OE^G�P��*�qU��LshX��1T�bg^T�FPwf�
Xf�n����s}�=��?�R��iP��=e��Z�t�Ay����r�&��b>Su�Sw�Pܧ��T��V��mA��.�9��TLW�=�9^�z�[1��������!�P�Xb!&j*���F:,���V�H���<.���o���q�~Tjn���w���{�Q>�۴6j~0�{Ӗ�8㩿�����g����{�I���DOg�NQQQ7�p4��&KtW.�V���~�<��n��J�w�n���)�����[�� D��x5��R��>F.;�I�W���޵��]�U\BWO].�/��ffr�v�����whv��\MP������q?�H�,�H�N@�#E�l#�R)2������h-oo����􌛛��ܜ�����r��������Cwww Bpqq� Q��+;:����u&���h��߿�NV�{z��&x��^m7������BC�0��o�B��<o��-k*n��_����WS�-�y_`���;;�i�f��/�]��š�Cs���Lr�p��Y��tF<4��E
����=�͹K��*]'2��ѹ~���Lֵ�/��*����v8\�����/�8,4���Ĳ�S+62��9�z}ɄnNqf+�M�w���?���E��jkW;�F� Ǿ��]i=�E�^,�4�I��r8=�=:�C���N�k�W��?~(e����H�ʊ��Cgÿ���M�*c:h�L�"�����/��^��c��p��P�m__T~�>@����@�"�<��YQ���z{{�?֭���p\$��y��@��o������6���ʹ�D�_�IZ/��5x�;�q7���7[���;��缝Q��[�� ,˹[�)vl�4�T�<-�Ƃ��9D���~�j���m&�#�T���wҘ_>J�,�0� A+�\.�-�E�QdW8���>�6�����S|���w�������a�b��.��oДH昴A��t��JkUJQ00�I�j �S12ʸ��"&.n��#ss�����z�;D#l,_�����V��c�^�I�����B�H��KX���AdVVV�]�MLFF���4D8QOO����M.��+�p,<� ����
Y�j���M��/Φ�]6���fA�g���(3n��H㛢�	�)6��<���# ���I����-H��!�Q���;�J��o�`�Bu�<�o��OK�*�Bh�wc�i�[�^�1�K[���@�?�<�j_0�N�����}�TxoifFAE��s�O��U��*�*��?��,�u{�Fʣ�y˗�!��͚�o�����E�W����_����JT�^���m�Ln[�����vU򄰙rSd�Oi7���z�$�ͩҌM�Z��@o++�<��$����O�99�P�4�$�����H�FI1/m��<&�W�|�|Nu33jZ��@K�k|ttȀP���+x@T^�i9D�P~1"I�\1,X�"�������Y�?�{c�e���u�*��\^ol[�� Qn����
-�P�RC{z�(|��-Ⱦd�aنP�V�
U]KKK�&33Sϔ	a\G];>m@{p����������mkk+���r��P���#1eF�o�A��|��v�1u�u��_��r�I�M�	���s\�m�\�K��d�|�ԵXө��n=�SVQ19�r�%�$�y�(��4�P2tB�Lu���1�ߕ��g�1�;�I���F@�	L����<@:�$�!��a
��%/�=�p��s��'|�D�|����AX���JEY�<P����P_�t�������SN��������xxzj��A۰$FA�-��ON�%��K����Iܿ�9Eх�J� U�5�%p4r���wԊ��}�������!�6�v�x�c��e0k�NV��r2Fu���Gp�@�+f�+(�T�Ԯ���Z~�I�^��KwC��޺�T��`��h8��w��[����Rd��m���ż���7sYX���{�l� ���P�O�$@�r��W<�%) �UT���/ж���~h4�J��>�->|�"E� z&�v
��^�*Y.�����6,��"&43��ݹ��_�ҞA����=`s��%F#��f��E& r��r��X^reZ�F%�.&ov&;�|Qc������}�T��a$�s��Viv�Si����`�niyǱ&���g�{>:
`Z���1.Β e�ht���
|��U�l���D�$���e[�������UK4L���[�����Q�0�оn������\) a��0��4]���K[W���:Rq{2�� �oE���'js�`  c�uDS�:��reۇ��An�Īݚ�O������T�J��0B�	������		utw�+]���9w0S����5gb���A���
y���}�c|dY*�����r�	��4�����OR���~'H]g���&�	��t�/�.kIvN��.��s�U;U���<���~:���&�"����;\��&�44sn�mw��Wn���0v��GIb�����ݝ.� F��l��Q�E���O2E4�R�m������ƌA	'pñ�m��U��OH�X�-LZcY�� c���󤶻��WpBM))		�/���!Y��iiA�FC��)7��2b�!y�
1�@Д�M�D��#�x?b��ܿ��v�о�+}4�j�hl��[�׬�^BO��3�*T C��p�R�d�oOA�
UTT�BDvqK��?���p�T�S���Z؀�5�a��}�"�^�\���<Ȃ�x�o�0��Zo��\$�v�υL����b����B��9AH�l,JSK�J��l�zҨ���MϷ��,QR�R��W��-�x�:Ϊ��O���E/[�9��)�F��;%˺�����P����g����/��f@�g0�7�����F�g�F
ՙ�f*�r�&&T4s4Ԃ�d���� ��BT��C����c�wX�:�<�a���/������!�gtt��^��<
�3)��
>&H��α�3�����#!j�}C����-���/�[A�{|! ֭���Un($o2U�g�m�ͣqK8������Do�>��A ~��E%`�{]�SU[
M����q����@�HW�<C�k����>�@P�V�Nęu�n~!�\)a��wq�m+��Ε�+�I��x?�E��j�ښ�?A�J���gN�ԕ
�G
��x4G�6��[|x8��+����j P�� �iw NB�������YYT��h�!v�PQ<:z`@@@�)��	Xn�A���򭔆>�HUa9�ѹm�A�>�U��7�j�u�W{n����<&))������33D��釧�b@V�T�Y;���&w�Dۭ�g�G��9^��^�D���)Њ���*[�6��!+9?���n����q��~a������n��-�S�hrWb�Hv`ڜ���h�ʰ,��kDA���������iA����n�����o�~���ǁ
�9���k��x��):1!!|Zvuu���	>P�B^�2'sd�����Ex�rs����2�6򞤮�c��7��d�!eg��2�'��b�LҠdz�)�4����1,mz{�↪�T�8Od�{�{}s#���:`maxZuu{��	��E>j���?��"<.g��w�Z$^6�;��&R��G<_��\�2j�<��e4Uz⹴L%����E
������(���E�����x���o
�̂2y1A`�hLJ�,��Ḗ�D�ܚ��ɠ�,�d�ٷAf�@�O�m��u�cz/X::��\��ԋ�ʒ#�����m2|�?G��U�nL�bV������ѡ�m ��\�Z?LW���L}Bn��{ {.+Ȫ2�X]���#��y���Bf��d��(V'��$>��\���VL�z~kk�HL�n�����><����h���.�i��h�`GΒ@��.*k���$��w�IZ^k�-+3l*����s�N����Vv{u�RJ��՟�6���_�m�6��X0Z�O�=*�N��W�~o߼i[\$�c��<yh4&!��˫�e����Y�ԙ����P�9V��wW%:�7Q��2����F�2i��8��d���&��x��P��~Gm�>Y�3�׏�J]�X~w݅p!m�R��'.%b����(<�I��J.�M�U����-7_obɻT�wHG���4��lɰ���F$�9�����۞�U�8iEQ�[��������(�g�����ʬ���v׃�ߐ8�*Ι�F*~��9�}��OD¬���������q����4������H�3����(3���$�э̑��E�sfx��� x�<"K|Pɻ{�9`�����f��AjFF��$A���e��]���������;�wZxNcB��) ��Ջ}=�#��*�����22�]�*�F�ɉ��@@��vgⷉ


`U����qz5`.U�}�@0v���atu��+�3���+`�ZF��u_�N����L�� $HVZ���R�x*����������(�3J�2�~9)ʀ��S��Y�M��� 97b^���?���ט����8f{�۟R�:�����noh�zW�[�]7��ȹO����Z����r_a����Y��]k�H��\�(�T�A˫aυ.��F�hĲ�_��u���>���5*rFM��A(E`{� �y� 6v�����`#�Ĝ�˓�/bj�����D�p��L�
JE��`b�w㷓35���P���O���U
�&��ʸx#�GE��N��֎�N��Cq�����X��k����c�j��[z��)D�_oei�!���uH���¤]��*I�Ж�B^���NNN����D�^/P[:b��]o����2�:������\i�?X?��fA߾}S?�{����Xd9PT�56v��C�O��,�V����H�Utn�����sh ���qs��;��5;����H�?3��w���Qz����<��xY�Di*>��nSA�[
��܊��)-�
�|s½�o��ܸV���ȱBG������C�2��:ܭ��|V=l@�ٴ��H��:L�����*�f+�0T��!�V���	����;�|���ɼ�N..�/_�ק��Z�}�� C�`��߿&�N��*�Oau�xA�ؤ�3��( ��2^�e8�	���ߴ���vQm]]
A�۲W�NwD���| �Y�$���
�3N�?�Z�|�bl�/�A|W�vUU �!�W�)��̮[mݦ��Lv"вN��td|�@��W�gɾ�TX|��2\s�b����3�*7Dyy�}�͵P���*V�S*WU�'��,���jM�t;�ܪ��H����1��V	�_/6�hoo_�a�]�B���[#L��.w,�C^^��n�"�g�-QJJ
l�Y�U6��$��_���P-��kN�hq�:���ǈΠ ����f�	�Dc�p�-k�cR��
#L�/E>�ڗ4�D���$N�� �[��0|W��+/� A��EY]=7��A-����e	�|R�AģPq����د_ �G���������wk��>s��wY:�:8=M��_�0C:*ߩ���n'��n�.7P%;B�Ǡ�H?����H�=����Da�N���(�\#.�QJa������ӳk����:��n6��e���t]ȿt�Z�?�kD��d�XMe�n�N�ldd$�U��@�� �� Ae���X.�su�d�K�q=���Xp��ѽ�.���w���陉�%Z��tF�b�L^߃i꣠����V�jrY:�~e_�pqs�2��ԁ؟[���ZE=8$��v�O���_,wF
z���Mg.#)*��D�w&L!�Y�WCԣ��ѫu	7{wd �~�9�#����*�Kݫ��3� SN$��Z���n��`yi��D�ivoj�g(+ �W��]U��y��Ϗ��,q�U)�>���8�J�t�U~C*o��`c��í⪜o���~
oqq��BH؛H�ft��ͣ>���9�*Ĵ�����e�T7P������_���Ͻ�����U��
������5�?>�(�3o�eT|�Ұ�Q�n�ߔv��W�L�1�K�C(li��|gz�Q&��p˕�ccc�6�8�����1x���^^^p@2v���m��:s��7�����BQٻ��CN�c�:�B~���'�y��"켼=�Ǝ�Pv�^�������>}�葴��8,�-�n��c5T���a����������/��2�ȁ�� �����Ϩ�� �Q=aY2;-�h�+�T���+��o�=Iɠ�p-��M�b�����*��'_�>0�g��5(e�c��ȨX~X�KI����������zץ4
����fy�\��`�����������/��Q-��1©�/�N�˲�ݘ�f��c
v��-������'z��Vf0��ha믋�G�<�x�&G���߅j8��r�E���Ϟ�H��ժt����Xa�6IIɴ��ۛ��[�G�u�zz����G&'o�����@�|��
���oJ��%��f�ss��D�D[tu�����%H�	1vK+�Z��WU�luu��݉�U�����ݝ�?�a��m��t��+�ҍ�|z������#J6�lٚ-�d�̊o�O��,��z�:��	O��e��Y�*yf��'��#{O:\��d�>��1�b�t5*���U�ҟ�����>�Ѱ`OW��'J�C��0���`$t����k�&WE��*��̥`�;*Ku|��PwO�����<��`X����_$�]��9dq�C�Z�������}�Z6t����y?E��-��u�\�nu�ot鳵�;������rdb��}���H�L����0=6��λ3ܒf�hu��6"� �ֻZ�Q����>uT[���ܜ��=R?��NR�
�r��K��:���1����߿Gl��ƛ^e�I���9����lk��u��z�A��+m��z-��ҾA��=�E�6^tu��P��oѩZ���,�v��y���;>���M�>>���I��@[�j��K�NH���$$%e�1o�����U�q��������W��|�*]��ppQ�wjmk^1�{�TU�]��Mɗ_'}�}>B��Q���R�)�	#{������仹��dr!!��Du�ն�H����pxFGFZ� D�K��J�f)}}⠧��%L_���Q�Oq��A������fk�ߔ������w�I�S��j�Yn��"���Ϩ�A����$��h1�� Bi�����>�z6C9�[�CNߔ��D�c,�X^[�8�s �u�@���=����=bUP{���Қ�����/��"��r�3�s�{Z�9:��(�\��sB�I�99햼�I���kx@Z��p�kd����zT�ٓ�/�y ����� ̈KJr�0ܾ��>���˂��?�&�>>vs_�m��IWSN�O���+~�ROʩA�w�{cO�k��|÷�f%�]z�Pb��h_i.
��?�d�m��VMY,,l���Nz/����>�]�:ي�G��[�w��˨�k�DǦU4�/����7�U{<�V��8*]�E�����}f���z�K���A���	����%%� �ŻYtuu��)m'�u��������(9���`7 ͸N73�������\�TS� ����,����������������}p�)55uoo�K��1��&���ȶͣ���H���d�K���8�55�_rrL��g�!��҂�L�(7��P�-��������?�泥�z�,�'X'���-v���/���٭�0{Sj�����{[ӑ�|�	��;�'�w���p6�J�@�*3��_hZ�m��}xzz;-���\E�MF����������i 48ã���*G�kن�뇨��m-�����g���q��gk]I].��6�;D�7�z
�ݕ�](%%�2��Iߴ�D=����6�eN���OG�l�`X����c=Q☯�&7���^�;eVV�I�޺�)������S��vq��Gs��<<��#��VY)i���|����/0��Cѡga�.Q�S����������BEHH;��8�i/k���>}�#oaX,�����(��c b�޾-J[�<��Q��ٻ35b`�MllB�:Sڟ����6(�e�M�@ڀ��$"*�K�@CC�M?��Ҍml.������u,��ddd��J���Fj�`���yph���m�2]g8>+Ƴg���#�5�Q[��Ǒ�XJ*��
�L�)1Ƴ�Pl'wwD�A�_c��fe�����}�b�A2����a�����P�<#=�v���O^%�
�S^*Y���v��B6S�����k{���h˲P�{��Gƫ'G1ǹ�Ƌ
��G*_�d�����\��|�u`@�,`�ZԝYa�u�M�ZZD.��Rֲ�����T��lOt�->��$Ĕ�̭������Ó�2}Ҋ�$�BW��Ɨ�M�nD��U�r3�ka�յ��k� �>3�-f��$�~��މR�0��ֻ,�LD;���u	x�������r7���L�g`(lw~��Ћ�/�� O}��K�l��Ay �䜜G�zuN��Qw�?� ��� ~w���l�G��l,rH������Ύ�2���n� ��t�.B����E�D��tu�z���k��w'dڧ��!��@��_߾����%��Uuu��\7�e�k���,�wG����&�FP����_v�V��x	:���3��V�#b���i��t�`3\����b��;Z=#O=��<���Ѧ7�u����������Ɇ�gv�E����s�2]BH�h�2���Ps~uq����s����?���X�񷝨~H�Zx��@���Y���I���y����L2}}}��qU�%�8�f��sv"{�D2��p����2���_H�Mj�0�Ϻ*
"�	Ϛ)��^���O��^R�~�wp z��E/,<|8��]c;�6X=Jj�vg�l�!hE~:6�A��4����vt�	z"LWZ�@�\��/''')�]蟝M>66F0!�U�/�h��ֻҺ����iyx��+���p{�����ۓ�n��22m �=s��p\l&q���hi�>A�|�{;��5�D��Т�n%�}8
X��K�����<x�Ob�OJ��+))���ՙ� �=N̜���j�l~}5v�:����9���J�80|z�������OT�W!��N�;�[�������a�zsss  ��v=��6��tQ��O��N��Cݓ�Z����k���ǫ��g�el+|A`U]����(TWW�\��ţ�����Kb��7��R��>��O2�}��^>7��z�GECCAAq��Bc�ţ4>g�Q>��h@�\�Q��3c����Ӗ��Naf2��jjjO	���ʤ��龙6DE�%0����b'[Ș _����}��"=�K?q�Hi�```<��F��C�$�ݺ"E��j��4J�������������(h!��4�����\=6��P_�`Ǥ�V��8�4=�y�$����7��S��iC}��Z�$������)8���H w�MILI�8d��"�`�h���]����/&s��Ǖ�<$�z��9N��p0�W����c��͞�Nc���ſ
������*ר�l�W��L��>}�ŕ�J6&���1������Ӕ�����Ο���u�4�4C"#�fj����>q߅�l���3�ب�RA��IP�?����)�^fff�����o_��acg� |l@{�<c	
xA"������p|z��`���]�W*$��\���+�Ya3� �Dvŗ�@+���*���8�� ��1�X3l��:40�����`K���_r�� +9��3 �u.�Ȍ�K �1��?ʹ���$x' f�]�?x�=)GJ�
�ѷ�T �cs%�D�� �LUT*o�q�&����Y�*�@(��G
�\$O#�CP�#X�OF|v?"��*�����y� i! {�K�\��0����Й�(\4[�a����Es磌��W$
��!W8_Qw�\=�|�����0��PTӣY�hggN���L��HE��J�|�
=���I�Q$((���,���D�E��ᧆ�$u?Ƀ@
F��6�ְ���+ / ?���
�8�b �D@\ _�wN�) ��g���`K����gaa�o������:'#���W��}�ޛ��ֿ�<�q��NHH�E 9�F|�ܰU������;�:�Y�"������P5����"&�y���G��Z��	`��0�"؁�D��AQ����R��:�b��@`/�E��#d	�/��f�{E�?Yl��`��<�Yo�]kML�e� �m�2]@Q#�����$]�Ɔ1��)eJ�zπ
ku$T䀟�ك��\�h�Sw!�3��]�j�} ��K�,fik�B���Yb�|,bdr���� �6����0����K���$[u���� ��	$&��9S�ʽ�q8ob66�Ă�"<��byf�H����Pm�65��x��V�_���zaiw��}��^�(�STT�&ow��%��8?Z[[���>c֭~/M��IM^^�i����Ex�&%%�2}���_B�v�V��1���3.ǹ$��IA��:�Ho��<�P��BBĚ��.���**uvwsd��H;�o��Y��*�T��'������o�y|=���aHJI�'��C�~/.^&qN'9�Z�@�"ޞ��5i������pХ:��(����u�6wk^kk��
H8��8aN��l�暞g��S߻w`N�`�_|��Z�݄q�R>>B+���$A��M�܀6��N�g����Uzz�����@�5�ϱ�*�ڽ�=j ,��:�VU�	}�l��X��}��� <���������Le]�G&ff���@$��F�kP}8����\�(�b�P�X�����c��R�=��iF�B +�w1�{s�� �����ǁ|y�����/A�i����/L9����<����������U/���,���i��V�U[�u��NӴ&'�l�<?ۅF~�q*���?�yW1�?SԲ��/j% 0ƨ��O;�T�B5"�;��{���+ׯf)7Kh*���od��^(��k�M���yd��edd��M>ʻ231��\��^�5é�KKK����_d1D	xK�Z�{F����B��[�t\WH��:��{{���CCBK61Qa=���.��,J��8K���t��jdb���/X$�ML~���K��)O�����������{x� �͠�:��S	{01?�z��O� (�������ag��OU���Ĳ���W.�6	���}?��og�x+�����~��0�.�Wes*�Z=O�x��@�������ދ�g#|��o��Ҩ�q	����x����GRY���$/�jk��x��+V; ����I�����V= S��/��G}Ā��Wr���5vS||�,d�)v�#�����8X��t�so�{�ԥ�jbx�����8��� RAZ�e�Ǯ�Z/& ������b����n�w[��|w8�z��g{ۯ*W�,�bZP(�VY����|���������*#c1l|*�vPk������_=�ؙ� �M���K�Y����[hb�Ї�����ְ�,%���''˛��¾��/��T&O^����Ƿ����{����P���
^���Ҳ���n�I2��ƽ˸�; ��Ɔ��Z0� Kiz{������������x[q�k�?|�8���㔊vg�eX#��jȄ�W��a�&�F8�'��]ܶ8v��`���@{@�a�|%���"-80�D`�����%�2�Q�&H_Q�[�~:<��n|sD�wy~H	g�ښ��$M����<̅]�WTT,.�}+RѤ7��y�L�`�a�LAA���і���98��us8�HJ�֖f�1j���|��(����k�+��G�`/�y�������H;�f3�84��^x�#kJ�Pl�B
pעK��=�ޝ�r{ L!dln���$�>�{:���O'3����8}@/�~|��W��ʃ
��m�M����S��]~NIA����'���<����&K�0II��҈"!�D���:ou�/x�S����v����������:~T�|x�޻��D�*,(s�n�"�
sm���m��E\����\���nҨ�9����I����dq�l�몕h�Ru��O�F������v�'s�}No���_e�9���#�˖߅�(��<�о��_�����2w���1HTo�JQ�K�3��1�p�7���~333�nj��Oh������\/c"��*,��)|~ݳj��;]e�nw�հ�׫�?P���  �����������[A �1��.��ݙ�jk������|�]�#}����~K�M�������x�NU����pJ5�\���i݇J@V�9�p�l�D&sZ���f�;C
$D�]bB�)�v�{�Y�t8�p��p�`O����ECCC�y�n!���m%J�[�C�B<�Z嶫��]�	�,�=�GE�>bff�\9<9�:?\�;��W���r�^f
�}T��<X��)bZ=������W�=��ӕ���Fh��L��4��t8����v�$K�gêkj`��QsZM���#�J�/�>�AAW�vy�ɸ㝕��Ѱ�� hHD���1��w7��������=�Q����,�($(���Q,�i��Srq򆹽Ŗ��S��"ے�6�^���W�����4˕������)0���--���e@��d�3��s.�L������1�QI�4��_�r޺&����U]Ĵ������lr^����p�
��6S�ث���E��m7�8��� e���B�77&��T'����;���,r����a����K��狁�C�kV�⇈�m�5I��9��ȁ��Dv`��}�A��m~�~����F�����}5_�m�	�!q�P]�0����@3���II����h�}�,�Eyǋ��D�����k��j���+--�D�������;RdO���')�?ϝ	��?~$�=�d��ZZ(���Y�C'<T��<-%�d�����}��c��
vx7�8�7i���޳����~�P#����`X��AB2��l:9$�6��g�5��b[\7zhz�(n<?�"}K5��.r���W���X`M�����ʊ(k+�׿�'0�2�R�A>��*'W����͎������;�el�X�ۚ`��z�aS�3@D͗\�==Z|�*���!��_m�������R-��~�\	&��L��;�f)�`Lޠ�37=�8��9C%��󣌑;8��s�&�+ه�n�):��q���|���Y�����G�s-b��h�����tz ��������'[�)����+k��t�ÿ47z=)����ٲ�j
�唗�q�O��H�<���
���˰��i�|sN���dC�f��C�hKKYq�6�G�,u� �H�hc?����H��iii)� ���l����+�!�jj����7���o�����(D=z$nn�+jh�	�u� bwVy9ƃGO�ݑ>��p�2�#5�u^�ô���N]}��uH��O�'���Ѥ/�##Q�_ F
�a;:��	3R�;��t�mw��H�NXĳ�� /ه�9��=�w!˳�V�����ǡF4;�;Oc�#��gb�D�%���>FE��������^XV+�F784�ki�8/���X
��t���������x�[B��u�Ȑ��m��������&��I�W���&��}�\��VMŤbmM]�_3�H^��د_��re�%-�}|}�u�Z0D����%��}JME�x����z("D����m���ޮ�&-�M�����Q���<�q�jϗ�>۟aiW�"���=�@	��ɡ����>����|PYU�A4k���S�Q�sL}��~�'ܶo�����k�.���W^k(��{8{"���������5W\7�.����<�)���4�$p#�IT��H���&_}I�#Lx���9������C�O4~"�ɯ;�?a!
z�*��L �������
ӭ����W�E�׵���}��;���*�톘f��ޙ�T��T;�BZ��N����[H�tSޓi���D��Ʉ n+@��Lɹ�����L�G�r[:y}}��_������H��KJ~l�㪷����ȳ�qxYh�����N��74)ED
�mK83�͍&������5Zf$��.�].
��vpz�$N��='�S1��?/.���Mbs8��H.=F�IK���W飛��a6��!�5���U�R���.eV�׉�X��3L��������"""�7@~�	LU�j���&�U�tv�ܵ���h��sA���7���^���;~��Y^[��su�+7�+}w.�'�(����؄
z��K��gwgdc�o6���	C���4i�8\*���}qe\�X�FG?$&��f���t�/w5&���Ƚ ���>�ǃ]��`co�v$2Adp��A=աj�âN�͠����}0�8^��P���%K�"�nu����}���kh���6��_����`E�J�͛�B����Q�f�蹟^�T B8��W�_����0Zz]�ɬ��ƼU򍵭-L�}�����w��:���JD5����\��!�<`�A�dQ B����_ܨ�~U��e�a�},������K\b��������$U�++�0�6���g�R}.�s؞,�� �����_h��r����#�����ˏAl�!�� �[�Hᱥ���ƃ���"222�?#�~f�0벲h�8Ԧ����B���Ɇ%+Ϗ�(aI����iR���7������ag��:i���Mi�ϟ�w`Z����P+�����-B�莎��N[2��yj`:?i*��%ީCJk}��$�J<Z���M|�G.@gz�0NPxxx�P��j�U7?�k2�i|�1!��$u�����ɰ1Icqw�VJ]Λ�FЯ���[ $ⅆ���ӭ�{AAՓ�?Z7��N�׮u$tR'����D8����P�e@	�Pq��rd�ۉ=���:���"v6 �Y�}��A��0���ż�Y�$�P_�+犝��W::���&������'[��)��ʢA������&���9��u�X�� Qx��w�`n�������q���y"�t����/�7�n�`.���n�F�" �3��Sɚ��$��wnV��Z�'A*<�l���D~ �VskG`� �VU��%� &�ʇ����;[v�'��K���f=��q�V�K��4�\Q7|o���S[6��[�'�b�AC�m�@0F��x��A�	,������g+� ����C����w۞T���,���H�E�ݾ�����X��K�����#�*9-�33D���啕�yyԛC
�ϙ�#���P��s�
�ƞ���Ww����juv��+�����
3$��j_�����42��D&���l��yE0�|�vx|;}`	�ǆlg:�ؖ���x\(���c��FJS�x�7�E֑�X�·+��x�ۓ�p�y<#���ߝ��11�i���^]�D�6L��vPI����I��:ޔ�$[07?_�.;Y5s�9''6$���鶛!j�,4��� �e[�T�[�>�����X�����pF��D4�
N�M��mO	#����|�"<�����a��j"ϖ��
�UsdDA���_�B�z r��XCrs��//�HF_z89���*�;�� �_*l-�����41f�g�/�=��[��GU�����=E����3�ħ���m�,5н�������ET������?���?�u,�=Ѐ馀SQJEu��Ů;�Sa�Ïj'�
�<Y^;`�R>�������oO�������M��>~|����_0��Pf�"yw{�>��<�[�>��\0�v���y����.����ON&��Y��~B�J͞dI��/ǁJ"�c��!''GײX%�?Y��uB���ɀ�4�0W
���r�����@ ?zJ�����>�_ F��o����&�rY�of-Oڜ���y�NW(�C%ۏЍ�(� ��!����"	�#��'������H��*��R���(x{��b�}����N����s'\[��}��x@��d_��+;� ��&ڐ�q֏6F�7o$�0���Wc2�I�R��L�R��i빏�ݻ�ЖX�W\̤x�"����xzb7U�6;����2b�_P�cnN߁�{���R�ʑdֵ����n�3X���R�oɃ[����֣ �cbg�F��mSwҒj���������N��,����ף_���! -���Y5.W>�O~ѴuJ���dI%&T�E�z�k��̉���>������-��H�R�}F�KE��R2⥭-X=��|�8�La8�e�l���F
x=|���拯�@�Eҁ���HQ���ܒPa��| �n1���03 ��sW<�0?�u���|r{���6���@0A���%�ӝ>m�����$v3�(��#��>�;}l�g�� 7g��З�a7���r�I�b٦o=<xLMMq�/�.U��R���u��/(Zani���b�v�5&�?�9x�'0ŏ5��:���p�-<[��Xõ��(d0�����_n�[%M�/���6�^�����i}����^���T�[�/s &�� �*kk�����@�\YYu�:��~�Y#��	Z羳{�T}w5���!)Jk!F�^ﹽ���}�u�Cv�և��OH��t(��t�B�οC�n��,f����Ր�45�-Y,�{O�<��p���̵���}Č��$��ű1�����˓m\��o��K燫N�ί�Y��n�'��@����D��>�{�Y�t��2�,,,�}}�樔��g���	x�	��Qn�F�/�C�d<;o0)��.��'�A����4HW6��v��n��JI\Bb��Ã�3�s8$Z�� ��u���l�|� v>���u,O�z<��nzzzic(����&>~O��`�е� ��\�A�]��J��B���_�LB��!GS=����~� RZ��;{{� 4���2#�h�����-<9��OR^���0��ӊ��q¯zE@�^YE� �>�'Z|�)�h�0��=�䥈y�Ã\P�ɉ��:���=l�h��.�P�P�(���a7�*��|zJ�&)���ֽ�Twr�$��ʅ�00����E��}n��j7 ����r�>������>f�y��?��H^�g�p��p������7�o�~���,nK��j 3�aׄ����.���_J�U4H������ք���E�o���P����	Nӆ��w�:0�ϒ��h�0�L���1Z�l`m3J���3U�yȹ��΋J���f;+��xF-xI��|��u�G��GK:�?[[{�xl��?q۶��]�ݕ��,M�Z鍡�G;K�ae�;��� '#���Gw1=�g��V\�@��=�� �mAUww�=26&���|��i0�o��fG++$AAA `�L+ � ?�9L$;�P�Nq�.!!���t+؏��ߜ`Q(���稸�Q
���ཹ
�Q�8����$�	U��g{�����h ��J�4�������G֣�º\EH�4��9%][�[�6� �o�Nr�\��m�zX؏u���/��V�*�9�T�G�������x�c�"���zJ&L��o����Ѿ���]���Bdm�pF#��R��]��w�>��[�0���z?�Z�B�f�}��v�⟖s�M��o��tq���:.6,�vD���7x^Tx� %Ճܣ���i��d�3#"�w��5x�z���*`� ���
p&b�NR �Ϸ��f�ÜJ�����>I�����Yyy�r�,}�]�S
����p1}}bS33�u/V��6�Y~@�A�z���z*"""���8,[s�%��T� �<IK`1�)�\��3��6쭉Rvv�%#J��&�³)���i����)^��n�*�lㄈ��Y:�d݃���(递���v�B#��+��p6����-$�DH�ȯ4�t�	�؄U�E�&��r�p��#�X����D:�91�D�\���+vR�
6�|��j3n���hs�ٓ��Ju�#���O����7�ŇF ��&���$��^��fNeÝ����ň��xw�%�*N����_�d���z�܁��+Dn�cg�qێ��*5 �l��']�AD�k]X0,�^hz�ddd(�
��x�bF=n{�_?&.��:���uʲ"@%"|VCqss*�6t.���%�E�����s�搰�s�
m�P��[ߜ��Pow��m�b�$���Ty�>���E��[������_VT��+-�3E�r$#U����/�tY�?(�|���iok�g����}K��V)ôxI���1�%<`U-|/�~�O�"�|;� wy��9wfy�/)�+���Ҳ}�.�4�E,(����O˨�k_=)�b�x�g�p�0�p��.�;�(�qqqQ�o+���dmk+JeZV�1�ք����5�5>��0����h!�(lU
�u]{�H�e�p����fZ�"����j�Є^� �98��L�onnN�7bǝ��Z[[3���Ӭ��5�B��zpp���]���"<���<3����+�����zc�]r۫3*9F[�II��S�sJ	�t��D�oi'�v*[l�Z�o�_����#�V���F������Cb3nEl<O���nz˻�3S�YC#A�t .��s>>�(�55ܛv{s���a�����՜OF\�Kj�<�y�����x&
m�-Q)��	��1��<b�d(( �(�~%������%'z�Λ������a)�T�r���FG� \��+��rxxH ����s��ȮS�����H�����f�u ��zWVUF2��/����և۬�-������%������N�E�&S��h��H��~D���N�:@#�ł]9�
���YN�n��ͼ3ܚ��nx~��I���߿��`tg�Q�w���� ���5��C�Ǫ�\>�$|�l���w��Q��<iq'UK�m�3S7@�1QW�^YU5h�����`I��r��M����C�6ua�޳�*� �КN�kQ��0(�
��{�J�Õ���{7�1��&@+���
A���{�",|��V�𵫭;��o����9q�*�B2�ФQ�gO5ok��-���M\|�s�P����������D���J�ml'�M�/�����w��u������m#A�Ezc�>��qNNN&���B@@`|{}э��G`�h�
���h*�q�Ӳ(���t��#���,q��#��֐{�<��c~���=%�&�fff&�T�z��hb$��[�[��f�N�L[},L�{�&�54����G`��*|n0�����;�����*��A�2�?��G��]z�my�X��w!��a
�c@�f��Z�����LC(�_�-�31�z�r��6�f��Oh���y����̈́S�%��]�.?U��,�`��*�m�':45���Ą��|ٯ99bA��$�?x*N�r�I��'	O���^F��[ h�*+'G	pJ6�L�;P��=��b�upp0�?���y��eɀB�?!_;X�"M�B[5#�uL[��(�$r{NI�gZ�KMz���cquuM���$�����F��󻊐��b:Υ���j�ٿ�c���{ ��ӏ�:�Ô�?�C<Fդ���y����333��_rrd<v�ޑ�x�x?����B�q�}Um��#i��}��ToOw�w��6���ÑT���^~�G}CC��i��rp0�%��!�v�k�n�0�Ǿ{���/\�d�~ٰ�[���?�l~}�3K�WP��#�LAV����[6��z�yw����@�f	e�nfkG`ߐ5��S`�ti�:$O*#�5Y$DD�I�Ȃg���� x��χ>f�O?'&��!�����M抉�����oMDD�9:�3[mnaA�����D���w̩ɬ�0~k>p`��⍨�,��邞4B�J���l���wS<]AL�����؝Ŗ��o�w9㥩֎���X#+B;��R��p!��Qa��V�q��䔔�_�|A^��}��;w�Ӭ�3�7��=h�����j&�l���߿1@�pii���.�#J
�*e���N�o,1ji����_^=����t�qg�U����o�[�/:���]7�驷/Plll`�\�ԓ�!�w���w������1a5���n��$���Oj���^�2�V����ݎa�������oO)Qbjp��Z�twVJ��x'����8�� ;�ݥ%:UA�'6�R�h���d��b�������`�g�o��������؄�0)%�^l���PJ�jkK��>�JpQS[�5}���-������A����0g<V���M,�A��'��mV�\���lS'�\�Bh(���_�������>��\�4x���RY� ��' �pӨ|�����"�p�0����8�����/W���GҶ�A���<���9Q�����M�Ζ�L-Qɑ�����
��MHH�����_0�pWq�tu5�9�w\h,8N�]ͬ��M���]Ns��y�^>CH����L��EtT�����&y���-���f������{QQQQG ��z�r�л7ӑ���mu����t���	֋��|�:ۿ�;�E��/���	^��d�ʡ�K ��g>/���1B��1�Ks��s����Lݭ��֮u�b�M�Qû(��Ҡ�GUU����ρ,��M��-/�TlА�#�~�	VYs�����ѽ�Q�[���uo�6��4~q&<�[���p�__�IyS-MM)4l��V���Ɠ���C��̉]uu�ع��l#{{�%��߼���[yx�%*]e9d�+��Г4Z
|<!	c"������Z�,,)Fݻnil�r���g~Z6����4r�����G� X�{C�aT�Mj�R�������[�u4��[�{���v�X0���A�4�:}��xC ���ˊ�r�K~�&ff��ۛ�J��^2���jKZ�TEg��7����YS�=����"&D>S�����}��A��C��'�N����@�X�6+�tUW��Ⱥ�^���ރ8�m�ǹ�� �5�o?|����-���z@�#R��e���(�c�D��/0�|�Ԫ����+<2�)�֒CS�����{Ϩ��v]��.���Р�" 9�(�A@��snh�ˀ�&HNJ�HΠ����$g�n���w�{���q��q���gUͷ��<U�s������8Ejck� D~¨.mq�� q�xW\�6����L�`���S�O�K���a �Y���j�L	㠇r!%�w>>��SP�(//�9�$	8}bڕ4��o��h�����~r��ݻw�~�h���'��=<-�f��x����l��p)�o 74��aր��Ҕ���d����*0���c��И��R���n�Ź�\��Щ%(����xʂ��̣DԤ`pn+��#ww�z��C!���k�o,�|}����dGY1��M�SС�[��� L�ruk��UAS%��˗7X�M���"$ۇ�*e��9�⬎kz�SS��{')&�1W�͇O"�l�Xt��7l%�@�G/0����T�h�Cb����"�m��v��
�=�,M>�*W���q ��tr�Bu f�j�L��Z����ʊ,j1/o�`��	b �s��3P�LWL�{�̸���T;Ϝ��U�|QS-�Nf���0���p&!)���ϸL $@�j�7n�x���R_�����?7J�Sœ8 .i4����(�X3�ì�z���ă��ZN�I�Z���7�$�ZFUSﭮ� j��u|Җ߯TSW@,]4pʍ���6F����PD��X���0��*Wh�1�ɻ�߿��'dg���f����m-I��)�!�����b��	���Y�7juXxP[f���>�GGO�u#8L�#�H�[l灓4^�P�. <�30�:�t�o߮����`_�vz�A��lcs��������RRR�9��o�܅��
����Fz�U���3������3���В�L��Լ��A�5ee|��i�����\q㺧H�S8��m�� Z�dnr��tv����op0^%[+E�(�Y$��dY��?撥� �Nz��9���|	tX�=Jt�z�+~ ��߿�gW>D��pQFF����˸�,�V�kv�΃�(��
���@�5��@?�*V��YZ7ˡ-=��G�7n���`�x�ͷ��}}�}}}�oWnuF'Gu�������w���s��e��ͦ�t�ϕ��<��{x	���fkk��O��>/��gn�7.�m�� ����c��9����B�w����U��A�C���56h 0�Ct:0=k��(u�o?F��D��u5�k�S�s��}�Rؚٸǭ^��cW�'xl��ډ����]Աb�k}G~��w�Z�o4�ih��F�F�ݚi�.�6,�vg���{��9�*�?�(��DP(��f�lU�G�z�t��aN���z�|�]W���u["8VG9c�=U���zz��r�߿o�H�\"c��p�y\`��ƅ�B��=�æ��A�P�`5nw&-�ڢXuzbq������e=Q�4>!a���row7	���{�Mou��*B����=V�{: c��zGX��P�AU;FEI��ot��x�ta<-=�w���~?�^9�PE[�y�XO�n�W��4���5J	o��Ni�?<\9�C�jM�L-^�ܿ�k]��X\�9���&����TE��x��DP쁞�H����^F�&����m�y*�V�����|�ʘǨ�>����
����v%)r�������1A� @V�ri�\R���Y/,p�q���G�������� ��bݭ���i�/=9L��UV
�RW�/,��n�w���Qҋ�� �x��BϷ�3��66��F��*���mmm���
	��d���b��f�����;�ݓ����Y�jν��D�|��i��/�e�	:U1�>C-o|���a��d<�ƣ:fW���B�""륂^J�
@���&�ũ&+@	&��z�l+5�+����;�
��x*D}�T{�U��(�+HGٮ߱S6�~�r�ʃ)fL��fuc*�/pp�W��ϊ2�Wōj>^Y��t�^�::427o��rg}}@�%����V>����)���y�����B��6�u�ɮ�M�O�sss�~�}N�-�24��&�����*=Y}��� <U:��|o��nm�yM�hC6�p�!���#�r�[�Xb;� �&�J�c�J���z�3�/q	yyy*y�����������*����#�h�����Ǎv� u�
��q/���*�RC�aLx���nCA�V��Lt�!���TKG���GM�k����.Ȏ�.����z���l/�Oe�� ��> �.���di;�`��P�Y�,z ���@@W-$x�!=��r��r���$�
6�C_]~_���9���M���t��!��#	�Ċ
���S�+��Cԥ��A:�IQ���`�-�*]����$IGv��1V�lk��F`T�q��^jZ�sJם��%?%��m�EI+�p��!�js��O=��_[����SS  �d���t=�*vU�����]��pw�v{����γR����!D�f��at�.�&�Qzv/G�FPWo�!�}?�'K32�uo�e���LuEI	$�su���6C�\ 2�F �X-G�QW,J�B2bu�ڞ��O�޽�6��t�jP�XS�e� %Z��V_@e�G�ׯc�V-E�,�B���d*ףWh �b�N+d�2k�]Ps�������0������V����2����p_h�a CV�=zff�A�k�� �ꭎש�Su!����~��u�:���h`�P��'�� I�0�r7K�=��f���)�v�r� [�baa!H�m���' T�Z[���3j�P"4$$$E����.ƨ��Lƒ�8��Or��!�$?F7��1���h�K��N�www�g�>|��Ƭ��|FU��C���#\���.}^q�ਡb{$R�i.�}S�y\�M���o��W��@����S�)d2]gª���y���Ζ�K���r�(�,ι�T�1á����хs��B�9�Rn�S:N����mg�]7�%�={v���_��B-�\�R�Ϣ�!3�,S���$����AC7��g��5��H\/u9� g�K��g�Yof�v�bh�"at�ݜQ�����g�R�`�7s�jd�(��*�����\���:&]VP�?bl���::.��Z�1��6�R� �1��b�F.�$�M5(�h�ǎ�#ՀHk�l�D��w�m+ό���f��Rw�3%�� �x�S��i7��B�7ߕj�'9�r��[�-��I������L{2x�6��yBS�\H��{J��}���@���q%/�
�C~{�<\E��}�W빛����Mv�K�[�t�a�h4&ʦ���[L��&.���'is�ۦ�ީ&�4�}��Diz���������[ ֹ�qa���í����L]i))YU�{�S��2K<���4�G��A �d�����
n�t�w�L�(�6�`;��{zz��lU+�kh�� >������E *�� 9��-���b����YR�D�����e/8���ܲq�����:h�Vnj��{rXs�;�T��i�s�<R��VO�D�_W����H�#���C��o�|p�r�z����8�՝	4&M9�u�\p!#Og�g���<`PUOL�������,��v� ��7����M�ʻ��a�҇�e�����u������������<�MS6�� O@���D����)���̕;:��ri �p �'>3s�+��R�2�wCz� 0Y�U�l���X��* }�hy/�%c�{Vs�.� �ٮ�7����ڄ� �+�ƺ��&r0�|�33 ��,�X�.�hyFDD�4^�ٛ��=<�ū�`w}b�S�?CW�ioM�B�m-H�T31(�`c�y�X?��TSg��o�����NW��M5A��WW�D��?�/-����{�Owb6�w��G�] : ��kiQ��wt\��}h���� T-`��Z�i�֪y�4聴�w�.ԗ�<Fff> Z�dg�!{�fW܄^	�o�FMY�$9���E7��N�@utt���qqq��cbb2i"$$$��ШD�I���{w2H���02�#��jjj��*yv�I��)�o,���_ ȓy+�"�
�������}�`S@M<>V���V̏��W�!fpd��{.!Hgoc��S-����$� e��ꪕb� �������и�T��	'�4Sm��`�n�@Q��~�l,�b��/�OpP�T̆K9���� �Z�рu��>?~̘`��ѧ�����"��RogC`����U�����Q\����e�`
\�+��pZ�8�r+�~����
�FΧ��:2k9��p���_uu[��2)'����
�mB�{Zj�'�z�����<����sP�X �&�7BS��Q��)))�0�z;�������E��pom�7��z0��565A/����de	Zi����C��CM�(� h#KK!��0i.;8������ːa��p,y��S"���C�1ݥm/�ܟS6j�'�a�M���)t�	
�ho�bu	���W��}?neq�k�/����7�l^g&k�/'�I+���Ͼ�`�?ج��fQEZi
�-�����/�t>�P���߼Ғ�<Řc�2�������O�Lur��M�<Ų��32\��ƾYlO���nu���C~�RH��N���P�C�CZ�>i�-j����#�\�hR�t���J|K�"W���ϟk?�6{20E��n�Vem�_����RW;�ߐ�*.�*�����]ɖD��rf"�6�-x�"ig ���2��XL���M�-�)Ԍ��$���@N:g�>�C���BM�����f1����p>h�3H&,񹨫����p#U5w11#��Lo��0h8��[;�Aq��8Zh���Ό7��ך�9��4���ks�_��D5*��o�P.CG����X^�p�ni7��.��O��*�m_���f,k�l��O�@�{/������ὴ���~6�����⽚����OZ��Ri���&.�l��Q�l��| ��D��,��m��qW�6�%�.�qً��+ �PXOE���e|�=Uy��Њ�f��c5����qH�O�gy~��&�T��VB�F�m��ړ�.S]�u��<��/����glJ����|�u$ȵߥ;��Ö�w�x���9Ẃ.�SM�.���Gؓ���ɫ����q��W3��d��XW��ϸ@v<������X�g/�\�\1�qi��N.'<
���Ȱk���3R�r[N=��~8�a����mv�L�j�g�I���c;ǽ �v4��\W(�ۜ��z|5(�Db/�b4�%�-���:(�̋����Øk�-ZI���(�f:Ɩň�cA2~��4о��M�%Q����1�����$�z�S�.�����9#��Ҷn����F/�;&ޭO���?_Ӧ,�k�(��߅�۪]:j�?e�^�z	桤?��@L�o����n������w���@m2�S�4_m�3l~t	M��=���#�q�E/���u|���t�D�$�B�sR���
&����nR��?z��B=�z�S��c��t^h������s�C䑯.�hV����"#k$(�oFXW[]*�o,I�\ ��O����px Q���^�����>?55ł��cfF�8>�4��G�x)!�|%�� 1�HCN��"�~��@O�buh�>H_z�����m��dS���Y�<ݙʧ*��i�4�x�=�\o���a�m�����p2 2tk�� ���Oɘ�!xU\��G��xn��&�[��0�[9Ÿ�A�%�p� �L�!r�8��ˌ�K9��1��{*��C󖓃VѰ�z��w8 I�]\A�E�� =�l�i�XO�4D#Y~�E=�v��a���D����A������XG��y��ՋV|�#�	���88(���6�Wǥ�^ �|)9D;�Hc����mU��uR&�IDέ�\&�캎�y��C���nwd\N*Gwx6r/���"���r�v���0�M����2.Vp�|������֓����;j=�9 .�Pf��":��Ãy�՘K����3S*�����=,�{��;�[?M$�ZK�]���vQ��s\��DLO�f�wV�>%�{d�3w���V�$C�����R2����64SU����h���LDV���FL������V�&�ީ�&�F�]��,1��o��B�s�(x0Fh��"88ZF�of��{Zr����J*z��J�k��=D %��ܛ}7������6�� �)������@��V�6�da�Kj��B\{?[��9�;�K�3nA��[ ����f�z��d�G�D���Ϩ�S4#�h������ >o��mk�G���� z2��β�mws�璼�-2���Y���w��
M�H��:�C ����Ȩ&�增B����^ I ���p���貽姯�s6GDF��A�A^��v̞���@F!*<kEX��T$�6FI���"�h�BD0ߎ�E��L��W�� 9XXxm�4���=�7!��Eg�)p.4����SMu��zsA�	��ܧ� ^�G��/h=-������%��	��iq@���Т����h��=����sfT�ap�6[���޾3x����>2Z��-@�F+�-��/�Q�����O����O�=�ۮ]���z/1�u��}�#�GL0�/�`n�c��b����sC�����#G]鶺9��~�Sp,m�1g�� �	�,��A2>w�a(V�B�]�r��٬�ɢ�;9K/Ο�_𚔒��L�'���a�|�ˣ`��8����j��.������wݚI`5Ŷ�*�w��K�166��d\��ȉ���w����+i���o�j��5P��=��\�1ET^�I Q��L��v������x1r�e~��c+�:F�hM�0���S,IK�UسGܱ!����wH��~��1]���t@izC�U8�2�5���'�(����A�P�������n�> ��h��k����Ԏw���]�u9�KI.!����mr�q����:�hr�EՁ���W3� �G�K�t�'��0<)΂��k/���ݒPq9k�^�q��%�L�EV�n0�j;�oe#V7ݎƹ����c�S����64DL�T��z�1B~a �fP�����;�����FP����0l�
͆o���֩RP�V�,Yo$��öu�e��I�\���{�~��.L'�K�B��	�v�T'ʩ|_3�<'.��[�_�����fx�S�1�,D�ٳ��hW��PI�"E�ׇ����g�6U��uuJ��,(�Z�����)��J��1(j�sU/�Y�\�}��>0p����H����(���a�}a�o��^~�6i�,M�+����1Co��'��}^<�Fw�!mKmME�
gM�;�֍�`�7�����q}Q��p�[����#�2���}]�ː��(qÏ���b�k�����d�J�_�W�#@B�Ǯc.�b|D��Q�?�ê�u��s3��W��p����d��+C���b�y3o��u�Yr�&�a�~ȓ�h<*����Qe˻�U�T��WxX�㶟,�����N�$^��n|�T��kB~>;T �����=�YM]D�����xFZV�@�F�����������rD�~S~�h}���C��NH:tJs�AoU��D�b� #��m��$�栭8����, ��t�!����@zϜ�d̬�b|���ȤB��P�5���ü-�(�WS�o&0������\�壢A'\1�m�zaY�Ȉ�꾘�g���R��7���z�
�hk'���2���7��#9,��"/A7>&S�b0��m�%*/��7���������,��ƶ��2	].�[#�y�'�4�@�9��_Zm,��"�����+6�1����08���`���8�\g~�s��6�K��
5�MN���r��W�uu/Tjf���x����бs}�Jޑ��cDlQ_�hd��n�;�
�����K5���E�����:յ���j�G�����6��p�<"�lC��z���C4K[�}�3���buLQ�醎�9$�������>� �%��c]1Z�H�zh;Z_`���p���i�� ��B�j������Z�8n����bMR�bo\ �%�1����M��������+E�3�b�KIa��|�q�����&��r��#��4j�~���;���Mj�PL�;z�E����B�}���Ts��ه�Z���/����]�ۚb\�UM��R����u�W����]��%�=����um�职v���w�b} N�,�r�	�]�n�%�z��<..���Q*���ő��M[�h�bdf"�?2�)�2���v�M���ə��b0��\�h�oF���M�,���Y�����"xv��s�1�J��=_u]\}���v�"�r��5��e�{~����B� ��G(����uP�ʁz��y2V�X�k���Kp��Y�5̑LBp��l=�e�AQ�W����d]���+v�$��T͍3\b"�3���}$|��I��{���ߑ�v�|��>+��#��?������5���xqqIO��{�Kyy"h�s~~_��% N�} rr�ZZ�}���A���	6�4�>�aΐ�=���P��S��mtBK��[K�����u�=��9z8�ҳ�H�S��^g�1Y���s�����{�{��S�R�kiży��z���d�l}���L�-��kQh�OQV�ڤV-0Qn���H �~���͡VP��B�������� ��wBT�v*T��h���fѐ���HWw���r7��h{{@cԈ���H�I��r�|��
���ߚw�����5'&&��3100H,���J*|�-���x��M��ބ������-��ο��6;A����}�
�M-��\�b�F�}��PP>?K��v&��k�=ۿ����@�,�C�{���5l{Lp�p{+s5��H6v��.4�Q��ۻ�+X�4��fp�٧�e�_��d�6��H��Z��x-��ѯBd���M��RL��.sR#[?�ѵ�C5~�x����7~�m����tq��4��fB��l��c�%o���e�H�[��c���
;��ѫaۖ�vS�g� ���d�:�F�c��\
����w�m�~h���$��h}a���6.�s.J�����f;J��@�ڠ5j7d�����u��_�~Ř�� �|\��MQSC9j����lmm�+�pN�jW �>��Q~6�����w����D�***�ؗ�(M��x�t���ϼ�����g�@Ob���O\\�(��8��'đH$`v{��8k���?t�:�;��N*���j��6۷B�� w�5zv�tW-讅��3_Fmr�@E���|��SVSw727G�*�״�P��<^��Q��[+��1j1����U�m�!� ��9d���v���_7���g�ZR����Wo�y�'� \u&��}$��g��
h�ν{���uw~�4M���nc���>�ò�5���ђڪQ�����2��j!mh�͜�:��30�NGRW����	�ѝ*Һ	���/b��ϧ���ee��V����3��,Ay���9��m\���O z�~/�PX�I*{n�� �Nq�G4���2�hvV�F)��}����U����||.<��}'�B\]Zn�zinn�w�{�꿰�67�JrG�g%���S�t���_rr�g�O>u�������~��2?P��n_R��a"��3m������)�ۭ ����S��F|2�g@�'���@$VPA~�]�BRT�{��)���<�O�;����B��� mI#�H��'-��[���xo{;�d `ƿ��^[�3� �b[�88RE v��߆ )�;�5�zg�E�3��=T@\��T�p���2��y��~�����WM�K������e�wQ��q=�#ץ����=�+�)�O�܆�Y.���/S��I��_�9؃Y���>�Hd� )�'�Р��$[%�ޗ��,p4�W��G��5��z�˷t\�+ �m���ѫ�yU^�7k?��z��&�0����H+H�ko�N�ݝ���W�1����М���1���K#���!->�=��*��e�oE���Q���oƃo�\���W��dh�Tk��������[�HٽX,�Ve��d�.���!e��[Rn۸�iD>�xeC�#^�7?��'��+�Y�4me�궀�q��9����y�8�!�	_�f̆CUVV�N?���6n^�r�_�m��Zz9W|�YŊ��a �Iv�xY�x�t��y=rԧSVH��g&*�U���M����W����v٨(�P��m��τ��3З�rl�OH�������-4؃�*�9y�� ��o��f6���[VN��30���T�UG�lm�F#�z�D.㤡X�N�����f�/��	�퀿�C��r��pi�J]�[e<f��`5�Ewк^�6wN���X�j�YuI]
��Z�WI�S~�
�������{�65�u�,�73�{�A���Y�,�|Ư%��w�a0����o@I�<:
�����^���D��.��oÝ�yݟ��g}��$�������g���0��:gb=d�������y����n���ģo��T�HC�_P�1�$� D��j:��K@_�;��r�:O��8ﮝx�����<��A�1�rЖpr��C����c[
?�j���?�H�]���?*��݂����e7w�d+��QPxr���:w"j���ʍ��M�X�� ���J^�m�B{�t��-��z��΅6M������=��f�'�r���.�`�?��� )����j<���>WG�mji��Е{�g�x�H�!�wp+n���)II
�����f	����+δ@!K���@�[,]omj#.�ޜ����'��{ 15k��
r��� �� �4T��1���~�&�\\���C�pq��m�;!��*�V2˶��t�?2A�<���pU�p�/�M�ސ�Y[D�:lm��{�H��/(�X��� ��S i���0iF�1�׌f���;���=6�EW��eE�f5;;{�Ī�tL����squE�C�U)���e��9��g�@{�4�ы�7���ܵx��ޭwI�0�\|q%%�.��ܰ�p{�H�|3�Ut����3�`u������eA�q@��΁���F0�3�;�Z��bU6�8�x�X,�y���#,	�}s[��y���4��ت&���@�_�#�?\"����Ji��nk
��m�>�9�R�cC�i'��3qNF$���_��AN�J�>���%G�ނ;ϖ>�j�r��=bM���@���E���� N���	J4$?����ߝJ�Ȉ�U�?QM��տ��/ky�O���������9H����ҩO^Nl?I�y�|����k���=�1�;u�6�8�����_�0�
�[����k$`��f��Z�y�_���ZcE��Q ���f���{PT��~�2���=�2E3��ؿ��4�v����Zn��f%�Bήڵ����,Gg'��nz��(�������1���bi�U\��(Z�;��l
��=&��rg����C�`0c�"�%�T̠���s���N��s�e\��(c�\�=��C�X_��HJ�?Wp�;/3T�P�Y�|�ፍ��V��Gr�O��GG� �F#^��4�?c]s�K0�����e��}�9$�:'�Ő�=�bS��a��a������+@ �^��Q�Z�uJ[�*�9G�qM{�Qe��( Y��z��'���%��0r�r�z_�^qO��/ *����-!���	$` �� Z?�/Gr��|B����+	, ���,�-!
P:��]�� ���n� ?�C.K��j�#|\���CŐ��Ǿ���_I���ۼ�fQ,+5 k�#�To�ť�/
�[Q%<��/��|2�z}���x�w�ȅ ���p��L5�v��(F��X�~ "�>�cn��?ɛi�.ʹCR`d+����PB�J� �$�����L�^�h5���q����5��c��)`Bg�/ީ<�2G�p�O�k�M 7 �7���Q�s���;�C��1��)AW�ߵ�/i���e�]g��#�W��{q		46%Co!��� �����[���z����=���� ������w��s�C�<�z���<�;A�剸�(qq�l�-����;�"|ډ=]w���)>��V/�Ò�Vt5Am�F̊^�	H�����UTྦྷ�t ����U֌�Giii���Q\��C�P�(���R�qC���XCӫ T��, ��RRMo���|nhhQmee �� 4���X�.�~���X��P��'tZ��aL�Y��GO�8ΞSӗ���*���d�I�Ę�M;p3Ԧ �ia�>R�3ғȤl���tȿ�Q�_oh��Z�ŌRU8���|`8���(@�^�c[�E!�F�G�Tbru��2\��cc�8�v��Y\�!7ò�_����rcV��U��ix;�����Tpqq�����-���)���yOPH�hjF?��?G�������]9��H��	
�ڱ����������z�*�T���pp����|<E��Ԩ�����:RN�'��b�&FF����cVKl�g��A-�Z�:�|�������$�K7}R�G�X��н�'9��ݿv����<����
�j�*�rYW*�����$�"/0�<���������4b�q:ܝ��r\���A-{����AG��M�y":������r�U�ʖy�)��j�vj���>�>$&��}��}��I�/Y=t����+&<n͎�2�mt��{1�uHҦJ�2�Z�ra�Κ�uӊ��߰�S{9@����u�V�1I�=F%+��\m	g��]&�vգs|~+�ܻ'���v���-�;����9�x�	3'�	ޱ,�/_��N�G�0��\�i�D��:�^_��~�cL*9r�B��`�EJo.��gZ����"�>�z~<Ѷ-�u���f�WD�����(�:���ʐ���>I"���-0<*t<w�l���3=*�E'��W��S:݂��c�;���ה���͑�qw�mع�	O�M,ֶ�ٜhH�P��Y�x};�~���G,��S�;�^UqZN���K���Ow��p�i�29�9�X*Q��%�=j�&w�Er^���n0ʢR�d_�0�V�$)d��3���0(���1=W�j�:b!0���>$kSG�B� �_O�h��Eg�$�f��+e�ڱS7�	����ñ��i.@
T6��۫����FNg�V��.j���)0i�`���N@>?�|��%c�����)n���,��z�������j2%�qޘ[~o������Ka�9p�U1G���iJ�1;��~n�ݱ���	�9Ǭ����޲��4b.���EEE�{E��&��,ٗI���Ƕ�����,G+of���i�o��J)����G��>���&ȹ���6S�7n/�Q����c��t.]�C$�}�S�D)�耀���!���r�칋����Y���f�x6x�2++�$s"޿ם*!eQ���'�/̝ �N����o���< O%�`Ri^BV���Mk6'V����$+����pS�D�;d[��`x �����<�+�f� F�Wy]�����ɝ�U���ɾ��2#�8�+�MK��~�p�Х!���GH������M� ����M���fY'Ê���&�}?��6-;[�����.��PR��e5�ع����̹� �)={��)va}���q�`�_���X2����5��d>�%L�`����cQhh#��[�F767��(�������Q4Ȉ�Ԑ�9�� ���K�����~s�?JW[��I�`��:]ش�	ȥ%&V��z^�H��H��h#rmx��y]�(�Ә��VB0�*�ر���6��N~��:A�����@6;�k ��G&ʷK�"
��tﴰw�ܟ�Q��`?^���E���"�4��*^n�|'ѵx�t���L�N�������������gN`�1��k�W\)66������*�r��/k�it���H����=5�_�ߟ1�1j4וi����H|������'��ƙsrd�7Q�Z���&-%�1(YW'�8]q�4�^#�)@l6C���T�!#c���6���#���N3�mII�E����R��c5�39���m:����y��H�7@Z�@� �Л]���?���20¯hIc�T�1(� >��#���{Gm�Gv�x�v�}{�p'�b�J��'�n�d�JB��C�Hp��X^���LMKc���}$�����_��8�5����?���+Wrw����ҐR(�T��|�RI������hx�y����� ���R"�[C������r���[Ԁ<����TI�t�	(�@s|���=Dqv�����ǉ�?A#��(ݿf��X|���!�� I�]�I�SXs�?��S�e	��"K.�)�N �v���Q��FHS]QԨқЛ��K 'o�@�n#��ebjJr�C��ų����Yu4�Xm
�UJ ��&R'��nkg�� B��
,![��wf����e�b�z�|�|}5<��
_��+pt���a����%���������u�rE.\�xOnyU`,�G�����E�N[[ۗ��<W;��68E�$�Zߵ��F����jlm�_���i�d�nм(5?��.�s��0�{c�S=�c��;� 1 o����%��_��Ҋ��u�%��;W��x�B�e�{o�S���wX��@T�T���PI��+7�KMMM����&��\�@8j��ZΫ���vĵ���C�]�k��@�iV�X�˖Z^�������񨋰���w��Q�+���j�������E�Ͱ�ߒ���e����r������ƣg�׬0	Y�)�P���]�{���§5QKI�����{�Unn�v��N�⛓A�����YY����oO�\�Y���b'�r^kH����ic��H�tk))>_��~���P���4�L�?�CHf��6e��~���P��`�lII	HJ?��ץſ߅��T��D��G�J _��A�-���'������r8H^��%���Ḙ���0��_f���=}}�׏w�Wh�gFTT0Z5�k�-N#�R��������ư�O��1d�������rL�S,�l�#Ժ�Y����~r�����V�ٰF���@�SW)����N�b�ן� < YNZZ:��iQ*����x�����ίr��W���*����q�����]7��CB"�����^��x%�w�|��~e$s�Y�$c{�����ͨ�5����"�������y0�Wy�W<#zRi7z�!j*Y��2��U�	)͚2��X�nSYsS�p�g�+�N{w�p�5�>ug@^U5����%����3�Q�sll6���@`���Au�
eۙV�MGH'4�@'����h����1�< j�n\��x ��U�k��7��.rZ�\���ߝrZk�UH�I��Lbk��y��nQR��wt��h���w����a*��G~�ü9��t!��,�ä�N}�=�K�k��9���[B��'�x͛�M{1j����I�nf�e��
�d�i�A*�~�83f}k�r���B��-##����`Ձ*]W��g��F-6y�SeS-p;r�g������������7��,�@3u�֧`歡ڮ�lX~E��fg��DW�:Wpp�qw��Y"�R�@*&��4�Xq���׋W�)) ������:��F��h��@��ş&�Jۭ|+�������W���^Ul��^U:�ܾ}����V`paJ��`��U��G&��������Z��Y�uK�D�Va3�u��*�A%@gh�J!>$/|m�ߦl�ݻPh�R��j���ω����G���₱�BG���£dt�u�/SL��JTk�#���F++�gW6њn-�����JɟR�[���_����7��0�N��hke��O��(����c����`�
�d!/\��q���*G�N���,�ɶ����á{X�YBe(�en'�b�r�G�~�ص���O���8E]�J7o�i*�坙��rۈ-l6m���2��X��j�6h0��
]��ơ�ׯv�<�r�Ogn/�s��I�U�w]�8��.Gغ˥��κI;�YZk2�u}Ѐr>$�I)�r�q%̴�<�6�V��+7��,�7,�)�-qڨu�y8���P�ۖj�˄��4p�;8=}��)���P�4�Hι�JwV0]�N���8� i��I�	�����}/�Z__I�=^�S~�7�� �q��ܲk��[Z���?x�-��KVcOVko P��i��s?k�M�i-,������D��W��>���S�b�(i�?�`��x��@]�!pŪS������x��m�P�KNMMA��&�VƙW�d���;�qoV�46؍GT�Ȃ~����Qd1�yhZב��7��w�gW����v&I�����lG���.��$�B��/V�kN�5�<����T��}a̫��yM��S~�cG�u,6����7�B�qη${(���s�t�;�>w�����-J,�@%x�E�p4MSH��=Y~�8�]S�5`*-��2(s/YY����K�y�*3�[G��n0�:��d�0=#��ȒM�4�D;=�?��߷�ݍ
̟�aV/8���Ed�E�$e����1PdZQH�gE�z��x�{En�\{�陥F����h����R���Z��S@��f�����j
����fG[����#?��1B<���aǂ���Ҫqm�%��?�ini�}���4𛣃��A�!�%()@� ��_����:(�Ay��4�K�û�Hh����-�o��#Zyff�^�l��Y�8bÔ��o��؛��}T�D]e]��J��ѥ���+��4L8rz�	���ICWY���Z�Lidd�v���, ܤ�e�-����]���K�*31���U�[-��:d���#��inR�u�Kr�ʹ; esp��m'H�w$�M��.�U�n��%$�8=_�n�*��_����G�L��Q��_�j���v�p�|G���!��>D�x���G������W^�������tK$ @&�'��؝M�(�j��r�J���B��L����("ⶦ����|�{�S��w���_y惜��߾�A�!�|-���n�Z�xǔ��ŗ�;_���&!%��海��Z(���AX�t���!��O��,�����-�bŝq��_h��C�x-Н���PD,�b��zlU��l�Pp?NBH����=r ���V>�
�vO�Z�A3����Cb���o�Y�Ƶ�̅���-���x��h��)wc�4�ab5����K NA��r�����e<t�F�v��^E%bc�ΰ�I�<�}{�X�aH��d��Ǵ��@e��x�%s݁m��o���֓��2��6���Ol�L����[��z'��)|�Z'o,���:=�tAN%�ģ��qzR҃$��NcK��l�Q<��8���OI�c�4Z%��p����q45��Rt�vt(���ެ��Ȼ� �~x�5�G&����QN�`�qP&�5�
~ � ���3`�����H������z��?�P �;��Ͼ��pƭp���HͿ&Ѽ�ۂ������{F\���zG&|#�m�[�~�#���a����و�����7_%|��1���� �s,��2Ɋ�1��c�a��� �vAۢZ��~ �o��S[>��9��vT�z�?���W�f����~���Y��ny��b��D��t#<��@e�Ș��t��Ky����&����� f�~�^EY�D���G�\�[��I��*���2u��TwFF\��3_<�G[tG8;�D��U���
��wO u#!&���9�Y��`���� -�?���:,�n�4К�
��P��( ����3�	�џ�/�aBn�Zn8D'K�> ;P̑��Ǒ�륹��w���w�
uS��ux���
���:.���EI	E)EzP���V��nPI��K��[���r�`�������������|��C?zf朽�^�Yϳ�:{���5��s�����%���:W�r/��MZ�mѽzT\�]�4K{Q�8��5/��c0�ԗ(��sЫ/׵�r�fr�%v�F��b��{>��硷x$�o�IJ���V�X���t|� ~=�0l��L�D�p���zg3 ��*L�����>��pȂ�ٵ0����<]��	.��ƃ��}w#h(�����Ky"�M��&=\T�5��4��U|�f�f�E{>=m��7�I��.H�l~�ɯ�~�@y�����Oe���%���.���?h2�yTB��{��'��W�-H�O�J��/��� i���gR��3n����R�?~[��u�꠴ W�����L��J��̓��zо~�������{S�QF���$��}F,��1��k������8攗�}h&����3gk�rku��Ȫ���F�`��3������Z��G(K([{��hy)=�3:ﴇ�i6�'N������lv�]��*��ý�(m*��3�R�^��>@�`�ƀ�S"����B�	��+;���Ta��T3'��r]җP�WP'�����'�T�z>��T$�ƺ&U3Y�;&�G=,4��h�J��k��#�5����>�b[cES�4>h����]�!��O�>m��W�������y+�1�a"YD|�����!� �|� 8w^-���p:X���3�^��-�{�X�Q4E������P�B�%	dSe6� �����#�p��#}�M��B�l��m�R��
����%xR��ۃynFFF���s\~)��8�L$��Ohe|^��ڶ0y�V��N�x�;şq��8��WOO��NbA��D���/�HS��I����E���*�w��qa�&:{�P�^۸��tC�5�L�{I�D�r��׼�߳ �! :ͦ�L��QŲ\��Un1z��Mƣ##����Z��q�>'nG�8��y;�Q����ej]�˫�J������^X;�?�#}M�cwd�����p��L��pYy�UBLTT氂�<=Pmuז���'����:'���ӈ7��ޡ-�T�c� mC�i)�?����pG*��G��ӧ�L��"͆&7w���[���O�E��
��j'��a<�� h�0U|19��$�}�xS��.LL�D'C^��7���z���j
L���qu���|��
I�^�xR�=K7R����>������-O
90���m��i]į�m�=�g�MʊB����6��G���vww{I%�A+�4J��%�6ǧq�?�IING݀=@�9KJZ���8�­Rد_�X�}Rg'��:�PR�K[0�`��WL`�qʺ^8t��X�a�q��������{�3�É=��O�/��:�u�q��G��+'�q�=.���1��G:�W齫`t��_4N�HV6�:aET�����I�����j�L*^��V��ؖ:���ӏI�h0�g-f�~U��3`�}Ij5���;���]�%���*�,��VI���3��a�YeTU���S���cb2�ݨj�ǲtT"�Aj�V���ܘ�{����ƪ��(�T9J$�u&"bja8�42jq����?fM�D^��覜�%HGZ������}�K���I��5L<x}�V�å��.]�G�:��1(�W��Y��)<t��7�8�4��V.rVY-೘o��^�(�[3�^�;|�"1�錠J�]�RU6B��/p�r�A�_�c�{��3$�ʍ�I ���	�~�]�}	x|����4/�׷������΁|�k�?Qc�J���\�b����gG����ޫ)�����p�ذ3�%����qgF'#��0�$9��kd��>�O`�K��
�L��HrU#��^y�]��4����O���֖�����z�h�	XyY�ؘ[�du�NB�F���ɹ�*����[�z�˺�kLó�1���ڼ:8����*��i^s|�͔N���z@!����HXR����U���OXt�:^_��6k� �@,y�w����s��sk���^Y��2���j�N��\-�����n�Qt���C��kZkq�(>�?K�Z�n�jq�Kn����l��������?�9�^o�����%������9�p����%O��z1v�'�7�v���M�9������O.Cg����[�P�sa_)/�%���q��V���d�u��ͳt�����D`����O��k�PG��JJ[�V��)>J3���v�i�R=��l|tg�e��[�3Cpiι���'A����W�z�l�!{^�y�r��q`>����d�]8�39I���so�˯Usv�R�Z7]�d�[��2:��ߊ�|�	�h� ��'�3=�ȗjr��q����;f6'���Vƿ��W��!}E{�'��Bt[�׻�N�X����� 4��}u��$TI-�z�?�}:��w��ȁk#����a����T?���V:��4�j�b��.�24����'�	r��a0��)����X�J�g>����-M'\��6�Ȼ��|熿��΢�Q���f��#iY޿���-���X?�gs)����ép�B�j�)�u�n4b4Fq���kA�T��t���f+�%��U�of��`i̤���p�᪉ԗ�����ٖ�|���J|��m`�=}�x���+L���K�e���^����E��L^z8{�M5�.y:u��}�H:c�x���&I���ʜ֣P�w'3rRBy_��=a�\�t�;3l7��Iҩ�B�H6�*%)���A�!�I�o��u�w�V��h�[ux��������bTt�,IA�Oc����Y��;�//����?T���qW)Y~f�8f9$[�0�l����7 ��$,w�>Ǎ�f�D�Չ�l@�s�"UTU=U�E���M��{g�Lټ/����g�bG�)g-�~�?ռ�U��E$�++о�� U!��4vR�-D_Y*-
@�...D�i�w�sDۃ!+��u�C�;w����~�%	�ٍZ���
�;�z*"�fhl�;*	�7���ej��0/m�.���V�+WY�Ʒ1�:o���.$��*���aL#Ͼׂ2��ڻ����L���o��bc�lj�h��+Y�9��M�髃�I�F�o�y��{���|��"$&���{����1�φ�N��;��I�FM%�b�����-f�A1�H��ϻ؉�PڼQ��Ҵ��q�V��&���j����7�8���_�)/_�����iQ�XY!����Կ�*���Ƀ� q���6Z���3,��4�&v�����O��v���J��H6�y�`�:Wi��$s�:O���ާ]��c�TUCąDw��5�����>R���+�!�н�ݼtDRFfSY7'�-�Vn?�����î��A6O�M^�F�PɘW���M<@���[?���	�y?�L�l� �͓�2����]�1�o�Cw�Ň�՟��z��G����(E���>�ZrT��z	Ѭt��o$GG�-�����8����rYi�j��@'�i%�� !D.K��A9~U�3S3��7�n�n�[�z{�����K�J�n�=V�J,���ߍ�|oY��-7Q�J�x|L�c/5�(O�8���~.�0U�&7��E�2�*�<s���$���0�F>1�~M�Du%�	lC"*��	���Rv��ge�i;]��nt�)�C��	WX����
+{QOP
�v��-�$n��Y�S�*�^�k���9��s_7o����o��NsI��+|?�L����.����Y���Wn��W�D�r���-��~�?��2�~�W�q�?z���K0��Z�
�ʶ������c�Uo�QnB/����Z���}Np)��[��G�8j��x/��؞dO��nU �O�d���������z��w��\�� ���ͮVH�ؾ ��p~���m1�����<F��VTT��F*V�DO��d��[f�`�-z��<�t&+ѻ��v���0�cv���i���:WMuN-�	�>	�|PeEOP��ήT�d�pj��h����\}���1�NdБ8=�%��<��G(<�\{z��y��2�&1�U���X�W�r���	�z��Yz el�5� ���D�W}��(z��74��<Y����i�Q=�u>h�9��;MCI��t��C�R�b�X&�5)�[,�੹+RV��渦8o���q��7���U3�!���U����j��������|j��V ��HT�iZ�BU�a8�_��c�������p����;�ȼ��%���J���aEu�np��ޱ�-^0�r�^k�n���cq��SG77"n||�{�������;����S��S������*����&����{���-�f�:+Mg~d�:��S������(6X��r�YB�}t�Qo`���R͌o���F�0�<�xOoA�1�p�,�tI��s�0��w�ܱ��%�����[��M}�'���ͥ��'F����G�V� �@��۰3�c���KIS3�	3�/�꟤�	�²qX)�wם��W�C�smQ))^�qr������ ���x���g��&�}�&�c6�|H��(w�_�J\ow�F�(�z����k�(��.S�c�mu�p�^G���)#`	���o�&ѱa�U@��e�v��w[�zݞ��|E��m�W>��'���58X?`���|�����FnQ�U/��.~�f1�����\� ��F��bf����וj���`�i�Teg'W��K�J�����	p���5��g[>��Y@����Z�N쇯E� "��r�S���֧nn���Y�|��w�j�
���J�a ���o���U��������~���Ĕ2.Ϻ^Uaf�"n��;��",K��:?hEk|e�}�6�����I��w�˛�2U9��[����UX�T�0��hUY�U���~����%'<�82*���G���+<�O��CLM/�wBV���*�ף�p��y����b��Ć���A���y�iz���wI��սCz�T�P�74/X@���_�ȦԧO�h5��a�-�[*��X-�Q׾���i鲐�*��_�Rc��/UU��ہU���]ՇL�u���=<[O��Ii��P��A%i�`�ܖ�����p���2����脝���2K������tmjSU1�q͍����>y��f����l��3�[�.�q��GW/|`�K�~?����Տ��9�	.qa?���ٷ��Z���Jˠ���w�КG�wn��+i�vy���I�WT$@w�����R���pZt�ŧ�Q+�(Q]�.��c��)��u��V��u��ۓ�����\��eeY�J�ԣ)����o5W�%���O>�`G:�J�xg>�ŇxY�m����©������٦��d�]�k5�!TY�9kEHL�}����n�e����+�L3**}�Z�A`�҇r�<�^�p����U�$����}�;���;z*fTv�T���� /Tkn��-��9O�{��]�_pǴ��s�կ��U�&�i5� ۫n5bbQ�Fvq�_8���rU�t�,��~�^�L�#ү�pٿ�:CG�jc(���¬�~t�h>V�￟Ҍp!���p#EI���ښ�zn���1�
��y�OEU�8��&{q�D�4��M�����x����}��E����j)�k��wNH���AZ?-�֎����$µQ��Ȉnw�V�`uuU-I=����m�֞I��Ɠ�����j�(�����P�[Ɔ����q���nh�{{{}���2""�ߤ���%�j�3E�����wQ�wG��÷wJk��.�x����^�@~n��^���w��df��ee��M�܅���MQ�ΞE{���k�����9M^�<4*"�%���+��F9oL禥1y����sI��Z�i{'���v. $���}|x_@@���6�dg'#-Mʙ y�L��@%VU>�gf_��;��(��:.��zypp��D�����e���b
����_�@#��G��� e�?r��O��?�]goF'&�����#��SQ��x�jWz�{��f�|~<���R��ڄ_���ܜ����Z7Mw��дo�N�I�P+ҙX�)�=��m�9����{v߉�uGf'��죉������QuG�z������ǌ���i=h>*�3��һ�<����*�N>���jڟ��g��N�[X�ҳݸ�	�A�ŋ�;�i@�i@dOC9[��}{�͑C�/����)�i��u�7q�N�#�&��&Iv��B�9EEU�����B�Ӄn/� ����(��[<�I0'���f���������������C��1T�j^~0�B� --튃#9S��]`��9dZ�Q�U'f�'DF�M0�O����_`+8=_���4�_�d~�,%V���.B$u���-��ۯ��M���W2/��o����C�\�*)JlkcVV�*��gisم�$,����!�io�E���V����z�	c"��[�q�N�2�� �7���R���kk�c��e�CZ+$�cj=����h9�P��ust��Q�}آUe���X8u!P:��k����q�ޥ�ꀔV���7~]�ٹjk��gD��+��r��m����ܼ����>f�.}��^h�B����2@?�z#C�$�
Z��T�߿<�Z(��K��/@o�#�E�ҽ�����j����F�c��C!ڰ�ԍ0�"��|K}51-4�p��5#�9k�-/]���ch���v)��KNP��
�9}�d!��N��s���R�׃A?���t�0rX��G@5+�ܢ�:&q~o�iv�ꠤ9�^���.d���m���n� ����@+����/_�.�(e����-Cz`k�x�Z��	�w���}*�_+u�4Y�5{��_T�7T-.w�=Jy��T̙~���
0�D���mn«�疔��i܉��I2l��:/���:�O�*�W =q�N�#ݎ���Ғ��=����ٟ^p���l�r�ULսd�x.ݺ�P�`�-ˤ�/_RO�O�I��>`�lz�3��
듕�Sn᥆]�К��C�N��4��෧P#��I )CQ�衴agH)����z�]�@��0��36܈��
��Էz.]�!���S�=b�N��̲!�W�O�j�y+]��f�FoX�u�� ]���M�FA�N�����
��᡻�۷9�]a�3��Wi�ޖ~��o�+Au~�OZ���B��T�n9k5U�ɅS"��Ʃ[�BΪ0O�q�_�+;���:�N�b�r���~���T��{��jUUU��������I�ѱ16 ��1 N��W��һ/3^ ~��PO���UR3ȇHp�3�Z��������
�`F3e)�2���^5/�Q�V���C�S<
�l��>%�VD'�$�ynu���Ԅ0{��0���]UY9`S�JZ9����>��6��{��'�@G�q/��&Pp�\�-��'�74�TVV�Ң��F�{�]6
\P^���� �z�d0_v�5ֆJh����C���F��`����F/���ݝ�P�����";_����e�v�[��@az���s��жī,�C Z|���M�d���?�ߠYn�[S��"w~WXX���Lc��V;y����*���J�l�m�Pw6f���=
��J

���= ����w���(+))�,��0?9]�q�TQ=������|vv����E�<���L�$^_�qQ�}FB����v������w����W��^:#��(!�,F�����n\��[��t�?��=2���m�gn�	�[1�ݻ;�����f}�FXX�2T%����ۈ�o�*�k�L��_�:J�d�t0>;�3�Sե�-QM�-�k9%C���+g}S/�kЧ��K�9��ז.]��=�$\�zgN�뗰VV�t��7��żu���ro i��j��_�� ��q�O�����{v;wR���������>�w�^�Kûw LbaNlX��k�璄](��0v>߬�	)�
2��>|��-z:��.��^�DP{2�ל�yz6(����%Q�{r���ݼys��./���n$�}�1� ���qr��^+t��U���Â9d�z�q���n,�q"�ς���}�ǝ,��"�����|�)x<�(F����R�X|�����p�D��Q��1m�\����/m�w@��=�|�(�&v�� ��(���?Z�F�t���ՅS�l����
� �����@L�P�����b���n�(#��\�\�=��ϵ0�(/��KɅ+%��!�PX�㑜[J�	�%�---5���Lu�CL�p:
�N!3������;
51QQ�`�����㠋�ML�6��������o�V,E�r���5�T�?�:�2-++�	R�Ӯ���K_"m/�z��S�W��˝1�p�q8�XѰ��/����j��J�λ�[����R�j��x�(��|��L]G�c��I>��;�ћa�T�	�Vccc�a�w#K3ec� 2"k�lP
���钡g^v��|+�s�����f�1��`d|�����!��BF� |�?L ^`E�իVZ:��J��,�9�̴k��i)އ���j��#��I�&!��Dn�)4w�s��;G��h�|�C�R}(�>ڡ��#��e%�[=��Ҋ5<��ݑ�NUE�2@�G�.Z�l@Q�J��9���c���,=/�p �B�������8�}@'.,ۗ�TW`#�X�bc�Ԕ�ۄ����1��y�:�s�>��y�DX��T�Ք+�~we;����zt||�0*�35�����јQs������,��P'��N�r�x"���Tt��or���)�E���Å���.�tR%�xT)4}�;��]��J~���_K�<O�������J��E���sp*C@����[�^��^.��7�2|�_-�g��U���/�Ӵ�.�-/��-�ؙcz1_-r
�J~}�xh���Ү����Z�N�Mz��8 �%3 õ+��[�;
v^��i���ZZ�n�<�Gr.!����w���>v¡�ҥH�{��?��i�U��L�Id�~zδ�s�;�i��x�hzF�KF�]x�`1��q<\\$N����v�B�}��m���bb)�I��߿?9'��b���h΅�9�r�����4m�h4t�j"0
BR�p�P(��⣹t?�{��8��)�¿e�s�N/<$�䰫�7;W~-�&e����Ƶwt���̑z�Љ�y���6���i��BW8戠>�]=���@�Y�E|oc�F���/ �^��^�>y�k�3����Kkk!��+k� ;��5�,o�+��Ћ�;\�,1�+� �\:��p�spwv4�a�&��$��F��*����t}#C�s*br
r&c���(�gw�^�I\m<��4�Y�rK����:��o2>wIKO�FC��f�?Ho�HC(�@I.[�-
:���Z��R�B���U(��Ʉ���),\l��U�ɶQ�%�ٖ��hAj���R@-�'8�{;	;�fgf�x%O+h�G�_��xupl� ,~�V0P	���={���ag}��͛7� ]?|�z���0J55{�^�W��.���k�.���
�rw�O�����s� ���^6jt�R�E�r(M�
�G
�Z���;'����f�x�%�$�ݵ	° 2�����}k��d�67��޳��˃����30�S�T8=�VQ�~(å�
�@����3hJ�.F���U�����<r�Z\Qq������;7n�ON�5��p��z����������+��^�ʇ����Awp���@��!o�Q��:��w)o�x}�k�=	�2�ݐ`澷q5NN��zP�-/ﲀ�g���b&��"7�W[֝���E�#i���]�Xv�|�1`�����E�����@{2<�#K�ut������g��}]Z�]MBJH�RM- �tH��46��[mu��e�`]u���g;W������>	���>��\��{g������&Al{}�^�����Axy�v��{����=;����J��l*!{�ݵ�P��R1Z���A鱷1j��3YnBZ�S���Hq�w�1�������U�;���|⌬,�JcE<����f��CWWW��{�����'��lJ�v_o 7��ۣ �[ �'>v{� w�������)�B�m����%��p����)�|�m7��<�|o<uӳ�d�?b���P��˄RW���n���ږ�,��YP`��I����j����P:�.��c�6��!�A!p�ZY�wg`}�#8снM�����*�z���l!J�''#\;pYW2�	�!���`j"��pp��g287���H�҇Sb�
������'W��h0��c���&�����!wn������0X�`�2M8�pb)zq�������y$G�U��n�S�0ږHV��mmmm�[CU. �� ha�����>�QX�tm�n�$'7,�Cv���������##��q/w�3�9���`�h]u���ژ�i�Ǯ�˛�pw!E2��G���N��Kh�����ꈍ��.��p5�;`�-A&���җlQ������a 5nw�::n	R�}&$��>�`�(��B*��,�R�YK.%%e9UJ�s��ݽ9�!SW��1U�8�˟�\]ѯ4��C��u�L�����ăj?K�,#��|M���n��&W�~�,���[S�U�HJ*`��G���w���ed�ƺ�ks�)�M�y�t���)/5��0\|d$9<E,��F�JV���077�ô[+m��;���K�&ɉ� �8�L,�tj޵�?�[@gh�l�d&[�DЙ�S����x�K������XAi��]�D���g�!��w��llQ�-�
�Dj���W�o�8�n����o����372��_{��'�'S�/d�5εR���� @GW�*̔#���ԥ���⣢nB���̜K�izjiY�Z�璒���5�-߿|$g�333	\�&�z��I$AC�IE�@��c�b��]{jo�B;�<���9��L�H���Qa��RM�s���@3TA`��z���r����-Y��O.�%�[M���t�n�K��2Ԡ��Ρ*vZ�T5!���4?o���[[=�c�Џ�[7&���>����SH��flms
Pnmm�x���BoBm+����
x�ס�/�\�:riw}�0xn�K��o���hNmj�����]mJt��g��΀Y
d�{s��}�v��p:�:� ���68x��w��A:R+��@M�=!���_koT��U��fe�MJ1x�'2���zb$A�{zz�iC� S]��|���<� ӛ�f����O����F2��ׄS�]~�F���jH�o���Xҫ0=��3�!�&��,����p�>hu��p�
�b����7N��8����<�mC���	�2����a�қ�7�#��e'��]1�����H_�sb���
�\���C�z����4�8	�dn?������듣�9�0��z�ҕ)���,G����nZ����-��I1���"۲9K+���.6��<��"�$؄�O��?9 �"���3��o߲�$�n����7���~N@}Ǌz�l�.X�Op����F�i巖���4���! c�$3ܻR�s�p�FGG���Ы��v��j�p��9�h�

$E��a�xbfɐo��/��\0���Z1o��NZcb W�}N��r���ĊO��1cӵu�[@��J{���k��Ї��7c�
��H'��w	m���3_'A)_�n	�,6Y�Ďnq�ܰ���|R��x2��9�,��J��ģ���+��3濨�,s=X���#@4]/���Yn�][S�����c���_UW7�ǏWp����?�.j8O���W��Hy�O��ܞ��}q<D@��S?�`fb:���rRRh(� t���{7`a�d8�K.iQ�&|X���<�eP~"�!q�z�;��C�%��&&z�eo/���C}V������'G�p��]�@�R�ξ#��n@�1/{^�5鳘��&����a�)�	�c�r7�1�mS)�c�#--��$�4`���;�H:}ϭ?��K�1�������٨��4�H��Ųߙ�TJ�y�%���:d.�A�[ۇ�?#�"Sʫ�:�.5��1)��k+ �T�c�8uj�3����`.���ސlM:�&'���b�ܤ���4��8YRU����zN#�ux[LL�d{�r��Ȩ(��r` 	)��lL��M]�P׌
�Xx�}�34�k/#�;?7�D=}����� 0����3���-|���H��\1��jjj���������D�"(y�=y�Υ���C�vέ�|e�(�mH��mi9��y&"2R��<���f�)g�ŵH�%�],�D5%ᴀl+}�r�b��G�vR8 ����(w�9�������NAM��!���W~6}� 	�Q�bw��I��@ �P@�z��z���G��W(�ځm�66�9@��2黝��I$k=�M�q��;������CCנL�#S�ngu�nL���KH���A_X~
6�7�&M��Y�J��X�s�k��������!���}D�O�ѻ��ŵ���:��Xe���@n5Y�m�<�c�M8���1z�%A�]ˤ���[�ΖI�Y5���.Xd�I�W�S_��K@�tDܑ�]껕3j^ع:�z��`���͍o���g���АR��S(6��ŋ���.�\��ѬB�|��)P��ss����k`�6�П$L	������'A��ЩY��|�D�����S�1f��'��Skk�%xR��|��Y�vL��/����a�|;+��ٙF��o\.�,'|�;�]�VXB��J��8��oXi� ��j����[*���r�TT���$����Α��@d
�1��P2����<�t�L�P��=J�փ	�#3�|�� ^�-Jb�� pT���r ~�:<L8t身 ����H6��}%~r��K?'{��A�G�,�s r*�3�SD�H��ymY:A�0掎�'��fjA�����ٵ��>�_l��T��(=�f���k�iNR�����o�*,�/..�d�l�tT��B����|��U��V�qsr����䢨��ԍ�/tS��}����l#`�߁Y%%	�m�! Ͷ�����sj��ث��n %��M�s/���
_?/�>90aaeE�8
��>`zG��p6�t��1�����5�8^`��	�"�"N�*�V`�����i��5GG?�B���x�H��x�>%��2kܶ�X���h>���Ϊ�HR�.X=$6)�ս�ew�|2篵r23�;=��s���������J���Γ� ��8����n������EU�����!�����M�`���
^�k�%J��x�K�9n�q3xY�6'�xP &ܑ&�	\����A���t�+��!)*~�X�/�/��� �u!=\��Y�Lfk�5�H�#¨�>��7��8 �+n>����3� \�����Ic��*?D� ���9�&O/|�΅�_Ǌ�p��:�`o��5dc=��_�= rq3u�Y�4�Go��ɼ�*���A�A�3F'�Kz����h��yd+U[�U۵qn�Ǯ%�H�׆���S�a����X������S+lP�� R�Y���o [��D�TTn��
�~�ҙ]SC�@h���fm�<��Joo>2;�"��ʫ މ��|!r�QQsl��ZZ�8���9��($���/_�uϾ'��`i�KKz9�zpwm�M3�kU�ɺ������\eV�w�F:����������xر���x2j���&�lF�[qy���
�			%"h&G�q��I <�|��O�l�?�o�����(sX"����2]���u(i
iΛ_����$�.�Oج�N�rѫo��7wu=K>a���q�A��j��*+�٠���
�j]>?�mg� �i<����n�P��.�r���L�����g��I�vi
b��I��!���&&��� �uݛqٚ0Iy�n-v��p+/+�,�9�=���Dq)100<��W��
��� ����I=�x�ʂx�Iju�KO~�4�B�B\��#�R�C�b�}�f���� zT�F�+w��*��tm�HF�\ê�������Q{����-k�*�$�[��g޽��k7v���Q�^C1e�N@�_�Wn�ip5e<75��&|&�)��^n�\1���g�f�dH��_}�
6��(�0c0�b����ߎ�CI�"��{Fy�mt ЅfO�H���}���j�-'�vj$y������mt�y�֭D�]����}j��;@9~���J<���
�ӠmF�,,- 2'b��7���T�y��.�����^N��8���ps[��v��ū<�����E�N�+���	�f9�[!n���8��K�AW
9,Q	R/�v� ��*))��׫��~���Cp54��YӋ�" �~r��G�9�D;:.�M'�~��{hq�~�7b����t=4_�>���9�p�7'�&vGb�
� �KI�MَyD���t�/@;=1A?Ή<���}�BA3QI���fE���,�h�RVns{b�����a"��^r���L�1%�99�~wո�����(��������(��:ill�dedʂF�xս�EM܊�w��k{�,'+^�ح������1}��ť��!���wc����u 4��C��A�
��Ǩҥ�%]]ѕ��[_ۑ����� Hۺ��d�1u(!d��H�	T��K#kS�=����ϝ�@xW��ى*�����#���J�$;�-�b��.1ec�|v��w�7ơ���������u���?v�N89A�n����7h��w� �s N�X���^(�5ve]�ua�ggT}fL�9;?�*����$��&~ � c�v��O�"Ê&����� e.�g�@.������˗d�~zp�l��y�.�Ş�*���+��n4�9v�P@�?P� �+��p/�h�*�B�c,�T<Q��j��C�R
X.�MR9 ����'���u;��)�54���霔������|�]��K�3��BD��K77!��9"?W&=L���^�?$�n:���O=�i�F+�:�@C���b�|�H��o��P��zlS�o��ɼN�o�N&0aO@�Պt.���1�ќ�Yg�gffn5ċz�!�k�;
tj#p}����n�ڪ���1v�In=�+?�=!�L�4r��ֶ�k���٤�?^���bߡO���1!���LAM��&���b� ��s�c�gr�H�ڨ�&\�(�Sa����DD��/Y�;cFQZ<c�ׯ����ڨ��+[=m ���ke3_!�����z���
4Z�8��.�N��0x�I* �Ez��s��v�1k��T���"���ВJ��h͒�g���联.h���8��B���Y�y�k)����Ǵ�Ra�Tۨ��}7�LT����	���aʃ&��@'����C���W"��a��A���!��Z< �D�H�S�R*�� � daRx1���[,�a��^�|�B�Ց�ϥ���@uAt~6�"����ʏzzzN=݀U��p�p��+B*g߁DM�n�:xmu�)�t�R��C��bnnn"B2����Tu��d]��I�Gg��2�Bw_O ��E�E�/Z���:����h b������`N���(��c�.h��"���t���P����s�X�4WE=	r��l˹�~��\����4h�{m�K��;pA��m�$���*��X>��Z*�5�S��@^$hU�d�2�Ł��Y1�ߋ����fʍ��ZZ�	ߜ%���?Y�nd�}嬒��vBD6T�ز��r���v,j5^�:�Y>I#b��yM����Ŵ���Z� ��������Z|����K�Ƨ&���C��kjj��CS[Q11�[�@�:Vh����ܚ�ZD�E]���7ۦ���/���s9v=��� ���}(�k9��]�Aw�0���+�@Ȼv5���^!%�q^���^���\�a�8����x�dT��Y@��_g���EzĠ��'�1�Z��+��E.��d��-�ݽ,���5�?p�X��f
����y�w�qд�������g�g�����<�����\raee���E	�Ё����!�U7<Ydj��3ƹ?���v!z��/�+��X0�Ty���ar�&@�Ƣ��r����Y��^;7����"/\��x"J&OyɅ�zc�sДX��l+A���/�`ýd��&nv�O
��7)(����=�VL���VX�s�G�utH`J
�>�As5���c�O��>V��|$$�	p?$��� +�F��,D��ʪ�
p7�\�Pze����\$woO���1���BCgGǷ ���bA�.����"N�䶤{'�x�ChG�j*��s$�B��ӐbAJ�P���r�:@�,G�45���EzNv��Kkj�p�,��,��8i !�֘A�@�μ������&"~vg�t� ��.�����j�����-Y��}�?�����Q�����2\K�i�v�N͗_t}���~ ����p390 WE/����\��&�K5���⢢Fm�Y�_ZY��`H񾦃�B������?�1>N4��E}++{T������w�h�L����5�"z�p�M�ְ���]>0}͡�"�###�௒�@�r@u�mll���^^/"�?��R�����454bǶ����ը�yB%���Bm��T��Ui������߇@� ���jH'U�acww�H��W���)A�F����a��[���p�j�ҙ�\:/S��.���o�I����S�S�b'��o|����O�������N�� �����{�.�xH^���E�;� �UR�_ߐɌ x�X￤ȕ�����$+2e����������t �8�	�8[]�D�NNN醨;fО�ɠi��S#�ʕ�_#�����:X;�Z��1<Ls|xt�9��n5uxjVUM�?V,�im��a?��->V�lBKvV�y�����K.���Zؽ��#9Jx/ ���~vs���a?8�\J/�O���X��OO7�e��K�����c���н3�>���=o�V��ca_�H�INA��|M���y��5FƧ�R@@����֦��%�8��෱���䚦���;{{�'�HSD����p��ēu���5&&$o�/_�:��=ӣ� ��ɕd�r�-E��!^S�U�8 �<>� ��ecz�S�9%Ŧc�������|���=��
gX��u �����)-�^� �{�����㻠]X��l�k�̟�T}��V�����,�(~�ǔ�����E�Ra�Ф��B�ت�Q|<��nVST���qjm����;x�0�Gs��ƞ�MWYMA4@��Y�Ɓ�� aG��<���F�q��nF�g�w0�$�d��Bs棗ec�$����E99߁�̔�tČ]�BL�� �\�]����:�����Z�4s�.(/J`H�@��	!�����������B��Ie�MU�67�_d{Pa�%����wwwww� ����=���%���f����ݪT�h^���9��~��~dl,Bn�����'�&�5,lf����n-� `K##!�|�"��6q@��bcG z�DU4����, ��o/�g+������P|�gO��wD�55O���W^ǁiA�Ύt�x�j*G�ְ��rg����^_t"L�$����@)n^��vϿC���Wµ��������������!N����=b�@7��\�M%ees�6{�1�h��@ȋ� llL"N�R4,ȟ,6�:�-A^w@�F)�x,LO׮�� �y�:�wB%TY99]�h�����v�ԸjY$43euUw꾈����U��%�"���5�9��TlfsTYz��	gJ����x�KQ�:.�+P�}\�1�Z����������
����|^"P���p��y��目���ܟ_z&ΧK�z�@��|^�_H��͹���9��~vFoo�y�=�&�%�/Y?Ujk+*z�𹜏fHj׃,�u"���Ҫ�8m��}���Ncjj�}qQ���Ȏ���SNiuE'B`�m�QDaHVVW
�&\Nn���S��0VQg'�7�D�~�@��%�euu	���mB#xyu�oqK�����ϊhhh�]]� ɍ/ZycF�BAA	�~zy���$zxxH�-�a`����
��Z���t��]?��a���ass���1�p�@���� J]6l&������JL00�OW���i0������=���0��H � �\�̂ȩܕ�r?����fA+w���@p ����
!�7��������{ ��������$ۆ�?/����� M��:���K5
�5cQn�\U]k)�P5�����.)!
�-��$�$XQ�%5�c���Hq�P2%h4{_��uW��ٖ/, <���/�Wܠ*̔!Z�
h\�6�0���Ly� }����6Ѹ�J���?x�y�%��L!��p�O3?+%-(�{�F�Ui�T�����E��m�8D#�"u���M�`�l��ki�z���L.�:2=8�7���¶��U����ą4��E�r���%�N���[`��u���ޙ���ɂri��u��LN}p���C�kG�-��\�������EF�|�Ӹ��,5]��H�!I�!���q}���R�j��Q<RK]��pA��N@�R�, ��0�4F�i�ο���|ג'��4ԩJu~=�7 n^���I�(@������X%��I�����7Krd�I\���W<��5'�l��ċ+�hKl��JS2Uw�����E��L@\�^6��Yg%ld�9HR̎e�ߎr�㎨or�hqqzZ�{v������������Q����v��NӸ�x���e����Z���T��T�=�����j$4�A*Խ�4�
92B'��Iz'�?���?2�� �8�4ٙ�i�� C�;Iz#.����٥��T]��R����4����6��w��m�0s/�y�NN�[�M�S��,#e�H��*Efgk��4h�FR�8��ɖSˡJI�-15'�xO}= 3�Σy��`za��� �NR9�ZwY���w�n�Q@@���!ֱ���&�+.��/	�~o��յk�c�������u�=��/�5	e�$��ݝ����m� ��U�c���}�������O?-����ޜ^ֵ��uqq|���+�9)+fԣj�7<Gnb�P!�Ɉ��R�0�7A�^#�}8���WG2�h)j.ob�>Ɍ��#�hM�vaW3�@(�)���Xi�V���vW'#����G�7PUP?�I�	yum��K+80	LI�v��w=�Tش�ʇ�3I��T�>�❕~�Ae�Qu�CC��~��P���*srx��{�(�D?C����Κ^�>}Lẖ�%[k���B
����J��&:)5':�Cə�4Lv-	��]/ ڧ������RewEB	5Z��z.�1@]��|!c�A�W�Gh���$đOyhꖚ�LrC�1Q#�E��{~��Q�	c	CL̪1x	�۲��2��_��|�s�I��曽��G!��!��%e%�/]�=�gF�%0�'C���^$���c_����3��l�����Ұ\^I�|9w��0�-IK�)ف�(&Z�O#��P^(��:8���.=���v�7A����IF<���`N�F��^���t���h]7�9ð�q�i������䊡�n�����ƒ�� Z1o�W=V\t�58���� �A�>��(J�+����,����SN�&I:�3u��;��/
��%����a������\]��jfJ�X�Ð��!)�x`˦�f&��)�bfI��YsEg��-�<� H�^
1^��c����Rha�ޝ�+o�.瞭��2�8 21С���T�ǫ 1�b �G�=�B�� 
tc5�%ҷ1�~�hl�����-&�8x؈[�C1e� q]��:���D�ي��y�(
�㎈޴���2�|:ev&�
�<)'P�BT=T(����ߦ���?�(A���=#�1�~l�)�X
d��"2(�3�e�c��%��ҡ��x�~���a�StD�'�f;��3����ڶL�~�BcݎhP^Q�Y���J�C8B$V�
���\Q&ݫ�_��?"��kw��(|\����C�9KK��؁K���gq��z_}
���
�;�8�~�	'�FGh�?�X!3�6�CT$����a`;����l�/��+�?�p:Zn�zn����V�׳Mi'.�5\./Dּ��������N����`fɡ̏^�Y!a����,a��lZbf��S¨)�y[.g3 ��C�@F���X���6:�D��SG�fqx�r��@)��~G�Z�b��#���dc{�Z7��KB�+姧��
s-�~�q�m"ΪY>���W�J-7�"�߱����P�B�Gd�1��V���v~�K�aAʌ��������d�yg��������Ì
���'|]P����0-m���שݾ}
:7c�u�sVOs���kL^�.�؝�4��߇���<(1�Gs���b%�0�����f�?�\�~���:��\h�ꞇ7)`C�V���sY���;MqԀ)�ϣu�N�X����]I�f�������m��<!���tl@�hȷP������Ŕ��p���_�X��Ak䝹��<AO��NQ�ym9'ly����σ�������I����b�����"ib��De�[NO�Ė��V*��Q�j����*޿�alٖ���5���3R� ��fz+1�$k�a3��Ȭ'l\f��AV���E�t�iƟ���׿X=؄P�0k�2�?�T�tԎ�?l���b�&5Mh�YQ�@l��Hd/�1TuOERN�\�(���ע��Εh���ֻ4>��Q+m�]�c+�`��y窤�K(��20~���0�.�Q�#EJ^�8g�=6l
���Pӈ}t�ݹ�����f���iص�Yi׏�g~~d2�4�%������k�ZYSQF�l����T>�9�5NC_5�^Oeb���t��_ݙ�/p�i$���Pد�å��6�{���ћ��/.�f�1�]���Q
C
c�YՍ���B�``W ƊZ6�9��au��>S!�4�"]�LN\N��O��n2� ,�Q��y?P�m���)<�k>��^Oi�;���A�RB`FY
pkɿ>՟����?qi�C��a;�v|}b��yz�j���֥�5�����n�F�r�ܑ��<�] �&�Eմ��@/�F���f�!���j�������l)-�$�y�?*�Y�G)p8��_�Qx1��g����,΄��������gDP
�8e'�ƅ�mV�8��q�Pߥ��'�ұ�ɛ��}c!8s Z�Z�v?�,I;t�`/�a�,�9�V�#�䈓�����=�]ҍ�W�"E�S�w��T����K2����:K
,��I.�u��b�N>���������B��o��ǁO��d�㔿�f
��˫�z�ʩ���s���/N�,���4E#L� .	�DY^E��QR��cak�����f'o�P����i�u����K����=��r�eV���ul=�?VS��ğa7�t�ꎹk6�I�i�� 8_C��av����}2�uQWW��-��x2�y����Y�9�TQ��\z��B��ç��]F��tdFƭ)�ؓ��Ú������_�^TW��U- �_�R@x1���'WZԢ(a
Y�,��1@Q��Ӫ4 �&	Dﺮ�� ҊNT�	v�p}B�v$�n����)��~󍽠�^�����?g@��F�^�{��^i��������iт�JH��l�P�
e+C�����[�"aV��j1'�z��
H���8�	)��ۢ&]>�"wfi�&(;��Tr*^H	�lY%;�[X/SNS_	��el,���R8�sPjh�uyo��y���Y$���������L�40Brp��M5��Tx��A�.83ɇ|�/
h���%¢dO������B��������S6�]��!�S�I"�F�t(�fQ�E�[c@g�Gw<Z#r�3#S3d
�)ƫ�vU��i����^�~�����ęi�t�?�X�{C0x�b2�&K�F����P-����4��{{ڪ�?;C��}|	�(�3�t`�&�Dr�~���0�a��A2y�70�?����HZ�X���t�Ë4�ӚH )9r�(.���O��S�A���'�-� ��X]��Ur�%c;�1�qH�HY�G�lT|h�/sgN�:]o�� �ɀ�)Q��B�����hl�B��(���0�
[Y2��1�� T-�|�(6??G��8��iǝ%I��ݞ8�.�����:)����<��G��el���]�4�l펇�� �W`�"�Z��KA~n[{3qJ]�#�y�8�d�@?���C�:���m�K�(Cc)b��g
$*�y��<�}I4~)@0��9�u�<!K/��ͻ��%�$O@�5�(��5��P�P9@} ��P	�h��,zwzM����T���
Sq����s���"A�����m*Ol��\Ԝ�,'��	? ��M��H3� �I9���ҹkJ�!Ma:�-���1���%����/@�~	�M����>K��)2�������*� �`'\8@��G�.��3���V"8B8RI (�J�˷	�����	܉�J��g��i&0:q���0�+籁qR�ޑ'����:U�ySS�A�瓄�u�%�?��7�}�Y���i>�X1�+-��_�)��,!�%��bw�Tר�c�G��W����L�(s^���i	�˱l������0��?^�Ώ�R�HJ?e$�ࠤ�Q��h�	*�ߎ/�UiH�M�osS��fc�h۷C�h9�P�a{@?A~3�fv�����m��ȸ@"65_'ǡĲr�q�g���	 � 9 Kl��� ���͋������0z���k�; ;Y��w
��)t����'�L�-�g�'Ce��'d?@����tU��O4jG�0�x��s�Ί�.��K���)�K�&��ͬ�	��4�)<P�n
��q�d�D��#+��sfWi=:��-j�0D�q�/���# I�
���� �ͳ
G=�Lcn�6��Q�!��K��Y~s���D*B_�act��7�r���t!bMay�K7h��� ^��T��ה6�g���= �I�a����+��X�IhU`��.��Ю9Z�����L�' |����A��l	AA� �k��u��N��ɀ?�,�R<썈����[����3D�2+Q���7�wS4v�Q`��{R鲞�Y�h ��.����}�}�  ���F���|&}�B6���V�X4r��R �\�6�[G�����: ���&���}�)�8��>���4G�#_�s�B�[U��`-���K IJ.�B�՞ck/B�'���|H�rpU���,��\�0|е�5H�TJtȁL�C��7�/�ƪ0dI0��wy��"��$�2�(b]�0c��`E�Ǣ��������>��Fm
 lu��@�P��b�f*
����7�`"!�dy�^;��|�1 q{��5f cjrv��(Gk9,��=nm=z���
�!4q�(���s"��$�&;.�X<z�p�Ӥe��
�Zv�^gd�u0>v�������8�2 ,u�?�(� ���t	�΋ [X++>��wa O��p@�*�ƉG!��N���+�\oH�'!�˧��S�W\^1�%��e�8�a[������ɨ#PA xp\z~���3�(m�C<�޹�FCBq.��ύ];��I�wD%�ZQ= �%��[gLP�}W�~�
�� �
8����t,T;�w���� �|vCt�*�GfxT�j��{J'N�_�A��nNC�R=��_��4l9�i�~V��۱�Q�����mS�I�`l�ܯ�W8du��r���UjK�7rh���1��(<�-�A�U��R)F����A`�bE*���Sָ��ȴa76o�������<ܔ�\��'�����4UJhk��4�����ɲ�ݗ�������F	����;�1[D��J���%�R�q�$m�l�:QR1`!����������dI�%;�5|L���uo�Z
N���~� $�+13'�_�*��6-D�p [R�k����>����&=}m����G{C���E�U�m����|`��)��BU���\{�.�{��-��A����T$&��-�
�7V���ܼ��9KB������I=U�c�,����(��2�%���ō�"�Dhn.��x������Q@`��O��~��o8��O~d�2�3C�Z	��Y�������L�Ƞ���?_����rG�ԥ}�L��Nk&[_���,�(j�%�p�w��P���P�z��i-��1a���)� g�k;����"Y��MW�A��|OfJ)��Ȼ7|E�+�.���A����ncqm|tN����h[�c�)~�0,T5L��E#fi��|,�uUL��,��5��J�^wE<7��EHF�k�õ�����ML2lL��-{G���g��<
���V�R��C�����bє�ﺪ�.��'>�/V͒�|�~��Dh!,�LI2Ť�o�k޴ =p: I\���1������˷��Z��H�<<�&���67�[���g�W���2P)�R�ts�Lr{|6d�7�/N��\��=5�V��X�n��L��<#����|���(Tt��j��8�?��4ZZKd�.����;-���N��ʳ�!Pk?�<��P�������6��#_�W� 3�	��C���UM:K��b�~����1ݲ4����ke��UX�����W9��Y�ߘ��:q���{�������x��a��wb�5}�����J484���E�X���MQӷ��AG?a�M��	��F���!�OG�s�����c_G'��Ɔ��12��G�/V[�'q��5&b�>v��O.lZ+e��HIR��W���Y!`�bp�鬜���9��Y�S����"�u/X���X^�7rsi�ǟ+*a]��<�j9�gtǑ��o�X������73��G����ɉ8�������mc���Z;d�2,�W��B�8	ba�, ?�O�!�O��X�5�5�_��R\oะ2�����K&�y\�3����O/j���^�}eK�^�l?v�}�����c���Ƴ}.���NI�S������:�Z/S����v?��p��|�M��kRt}:p�o��:lao��@�cPxcy�L���&g��;���Y<�/��">�5}t�N�J5��JH&.�;7�\�7��7�u� �l�<7)���J�� x�2���:���$[C����`��k��Սs���� ����E>o:��4��I�P4�̣�S�6�F�a�K� ���g��_��F,^r*e)����Y��t��?�}tɊ���b��i&:m �]�����"������m<8�~q�!�B�e6�@���m;�J�v�E�̫h�Xz��N�16�]2���,�n�;{h����r0�G�	 B�u�z��lX�1�Hh�PM9�q����*x���#��-��#���y���j4�4�΅�|��NC	�҉.���Y���&�nV'x�Z(q�p���L�ݺ�v7�u|g��46���*�%\]:���̾}k���+�\U���5��A텠�N4�!�b�������-���V�F�N��?�7�Iy��*\*�e��E�u�(������n�D���j����t�t�ۅk��ۤg��\�D�҂��[�1��[`�������Ą���+#�Üo��m�M�?��wz����qd������V+To|���~�� m�0�K�ВO�^b3���ߘ.*���X�:��)f��p�÷a��7�=eX���%�w)�i�x/�*OhL!�j���u�U���fæ�1F��-�h����T\�|Z��x�T�e�����&�aV��SV���4H���b|βw�BGl5V��ҍe���A�-A^Bb=��tq^'e��-�H����x��@,���j����]��FM0����/�ڮ��7:���/�}�1j,��+u��ݶO�+;�f˚Pʩ��ld�O>q�k~��s헳ퟵ��)}��иTH����Z�u��|gJ�z�P��k����ӫ�0�C>�c(V0A�#B��G��H�cRi7Y�U�Y�����]Uњ_ֿșUm�?y鼾�q��U:��d%�����Ҧ����b7�����*}��a��~��2�A����f,=���*�$��ӓ4���Y���t��٢L��
�\,0a~OSE�"t&R_��A�盹h��޺r>����֔՜��햩���V��
x���bO2�$B$ѵ�E�-T��E�:�=��:���?G�"e�̸�z��,�LWB!F�UO�]�9j�쌱�Z�8�u�(3xe��Ң���'���SR�p�������2�%v[��e��b�4��p�"q�b�9lx��D-D^T��J�	m����rG�����J5��z�ɩ��������z�]��o]F=*,X�z����Y�\�b��w��:$���!�ĺ��	�j�.��R��x���҆_��5h�<��F���W�{�.��#��Pe��k�PUZS!M�g�4�H|�v���l����}���yt�@���)��R�h�7�ɒ@�	�ԗ�e��������+�`$'?�	��V�vw��Z|�������t��
w��%�,=[��?R�#�9����92s��Ě�!w��w
H5�����uV�
{���;�<���M�fҡO�[�)�1R��̹]@y��a��\�:����yO��v�l�Z�\�Z%W�K_�1z=AU���szD��(Ġ�e�=}�2����VDK*�dNp�U���A�3���Ǔ����sۓ3z�j_]*t�Q�]{��qS��ՂD�	Yv[��m�	"�v~e��q����7�5p�o��t���C�vwg0�Ò����<��uH������Jl��j�e�=�����xY���G\?9��Ȩ��͈/�7��g傟�� ��n��*z���X�`mS]cS�'J�l�:OB��=�I��=�'�����"�/���L��D�?s����F2�Z�_|k��.�<<r9�<������.>e�S��X�}�DC�g˛/��e ����}�	KW�WU��BM̧��+�P��޴�Φ���7	���i<���܄,��������������cH8TLJ� z�{B�~�}J���>o���<���<�d��	mJ��)�,�� �~ڤ�]��O�Z�i��Ά.�
����	{���D�z�yX=�bQ?���o�5}��[�y���U��v|��LK�$rC�c�dI�G"�t�"N[,Ms_�0�E/04{�]��k������5ݦ�el̆��2��T�m��O1mGk����5KHmbh��܀hO�B]���?<c	4�.�嗜Ϝ�/)T��D�hX�K�r���OԶaX�x�(�'�L�{ĉ3�E���u�n� �����0�I����D��WB�z	�
��*�"a:�vOp��x!v����R�!_c�C�X;�v�DƩ�r��l�H���udu�()�����Z�>2�J���Yľ�B?���?^ڂ�\��P�x�TQ���*���I��
�?6-�^n��o�[]�}/r%���/�g�fwU�i�4_hg}��i�T��yk;����u3�o~��n���»�Q�M��/����1MV�}�a�<�eO�%�B9�/L�A'���%zsAM���?��{�.�*b�I����wWpO�#Y�h��<z��W#FPf�Iu��[��8z}�*��q�����ƶ+�j��cH��a�<�7h��BN.���d�w-�L��^;;Yz>���Lfи����L���&���	5>�;~,�-_��ಽ��=�aD�pOp��4��כۋ�����\��c噘�*=�'0��z�2�z�7�gWnM�v~�.�eצk$L�~�u�,'5J<���NzJ��l��E�9>��*�3�C[^И�������ʿͤ���:���M���.{R4x�zǄ4ѭ��|��^�"]A� ���,l�	+�?��'��P&Gl�A������v��`��3"��j��C�c���K��2��͝�~,/#I_�����J���ihjV�\S�,��*�{�HD�#k����Ϋ��j~ �)ڜp�/KK����wFd*J|�R�`ٹ��-���}\	�;rrL�{�L�Z�|mD\�M��=�Цc)Go�t�5G#��t�>��>��!���&�F:$��ԙ�e�W�HR�a���v��m�1���N���!o;	5�p�fc����F�1�����-zjڳ�Yv��>HG焞�K|�����"�쫊ܷ$����b2�(���F�B�d��B2�	�K�U4ݝ��8Y+��8U��K��=���� ���V��~���	��p����]����@gz:V�B�/���@�2��ؙI�f��K/Q15jد�~ov��$j��ͫ߰o����?(P�K�}�2���UG�RdG�8�N����o!�<��%���r��fӪ�2���y���4j��|�˵��`��( v����������1C��>8�%��7����S�� ��]h>�l���-��\�Y�;d�''U���m4%sŔ��:Q��ty�k
�N��ӓ��q���m�@�gN�
SDk�D�7����^3�-(2�,��������_R��c�8,��K-��|�^@��쿕�Mj&&RMYcq�D`}���2�vb0��&��H�[���j�n���K�0�rv\wwH)�e��!ۈ�j��M:Mv'kkt'C#�����������#��e�w&PD�q
�g�G����E�s�4l�������ɝh&�]��P�xi����&�y�j��|�U� d�>���4���^��L����c0���ȇ��c�_�����d�����2�p=Pdgl�S�������j���Q�*�R�l]H���������<B)�$���i4�@/��O2��d�K}�{ψ� Z}��$�?�ҔZ&�%;�K�<^Ȭॉ7����>1Y��u5����S�$%�����b0��M�[�Ӧ���/|<$�a�ԛ!R ���N��MC����9v "�n������p�5��)�ܗEj��J�%�f��h|��1i�'��ikR��i�U�����=����l��[c"�`�oK~�^�N1��
X�p7ׅ��֓>%22AĳM��U������jJ�,���R}5���H���������3�[$���`�f�_�d@^�ܛ?(b�1.�>tu�G>�'�����=˜�� $-
Pd�.�]�M�c*���K/� ɋ�1u�ߩ�`�ŕ�γ\�]S��:�h�q�%�Ӵ��t����=a�d�q��y���d��<��"��W���)�#���
q�{���S��{r����A@����;�8W���|��B�����I���c���Ft��3C
!ل)��҃1�����/�m�nt�:��nF$*��������D`�͓�`��Nd�P�T�5]��I1�^v~��3b2�{�}HN߾W�[)��QY[���z��3�_Y��YE���wxk|-J�KH��AҦ�
gG��5Ă�aT��k��53���Zl_����q�XT)�s�R�F�7�r[��@1k�A��>�y�L�Vڮ��y<wn��'�$�M���:5��,`��gݫ�Ĝ�#����j2(�j1C,�n~�]]S��"�W<���=���܍O�C��Y2�A� ��ә��W;6�����̬�f/Y����� q���C,Ӳ�-�cM_�f���X�TO��t����'LE�4��l��^���+�v'H����}˱q��<�\�@�xaOO����y��t8�$/8�X�$,
-z��N�����0Tg���d�8'�ӱb�L6zoN[
0I ��N����s^�Q�C�-�����!WT�˧���O_ʞ��t7G"�p�%!���fj6�2�;�k��1�U#�=V�hk$R�����.��.�_��l�w�gQ�%��d���;���_&C(�_�L�3��#'6�`Ll�d<<<?NV㛑��o�Y�C'�@q�*v�k-;��|�����/w��&(�j&�4�mj��ֽ�;��kW�t@d�T�nF����0�%�
�$*��,���c:���Q��~���0+B' ��&��AB��1X�	�e1%�X����YT��!��ӧ��������%vS><�ۍ����ĭ�����H�qo�� ����r�:�����E%n��=��]��i���#���Ҫ�;��p��W�ZX�+H�{Nƃ�pW��tVY�]�O���A�]nDn���J�n�*S�ԹKA�9�Q��%�v�N�乼���]i��e0�����;�D���o���1�䬓X#���"�����
��Q5����VW�8��_�JXS�wWg��0���.Z�=l2��ѹ��o�Y��7h������z��o�v��D6�Q��rpe�w�$���M�5g������ԓ��W9�}��B?����<9!�f	&80j"�����M��v�xr�K�h�{yݛ��-����
��2�g�?I@�'�Fc�]��٢TBQ4��QI���wVY�$N��ħL���s�&Ҕ<)5�Cr����R4�
q�$�6��jp���8:�̷f����ٸ
\˙@]��T
0�2M�5dp��=�z_��<>����H�(�w#��q��^�?�4RY>�yE�<l��Of�D��ː��"���-�����U�k,d}DV�#�9���ˆah4���'>:鷺]�8��1�a�?/	/�]��"ND"�&T��m]����p=�syh+
,�����]v>q��`%z0\�S��.=���)�F1$��p}��[wy0CAs�!�rvo�F�[����7�&pc��U��.���!c�-M�������̙>�L\4�6�V'�|���bN���^��ObR�=8��,g�uK�y	�nzFʔ�qs3��d�?�G��P'�f�|V,�������VYB�oI��2?c.ZB42~`����M#Q�����e��0q�:�������w?��ow�g:؜��#�qd�Sj��-]*Cꈫ�aۆ[|&���s��4��7xsW<��&���+M�Ia/m<Xu����/� �[�_�Ԙ��@LU��l�/CN�Ĩo�B�����'��ߋ��O��P }�Wg�]h����9�鱴>Z>R�U�Ȉ�q;�{���/�p�rY3�}$�]f2v�GX��M���|��e(�i��x�5mr�x(���o��#'�mF��H�?H���D�'b/���Y�M��!T��[;��ë%������^^��co�cZ��M1CG�L��3a�ZA8{!E�ÎhФO��5|�d%37j[����4g��ۮ<(�a\��E�z�g��Q��<�g�[TRF���e\�t��YZĲ�}�>\��|c���z�����>���@:�-s=��WQ(}�T�wM��z�2}��1�I~�e�,?⠧�B��Af�X f��z��9)9x��S�n{�3#LX[5k���d��|;J��O���PK-�ݷkz����UY�?��.$�[�싶x���4��S�S>�o�3�4*�:����y���T#���PFrv^���"�m!j�z�w�H���!o=�bV@�l���<�����k�'��64ܜ+0��gfC}�n����&H�~�5Cb�켧%Hl��L�!&�ǘ�us{{^^���*���P�� R�L�1˖R��"�k�,�����1�=��?ELF����g��b��*� o��?L`��������Q�}^��I�Y��z��'�22ѤPՈjCcmSK���1dC#���KDȯ�	n`��e��A�t7�Z�hh����+������\�����O�P)Z���rF�>0n��g��&/±);�J�R��9''���y�t_��wB��wOd��y6(��>@��"�[Q����3�6d�ĸ&hW{6�A��	5��c��im�PV�T"'G����k�y�����(>�<��e�&���n�췷A)G?Ցse�������?>&�\R��(��[J>~�ʚNDl����ż�{�~�2��Q���$-r��Z�uv@[Q�Q�#}��v��~4���~�/"~ߢ��=)	�S�=��������l�]^#.w�&��7+]�~�5�]���$(�����cQ\�#���j��kcƼ���P�Hy�bU��l%%%-�� �v���8wm��;�����bbE�+6�j��ճ.e|2���i�Dͦ�<-)-�UϳhC�����~3>�/!������#�q��p6�GN� �\l��SL� �J���۱
�����뽵���6�n�t~:��'n8�Z]����R�/���;���釼BI*��7��&�1T�k*�o�����+$�s�djm8vX���@C�����Y�
��~D�J�<0>(�#C7�)B:%�@��1���s��<;Gv'��@,}���Q$��*��<(>�2n䛅*��@C����[?��h����5>w�\0���}~�ozl�i'�Rk7q 󲹄^�3�c���+��yzBL����� xJ0>�(�ن90�m܈��5�x2vV!㉃��	�*�YR���佂��d�	-�z�3�?HAې�� ����=ڔ�����(O�`|~�Kbd�����F�	dg�.b��(	�G<xXӭ�^�S���<���_uM�O�� �R��N�N�}��djs�xĈ;�1�3;�/Ԥ�YN�a�cIl��:ބ)�?;�x۝wֲ׸F#3��\S�������ٳ�l�MA��VL]$���ك]�B��]���8d��+��HyUuk�փ�A��(��56���n[F8�<�uM�Gg�0��SD�8<�x�A�Iw �k)�H�8Yr��������/F�`FN����{ߗي\�0K�ۧ�3��O���Wr����o������%Ӯn������7�������v������W��J���6rY2���ںAO�mn��+�����"n{�1�ޮ�򞞬�©?7躕k�GaSÔ����gX��s/4�Eu����up]x����u�ֵ�t��,�Pȃ͑sϢ���esq��đ��[�U"K[20��"JA���D��#�y�p�,\?[����^�þ�*�J²$!$'o��I�z��֝_qsk['Z������V���a��G( \3Di�R�ڟ���zL�|ı�	}Cj���x��/�w�`S�I�怟��j֚� ۯ�QA�c���������q�k�uG�I�nX��^���!��{��d��{xQ	��C��E�l L��,��'@�f�'�\�^-����rB�������B���HX���A������<x��W��^�R���lEIX��P�?d�z*��e�tÉ��6v�����0a$�Y�o@#lb㹏xE��˒;��_�kh	�0�d�C��qAꈄ<Y�IJ��|���iǲ��*\K��v�[�q,�V��J�+��/�w��'�`�� w$�"��C�g~�M�����M�̦h�x�v�.ܪ@����5�,�3(/�(�|��#��Č�f��A��A <پ�e`��d�*��!����t��j"�J8����[�']�X��ێ%c�hs�G�n�M?���.l�#h8^Ej�i&�<�u�@ea�6�����]�i�"���J1%�0=��n�X�O@�������"���=���|z=�ox����+���vTST�h;` \�0!��1m�}�cmW7���S�xpk-��Op�{P[B��"�LYB0�A!5w���WȔ�Of�c�=����M��9�<��Wσ�T TY3�`���<��J�u��\\ �Ux)0�f�I���������_���rAG?������8�[ZR�l��݁�Z�_�� �9��S9��׊�KV�da8�%�	ҏ���DJ�NŹ�|�����M78�������"~��~}جα0���b��a=_���\eq��b��0��,L�0��O���Ǐ�����]�UDH#�o�a>�M��,��X̭�'A�{��E&G�Ir������9m|0�Ӕ<��������s�<d+Kވ~PZ��(��r����@<R(Ts4��I2v��n�%���B��=`��I���H�}zo!�p�#J�S�ޢ�7m"� �˃�5k�."$L�[=��p�#x&���1�	��	0H����O �$���my�WoPE���-���"JJwwJ*!) ]"�]�����~����~�'{�^k=��u���/jf�8J��N�q\�bO�'P_�!݈�����C1A�"v!P�,5��J(��=ǆ c��L 0I��y=����mh��S���x�Z�I"�'��\�z�U<��Rb���}����6t佫���IԩA��p�h�id�Ȩ�Bm�
����_ѣ!�~	m��B_4v�t��]Qz�bNذR��	('�l�xy55���?�O��2��ya�~�-`FHq�}�T�p�H��:&�E�� IY��Im�p�$�Eϧ�����#����*`�/#��LM�-���Ҹ\{�E�@ђP��=>�j��M��D���o��L��H����bIUN�8�:����ޡM^`�釛��@e��&�����WWR���Z�7�lP52�&2��,�_?cE�LZIw@A�@3���.��-��q��^]B%Q�ƙ3��H����~C�ꌆ�m�����6 �d60T��������_h�\7����ψ��K��j+�e��xk�����B2���n%3R+���:��:��R���1�����%��6�~�����6��+�����F���������\�C95#t�:G<��S���f\OaBe��I,�=k1�FJ�&?�Uv�S4�>�c�Ӣ��#$X
�d���0���썭��y!���4���3Lq��΅��
|�A��b��.����j�t���c�3��h��0mw`8�((�2iD%��)����t?1�G,�8
����:4�T%1p,�M��Tmu��)��˒��H������M�D3Ks����@W���ϻ8���ՔF|���H h��L�,������";@d�V�$�BXsj���YY(����,q�� �����})vr�gHaL*E|,���|�$��v��8L��
��lZ����p�B�R��<�����V�#�1,�L�`��0?�R��� �~�K����h������ժk��>봹[ֳI���}N)�R<!�ɳ�j���Üs(���i�V�7p��W����� �)��r���m�VM���c���Cuй��ot&�@ب����
�4���ĸ�x�&\,Q�t��.�*��� ��s7�@F)�g�#H�\x7�f��G��i}��ei4i��H�Y3F��X���e��7��'�UAP�w=�A?)��r+��/9L�ٴ=~��Ýҏ�%�^���xE���J�Π�-�����r��o�'� ��q'^}�ީ��b\�O�����LVZ�%�7$�&U٠s��q�p(�F����j݋� F�%���ߛ��b�"���<?AE,��B�0���� ��mc�IP8rU&ZVaL�����^o��9B�K����\qӱfL.fXF�UdR����S.f�{�<�$��$�Ɠ-v�T����*��q� 	��r9*�d} C$���kUeec��a��uҕ�^%qw�h�-������B5DM:�Wt'��}ŕ��a��ox�{��&ic�/��������(ȟ��X(h�&K����V����k�Y���X��x�6B�O=�o��B�H��и��Ջ�zc�ǆ�5:R1�ԛϬ���~�TT�s��B���/�o�Z���ź��5[|z6
s�bP,�d#0d��rA<�;��a���>r�}	���Aښ����犙�z� ۙ�-����`b]vn�!xc+�J0����k4�wA�GN��(�}�<x��̮�û�+u�.�X��ꕒ\���#TL+?��o#�%ʼ2��<iT��e�jp��Xl���+hX�����֖1'�W[�A�OI�fAHѻY�}��oOP] ���JX��w�7~��|�.���#l��*8���a��^�����'���J��<**ɷFV�Ӻ��x@V�p�o���{�9�j�l�	]���C�v�C�ްwǳ����i�f]���c���>Zo:�!NE�`�ot�@I#�N���]Z���4��K�{��ߙ�\(�͚� 3s1h���t9�t����ƕ��:M����T�"DN�&��j��n!��"��Y3�u�Ǽ4%�W����q �Hs �����8�Rb�/��nV��u��DtJ!���HW�B���<7��W��s ��ڣ���	]XW@���(q��i׵	\T`6vs�9<l���[i�����8�t����&]Q�S�b�+b�٨"��2���@�����}_j
Hc�||�p	2&]�^F�n��t�R���E+'s�8����轱w�s��Vo��7?������yjZ�S��A¢���m������T�*���1������'�C�X-�RΎ��|͹�tq-H�w�T ~��aʘ��<�n8�B8�� �'K��4 ������M��qY�}v�����_\Ұ�ҏߍt�Έ�de�g\O`�"�A��AVU���K���CF����VӞ���1���]��	�������=x#O�fY!B{��r�á꯵A����Ω�DI�a�z��� dnȔ^�|x9~�&��畘�1�b����It�l��c�Ϯ4�]��|�W檩� ��R������:�iu��A�O@O�ŝm�ϩB����9U>Gh9���b����-Aȶ֢��Pe�9[kQ}0S6��u��y�w[	��� f@�/��/�b�'�FV�u�G�(�h<]��}��)���?k��\�/���~ ��?�����v�7�n]�42�t���.O���w�4���3+��ԬUh�D7:0h}Cd�R3��Ar�Tcp�bvW����ć\�O�7>8K��}���"5>�Og�e@C5GD�P��趨�97s�(9�B7)%
	���T��0�F5��Nv|�`L%�s�I����?�mf�k��p)�И����~(����'r6������ �T7��-G��0��O6��e���`�O$�J'��Ɛ��х�K�(QS'�ͱ�*�m��WVg��,�Sr��w�<���TOK;�	:���*-:�?�}�G�ǋ�H���գ�-���&�������v�2����	jW�����&K�|��KI���IV)��d�<�$��>-�c�[���Ɲ�䱐���aMe��ɡe���؉Ӡ��D�_*��Ci�n��q#/$�dv�"�)#�8�W�6��їA��})�S:||8z$ldżYi�'u27�;��Ԣ�6��$�;�ԓ|0�B��a~\����l`�� ���YJ�lt�a�b���,:�r�qiǵG|���H�/a'M[�)��L8Ĩ�ze�{��B'�B�1{��lM���j��S��}�����_E�Wז� ��OK���@W/��z��'б�?hS�E��H��X������rA���9��3�Q��񯵞���zB/R@�E_�]`<��%�ʡ�����+'�WP�^KL\`���NC�s����ӟi�v��:,�-�g=�4n�Uk������������1,��덾	�Ũn+��q�Ql�ʌ��rP�Z��?�ݙ"4�r�e�w�.���xSn)y!f����ݻ}.��=����r��/i��H��c�n��)"$�1Hxn��������f���A����rZwbp��yw� c���1����Ǩ��M����nPE��K����{��s)(*���x�ɐ~����F�
9/���v����Y7WpFgA�̉C$��^��-���
Mh��CC�q��}@ F磗��a�L�[���^O�#ie2�r�DƜWd���QO�͝6j������3GoX�� &WKf��T'=ن�;�z4����E���n�}B@�1�絿�b(�7�qrі��ի�Js��5$I���q��a�ㅚ����?+qx���	eD����n�e,�B��܃d"�|T�#+	�]kgX���zQ<��&~ԍWϞJ&TQ��W�"Az%�s�É���CPp�:O�_sd�v`����U)$�wG����b��0�w~__+�%�W�*O-�=|
61�GF�|I?�k�QkFI&�Y;�����^3�/ݓ������U��U*͹�Y�K]�B���zN��/)*�{D���9.i���0D�C��8�w��h?{Q�*���7��Af�@���	 6��*3�H@_((��-B.&�/w8���K���r��w��t��~m�.�Xo=� ��%�ه^|� �Y�����c�՟�ؔ��|��HK��N�M�+-�=�Ӄw�����B���a�(�:\�/L(I�-B������D�W��N8Ҷ��]�䇜��I�B2{�K�G�����-�7	X��w61ĩ=9%��'���{�<���*�W+(��@�����
��0	�Sѯ'�+s��L��j���*{��O�g&��,)����(�-N�ޭ�)�l1}0E��gƒ��r)2�8�œ��K���>u6��q�Fҿ�5��?u���N�O��i����;� �3I����d�m��N����,BV)� �X&E�y��_ ?^�'M��=}��⭌y �}���*��x��-�&b��µcg���7�t%���g��96�2��?�'˷ �h�Z���E�U�%���>tH�G1j��2j�	��e�&7���f�4�XoN�Tt�z�h�GΣWeD}WɃ!)��:��JJ3ã!}�י����頼YIM�O}d�3 �S���s��[�\\��5���=�'��k��g1���Ϳ��u�q�3q1m��Vvغu0إø��F�h_e��I��"���1K�\Z���$ZG����S��TN$�]�C�םTj5�����J�Q�W@*%[�E�6�Z������[�\m�k>ʮ��dD*l�{�z>te!�A ������Xy49#�ة ��IL�!�����U����q��x��[w�Q�(��?�]�8�
�= #�y��3쫝ď�m��#��Mg�ؐê�d�3�/�f�ƺ�^�JNi=�H���%�� $�:�)H�����oձ��K\& J��p��CN��"�bM�&�
�T��d�g�{�3#R[�8�y���5�ݖ'�a���|�|D���2
�����{�453J��{8E:$t� mؑ��:4.��[tl��c �}0�e�8�y!��j��¥S������T��}���qi�'Bi�3�����,�z-Oæ�|Ԇ�N��,W����I���Y\�q�4�Je�XZAC +��KTqͱz[P��z�&�� ��:�;
b�d�&�D�'�D.3ǖ�Vhpp�?���cW��Ξ�+�ϵ��U��.���6dWX�z�m+�B��ڔn^^F��J�gY�~hy���1��M�٪�GN�w��o�X�a�W�Ǘ$v ����C��fpeP��b(�J�k�O���S�u�pTM���t�ͩ�F
�'%*��"qﵡ`�=W~G�ʓ��q��;z�ū�G�L����뗩�-��4>2;�h��`��������0�\���4nm�om�dL��H�&XH|��R�A�Ъ��RXlm~��"���7����DG��R���F��Xu�>$��'��� [���M�w{u!�\E��<�]ӑ��Bh�xe$mu�Le�.Q�z���J�a(�FD�����7�褂<C�N.��[�y��pZ�
K~�$꣟1p����oMm���O��Yz�UN�Y�۳�O��}��&7(rϥ?Qym�ᙛ�wO��̃@� �:r��`uZ6B^"VS���{�2����E���#�;ۗ�_�{v�$�jrm�����f��&���D�� �H�UMe�Eu�Y{(�OD��D¨گ2g�1���R=d�Rjj��;����m����!��1]͛Q��}��p"f� *�M�#q*\g49"݅~������Y"��Bh��^[�"��=�B
n��������yf�{$�a���X����Qe6�q�վ���������e<�:!& bJa[��x�*��a<|�4Q�L> ?��F���\���,S&���l�,/�^H	N��ϟN�]_}Ti�v���&�)���1��ㆉa��K\_�NJ�ĭ�S��~"I���|y�o���E�,piR?3��5��V�]3��w��%�3KJ����,0���$3������;T�$�*��w��j�@�=�h���g�)��-��bT5��OI�k�$�5��M�>�c7`T3��Xg��IP	������x����n6 �6�IM'XR��xԙ�^�I��JJm��l&���[���0��ؖ��p�����L~��vb�eQ��'�$��a�����4�b�D\Z��Wm~}8׹`�rq]Y����B`�4O�n߸��~��]¨ºȹ�)��c�>!f��:����5g7��7}ye��s��� �0����s�f�ҳ�ΐP��͛�v!@4\�<6�]Њ}O렫:���Q�r�u*Jfɸ0��mݟt�Z�a��#��KČ�%�;TYI�l�)�B"���Y��������kW�?�^g�ysT��	���M������n:#�溡n ��L��^1� �k������e���0_��w6����I�a�k8�JK�ei��U`����Tr������������m�q��ߏy��f�Rß$Ʊ�����������"� x��1���E|��V�)k�������� ��0�>W��;�ڼ�,k�\�wR�_���ԯ�XITmx ���Րde���*µ3Ocwd�7�߸a�~.��a����G��VK;���v���C����xo��9���Ŝ�,��MAZle�+���D��X��S)/R�83F�$~-�P�m�\��b˒�ڵ�hK뙥�ӧ<:�����8d`T�($�@@m ˾I�ȭ>��rl_��~�:|�g�f��jlT��_)R����N��u:��Ah�Z��e?U�����*����V�$��[�M4�
��RYV�;�Qe3̞~�r�?���?��f�CU���u�U����aH�¡�
?#N��r�8e��,%맿s�_C�n�,���_&��b���H��3%�%J�_mN� �7����f�N�ƒ_���,�?oǨ�|،�$��[��U�4��	Օ)z����KDDVFǧ��F�m`C��E����u3]( Jr([�V�s5�������7c<���r['��o5M_h��2�%.������Ƨ�MlN�����I��Ͱ)���
��.+�k^�8��s�nk����b\�L�o�}��� F����������������[?*�^�vV�I�y�'�+���D�	W�����-�V|��gF6a��M�}卆˓k��5�՝ؓ���'xD��u�'x���cհ�������t|l&_t�h~��G�'1���AJd$�t��q���.*�G���f�w����^x�1B|o��x�J�g��
���>�ή9w��>�����y�������(�\�;�{���F���5��O;�Q��iI�<��/��-��*�����}�|Ƴ���S9�r��Rǽ!r�飢�b`�Gp�Еl�C�L���#�o�z�fä�Q7��e��fbֺh��	x�Ǻ����]�@
0����>7iuD����Ր.�3uzoi��ϡh�Ф������V٭�B��B��T�����'ʤ��J�l�A��OUM#��P �-L�Y�z���p����r��ۥ�ئk����=B+����4^G��u�V��k���slh@y��,�
	K&�5�#U���L�	����ՋǞ��e�fέ�^yPt@�C�fm;��RwP���5\�E���	�ޯP+ˣ�jg�f!�:a�Gw�PBnƨ�~Mp]&&�a�d�F�"�l�[Q�`	:�F�ė��R�k��^�|�:��s>ٱq��1��շe��WK`��BIm`'Mv�Uװ��D�����	T���Y8
ٞ.�>��}g���WYV9R�.��P"76��Z�4%��	֣��a�DT��R]!����RG��i�����2s�KC���������9��|b�%A�7����xw���3\2��$u 2�G�o�_��
�	ĭ������S�W����t�q��I
j2��î��)�.����f�?���h�+i�|�Ϸ�y�&�yýE��keJ�\��o��e��t.zx���b^n'*S�S���p�c<�}o��̗W_?_����'�Kѣ=�� ٓ�x�r+����.)踩BM��%����5m~`O�g$�!~��	�ZP5j�I4�L��Wg#�Οu:8y�����e�����MB�i"-(>O����\7�z0�ÜM������􂀞1q��aL y��i��t�B�C�t�_8_z��ve�a#�d��w�v<~�t���'A�L��]z��.�V����܌0�`��NtcƎR:m�ǋ�B�e��o�<F��B�|x�zz�'��uM�"��������H�q����so8��y��]_G�;m���� 7]��#�n cؕ$�)�L�~�L(>Ul3�ǳ��g�/3��e�8������|�0���ޮ!��*�悇�.�b���C�r�P�a���IR( ��N(��IR��
�l�UAn±1^쁏1P�Ig"
���Ѐ�;�0�;�Y�)��EV3�Fb�䅍��f�- ��\J�˷hL��uW�tA}�y�iJ��5?�z$���؍�"���8{
����z�!��	�2`�CC��&S���?T03��~�e��Q��ڌ>�3��fr��&ǫ�l�yhρwɶna�\Q;H
�U��B�"�E�8=��b��s_H�[����~�L�L�y�1lh��������f h�gA?���1
I�A����|�����#��(�&iu�hP6�,ўWoh�{׆�עm]ߞ))�?:b0E�hV\ĝxv���~U�F�^��(�� x6�$Vf����%j�/�$h�6v���]���B�v�3"�W���o=t��8��/;Ң-��Ŭ��ڬ��ڸ�7ա+��� \[��F�z�a4�!&�dɲП�X_>��w�p8��z<_���%��f�� ���*�U������ݢ��K
K��
�N�o<����D�%C
KG�ͯ�K�?�<�=4i�n{";?|�d��Hh�Xp@�}>��^���n����ilp�U��V�5�j����{J�i������28�`����!��+���"�+���i��t#�v8���/�:�܀�l0����;kB��L>7@���#�Di�T�\UM�=S���,?�W�'��y���/���;A˸4�E��-{%PEUO��chp1���A�l'ĭ2G����7�a�>�����7�j�F��[C�d�S��n�.�������W�x�;O����	��OC�Ō	��x���ڟ@��	��&���m�=(-)��ʊ�f�^�骀m$� �g8�I|��kϱ+4�%��z�:2}
���u�}>7��D�Ȥa\&�Y�#5���	|�i���<u�|��Z�d���P�3�~urN��4�k�hBڪ�-v��W,��v3��L��	;��.��mcЙ= +Z�FU|�ߑ�Ժ�u�'��񉢟�qh�!a$�q�b�;P���FN����s��I��t�������`�%�A?��gG����.�oX��R��f��3���=GN�w��JX9a����h��sSYxl��fU��G��k��ĥ~�6a��-�*O�|���zq'���|�$�t��CS!C��g�n8�xa� ���l7�y�vjl'yY� _%NP�.-}Y��X�:O��A�u"S\���[��mh�&��GU��~�^�T���g��81��˒� �	G���]�^7M�
<^4��r*0lچ�,0�O7:����h�O>����4��ޭsQ�2�$f�\�8|� ?A/��^��ſ*3�XMA霫���J<$W���i�	�?��gOք�F��������lҠ^(S5f����l0�tXX���5}�̾L�3^�c}�"+,��AU�Wy��iK�5�-V�錆���a�r��B���i���؁W�td'& ��G5��'E�`B	�E<q0����,9T�CLY��O�jW�b��K��f�{\����>M�ni|Q�b
�ӱG^�J�W�s���fp����]i^q-���~oV^ܫ��K�(}��5�A0I�ڽ#���k_�Q��<��o.���tA7��Z-��hw��8ȃ)2qwG;�?9Ы�E]��g�>��˟��A��:�4㛘F��D�����		�|#�n��]Ҋ����oX��P�����H��{6�U��;Y����e0�sT�iV��0�ߥ4iI{�"������o-����tɸ�O���ܞ��k�#$ie��M��u^��A�!��ϱY��r�Vx��VRo{&�z�M�v�����әy,�!cZ�1v�C�.�G��S���}�����\`P���!'$�t��f�ȤaU�~��Ro��uAk"�j���7��A��_0�x�H���B�LĘ�A������po����V% w�s4��7��B	��"(GL���'�� c�3����~�*<�)
�H�.q@_��3҅�1z���8�$m������I;Z����w�����ڣ:~gg���S����cu�����@{Hq�n$ay5�4WF�~���(�(�5F�����l۠B ����`S�ƽ��}+��y��s��i(�ߥQ������p�[�@�:K3"�����Ս�/�V�U��X���4%$�'U�AH�뎸�?���*�����"�NϘo�z�����au��W��]GbI������@�+�Ey������d&Oʘ���A�$���Q�J6�Wߖ��(�;-�G��T�ڞMaq@~����[�n����p�b.���������g��K@�'j�8hLqq2�`j�T��FxhU���-��Z)���R$�p2M��<�QD���2'>wO]��^4�N4�Ov�v�9��n���n�5(��k6��:o{��aZ��C�U�8{r_<~.�3i�&��~��x��&]�",3���s:�SF˴��^C%P����k#��(k��A_)C�*6���e;r<�ϳ��s�:�'0�LS7�%.�.�XT
&9��	?�.\�>���6H�o؇���RHC���/��	�y��p�bF�,:5�A68>�$+�+eI���I�i|2��H7��X��		�9e2�_��PB�J$���m'� ���uk=�鷟Oy�RˏC4�_.rB�� �D��-���!Z}�d�Iy����}i��DŌ���œ�9��9J�T�tb`^"o%�)�"@�ǖ��⌵�tNM��a1���ʚq�*�����?�r>�DTF�ߚ��	��=O�[��5T1�C�뮻���B.Y��H�U�|-( M��f�/��ȏx��6H�����a��$�5i�ZS^S�� �	ix�.p��e��ƞZ8���a��F%��*]X�X��q-W�~X��`d� &��Ű�Xd��$M��C�jTQ��v�"���v�dGf1�,���**���d�#��?xH;��C�t���3w�9��#����Ԧ��gb�]y�����\�=�5� ��o	���eZa�"���K�o�Yh;��c�LG�PU��u�x׸38^D�:S|��P�|�����i�y��c�'����hb���v�B��2�)?�IW�$۔ı�u,�ǚ�z�GG12r��bΕH��Þ��Tț>�ur��b&��,\?����<yr�n��L~WR;a�b�)��#�t��Oq�b<�bHb��E��F:�0 g_��R�Eӽ5�������d���m��~4{�����Y֒/&�Y9� �\���Zh����Qe8o7]�31MF�1B�8h�C`�ʙA��!�'�9�����#
g�Z5@\%ʈT��%p�OM��f����9� y�"���F����o��̕_�A6MJ�"4�zz����No.����jҝp��H��1���'���Bݎ���\#0㒬���3�f�r�c�������ݧ�'-ZEm1x�8��Ì�����7��J��3X$Ӕ�jŰSE.����%�;�+3_��+��e��Y|�L4����7qh��kr �~�s�ȵ�|�5��&LM@�����&�ԥ'T�!oL���E��#M:�E��]���\�u����&㊠7��[H
F���*�1�lV���ʴbQtc���%
798ҵ�̈́M��R��E�m�K�� S�ӯu.*� E.Y�ݙ_H�GS`e�\p���O��*�E=�?PM6�MG�n���](�@)���0�ܖ��|J[j�.�;`�;|;�(�#VJ��� ��g`�p	{�0c��ʥ+~Hn��{R} VՑ
��g��HI��[(�4��ٚ\)�Ż~��?�Z�!�v4ց⫿�y΁�-c�v?._���Q�i��-x<���yV��}�4�L�ȿ���d��7%w|��䃯���$��4�����<u�<y�ŻYk��M{-��l�"�
Cww@P��Z�GHH�l�m��:oI*�Ed�Ou�8P��!W���q�������ߢ=1���`��]C0���x��������^Q���MG\�>�&#�A֔q���1���{jV��b�6B��4`�nn�ut�<��'\�?�4>�`	S���4��/f�,vzc�����'\���� 뚙(���a1���L�T�����>�
�Sr�Z�
�˟�$�f`X �^s�8=k���JyiJ�r���(R-@���I��7��۲��bt��,ZB���g�*�{�X��Bw�{�G���r<�i��1��OS{��N�D�G��r�k���H� Q����r�F���Z��ϋ#��<�(�	Eۛ&K�/.�4�YV�����a&U'�t��F�eؗ;g*��#+/p��~�>�������%����~	X \{�F��C��X ����������ɛ$6%	���+��ټUx�=,����=�L�;~5)Q|C�,I����{w#�w�-���n��t�����K�9�7)!����^�$�|l�b�1�w��I�������'����v)n� 
~`97���fU���~v��[�@(�>bM������]���;���w����yj���$S�6A��v�):�R�@~M?�q���t����� ��V"��-��P��qǼAr��V &��	vQ(�����Tz�ӡ��G�x2��b��X$� G�e��L+Ѧ%٫����9���y�R�ь��>�A�(�aa�Q�]^Y��a�[�Q�_�\��F�0>(O���l�����0>�:ݮڞ��>`���O�JJC����O�	�x��j�/���ښ���&��D|U8A b��7��%�������KlYvoa/������(��Ԁו�p��ED�x���.�і)9wb�A�� ��տ>�P.Y��T�T����͏����؟4���_h��DX	rP��X?�:�,��X��m�
���%��������Dt� ����eS%$T*�~Lϸ����� ��%� C}���$|��A ������,N�N:_r�Oۏ��I�:��[w�~��_n�8/�J���ȷćP�%;l�Rih�'0���	Ü�)~<����Ї�Z�u��[�>߸���x�``(�n�����#�:f�7+���4�E�t|>ߡ�"l4p�����P������nk=Չ���&��%��`ʒ7�����=�;��{�3"�x��h����:F�����W|���$TT�(
��0Y�'�����ʯ��P��x@)���A&�����9���|���D`؄�rֽ�]6�8��lv���MX��cx�����r_A�糰ߌ�"���aq�13�;#�����o+�Z:ӭcڭ�}L�m���mUlq��w�A�n�K�i��C�iM
�?+����?t)u@����X�ot��&������J��-؀�����C��G�nt�����7z���7�"� ��T�|%3��^|8}�=�4u2c���9N��cB���b�,-߿�����J��3Ƭ���oY�<&vV�V��l�Ϸ�-!��D��|!�3)=�r�;͇}�"!6mq���mB�!��R}����U�N�a��P|Q�Ɋtd�g����`ZKR���r�h�F�$:Hn�VF΂Dppt^)�V�H���x���|-]�$����]p~��2#�&�Lz1m1�g3����L��f��t^�;��?:�"?��D����9��j���y�W��I�v+��1ďlx�������`~+��|�;���FA8ڪ����+�dFo��9>��ɶ���5��|ۧ��'>�%c��ǰA_���@�|6�Am-H�*ߐ;WTJ�(��D	�֬X&�PXQ�!�������c��U)��᭣#)��`:K�&��`^
�P��ŕ��|x�m�	h�G>�2��������3G-�|�\������K�O@�}P�U�^�Zm"�@�;>G�ok������U��蝧	{�y|����^�-��*��9M./�
uh���O�S^|dYE�Pgw0Tu#Mu+���a�U@�/$�������|�kjҽ^�,Ӻ�{�~��q �8oP�����x��E^�+
ʻ� |�/����U��0�s=��UT�Ђ����).�/�/pM���r���V�O���nҡ��I�]��С��g�gޛ��җk�]�3wr���b��O��B�'�\R�$'���ߘ�ԋ�$�\B����-t.Vz�ս��0i��^b7w�µ�li��jPHN�ޗ�sĄ���F��|h5�e�-%�a��p ���<V)�(,�in���	G�dKdyDrX<O�c�j?�D�}�������dVuiξ�n���8��ji�A��S��f����Z=���h)��� Y���[P�E������Om7�W^ե��u�>z�.B�|��oJ��[�W�I4_��[Ci��^6�JC��X��pqq��52�@�/<$�Zw~[���&s��H�R�����}�A;�������iܥ��L��[ �������
�D �_U���FB<~\���r�K��:��-��
ȗΆ�����nx��Q_-��T����RJF�����=������|��Wiz��q���$G�?A���*F{1��\��O�ӧ0��@5D��q�-�}U6�R�gC���Fr	�
�7�C�Zt=�c��G�R��p���P� �����w��ڭ�S� ��~4%�g��!���"ĪXP�[�}���hZ��ĻZ|�����pH��<�!{\��&���NYfygQg�Ay�9VI^����S�� �C�.�Ǖ� ��[�pF���;F �-bC���u2����]?�}Uf`U��j�.T@�kP����@���oҎd����OeHO�@���>��ra��-�u�����"T��k�	iߓ�2����\:�.����rU؋g?��+$����W<�+�4�d���sf
L�����2(�aQ���&nG#��ަ�E�Xͧ$p�P/����c��A����R�����ݯ���������lB	�,��\�NW��_=�?i���Z�c�`�O���f�gUD �X�W�2m'!x#�����P+y*�L�����0�~��HF��7r?!����֚�C�ö��5�4��Υw4vuX׽w��P?рX��u�&� P���0������?]���y��pF�6��i�֐do4�N���I������a�S/4��A���p��U4��,�Q����]S}�!hg�s.���>�
ɋ�Uȅ�ϲ�(�!�\>��e���\"N��'�*���s(�sy� H Xz=���Oِ��!�@����>	���Y���<AX$2v��.B�!��	���S���@�1�%��>oA�C�V����b�9���.�HS�a�Q�������"	�9�U��X�7*���A�h��Rc�U4��TB/6y�8�?��F���� ���1<2��D�" ���C�����ϟz�-D999����:e�J�o�����pZ�C�����Ӌ�8::�??z�0��c�w546�H��Z��
�KH�mm����jhhdee0002��=)�q?~�rnpS-�r{:��jyҹ���Ï���ef֪P���b�j�2��g�;���9��.�'^�|~qѵ���~j$)-����b��Ι����	��4v�@�t��FFN��8֮��o*�|fjj䌡�Ҵ]�Ɉ��t�q��b���L��'U���e<NtX�`ۥƎ���g��Z/��{�N4�z�F����HH]�E�l��2��SH$$$\�?'��?���e


L�e��oƿc5���XZj��QSS�?�e+�ozj�TPՀ�(�r0-��m�,��f�e�Ԫ����=�N��!�m�|���2O<>�v����7CSV<V�iƄ�D���$&]��@��/,�����������Q�A�O�}}}�O_�}�m�"\j�F�p}d��ˆ����I���%���LИ�Э�c�̯�6�G*N���e/�d�ZkC0� 4M��s�=H���B�QPR�|�����!��=��wN˯ IysuՃk(SkΊ'iaaQ���be�\�yڒ��}���ň��X�\7��P��n}S��9��2����r�¡S8.�v��s���SI⼐�`w:����I�ߚ�������s����4�t�������<�ys�+2=?l�0�d1}�@+��p��x��j:�x�����lYI6�
�I��Y��##��BvY���سcf�=�9"�8���z~���v;�u^�q]������n�����,+���~h�����}�w�4]����G0kM�9�O�D$�Xd�[M��jk%�V�5�1�599J���Hy/���C]�nT|����"�[��l���.�Q����=<44�eX�hu<U�f=U=�]l��P�f��W�Ҋ���'����x�Ls���߹�I(9C։�3z��"}�r�9i� {^GW�G�Fo�"��g��go]��P��[/E<v^��ƛ�y���4�2K��Y'�h3[�u��R��<�����M4rҮE�޽���U��m����7���-���{�����@VN��`{bp�Qjq@��\԰5A�h����=*�Ђ������(�R#�,55�N�2�Xii��t�$��-�W�V�,���.&�c�Q���<\��f�Ђ9�K�_�Р�TVm�{�n�S�Gee�PԆ�S�������ڦiFg	�2�����]��R`N�ii�jjj��߼y���s�Z��������E�st<i�zz�j`���TUU)��D����I�7-��K�����K���|%o��,�B[W��ĸ����0H�t����e� ��tVY���� �	E��$A|[ݨN�����̽2q��@(9�	2�:�jc�����h��T���(eΖ�W���^1����kll,;����}�S5�J���7��ztO����TE�&�l&����l՛�=��~��
C�Y##�� Τ�y�����CPP���;2*����m�<���� :j��m2������ tc�S^�lDN��b- �@+�Q���$�J���/�b@/�.�ʣ���a.1))��#�o����9
�
B�m���]�n������N�L����.�D���Y&��o��;+،��IE@8v.���K>�L{�^��G0�����7�}�Y ��L����|��]�����#O=�n���6#��w#���~�f���0�5�ɘ��H 5��9��`�����z���޿��o�2��e��u�~B2��+|�܋��.�gqD�*B|ngo+��<Z���Ջ�뻎����/6��є��6X9[ĶwdD�`w���t=u����xu��d1i9˿�+�š��iA"�VZ��l�>��ލ����VKK���h$���s>�A�[����ܗk0���_jf�<�~���3��ҩx���ǟ����h��Ј�"~�C�ti��o?+,{������{�K�*�=�R�H��:��{��Gˣ�w��f���P����:p�Ժ���S^������(}vqq�]��8�k)�6�K�A1���i�O4:�A��S����V=%��~2�t����U�c=��a�o��-g��*6|%][��Z=��;��]4��]-��J�v�U�Q�v�ZoR�}MQ�s߳�?��A��;�]p��j����P��h��rF���& �m�-�,L�d�d%&������DQ�۹�Q\�G
yL�'��@$F����]���-�뉙��i�̵�.��*���Sn*�n�y�{�w�/ql� r&����&�)��2�GA���O�DE�f*6�)A��1��r��8��������6?���k�<�)�P表�h)oC��D$�7Z�����ٔ�RI�o�R�-F���bÚ�jaz{��f[ޫ��kVr�ns6��>��Sc�V-��yѩ����'�^}�_�^E�?��o�������9��� �l,J����8�40���nPf�����%݌~���ƪ�}؂�)�h����l�踆��t���t5�]LNO��g����ͳ����^of��E��]}�����뷦�,�w��Z��盛p���6,�҆�1��dx)�7�־�rZ���t�R8B���Q|R����������>mb�Q�roqH�l�yX�=Y�+ZYg�����W�]���$�׿��vب{��M�D��c�a�蠟���	d08�ggg��K�LC����n����
ѡ�(fc�gye��+(X]kEQ+F�>;�������F��!�e���>���������_������NuD��6��9��e�#�ݩ�?K��X�i+1�t�Ň��*��ѪP��+���o��`�
�X�;6B�]�|v�L#{����P���[<�x�b8��%.M��6�aҧ�1���C��:L�W�c��	��B�]�L�շoߞ�?.6����Ȕ@��s�`zr��?>�����$�ZKJJ����p0�)`�֓��=���(������W_0B��$�5�����#��� H��3���e0���}�}�:^����9~����eMsP�#P��M(j�޼}���ic ��dc��9�~d<�T�|%MUM-�<�����	��8?�꾝���������l��B?�xy��,�]�-8Z�,K6k�h?a��o>��#�����?MAR
$�=�>�Z���]���+EgP����Xg>��MJ������3��Y�Ǐ>s@C�wz�QL������)\��a|�0��w��M��:�_yDULZ3bhr�����Z'eeR��zR w����"��8������vc��@���^�,wF�'�������VT��#>�*��Ɔ��J� ��?A�GM~����"�J**�;��LN�!l�

ĉ�	M:�n�C�a�gx�h� P�Mw&��J���7���W���ţ������{��"���1�Ŕ�F��y��W>��>5[Cyq$��H.��5���z_��z1|� �(�Sj��؎7�iVQR
��)�ӭ����'�0�?�y��{ڮ&�̭�xGZ������33��v��W�Q�)W�q;+w#��F��K��t��$!�:�'O.g��7:w�	���}a�_Q��>������72r/7��4����,4��� ���C��.����U���1d����)D �h?/[ͱ ��ɷ�����f�g7��oE��ݴ������~EHHu00?84t�USd�n+`�}����'G��&B>���.����L���M�(\�����[�	���-�������Xa�x{Ր:^��hQ�Y�EO{O��� ��8-�<�~�5���o��cz�F7�֒���t���D�� Y�覆I,����y�����O`��# п�$%%���k�h����"�7���̪��ɹ0a����ES9����۷oAh<��0r���#��`�c�03jM��K
a�O�����LU�q�|�[]__Q'�n��;���	䢐�@'`�2�cǰ�Ǻl�PQ�!��������L��:<�N��!��~q���#�:|�I�?ߌ΄�@�U!O[i=�%O8Ռ�mzILd��	��#��A���ü�<))����X����N%��Yw���y�z*�i�ګkto��2T�ߵX��	��!�s`�r�(AbA�Td����*_��dE�`�	����������6�����K�~�w��M �H�v0���A9>iO,����)�TE(J9�X���沲�ۗŢ"����98�			Q.-5i�_o2z�:*#P���	���0b��>�
=O}X<S9�&}�֭�iB[��8�`������׵�2��7�`���=���>H��;��3�c�GևX`}̄飦E��9�����3��C�l9�C�SSS9�K�S* ��t_���FK8%7'�(������j����F��R��T��_F����'������pG/�q����$����2`c؎��k��fBөٱ77[��},��w���韶ї��S"��T���+�9v�m<�!w�l�!��)��*�;K�t������1iT%����l/T�l���^%�`�.�.�3i�o�ld�����`��;�a�t�$$V��K�||��8
M������a�����1����<f'"
X�I�f�Ws.�A4��k2���Dy`���ɽ���(zW\,�
��MK@#3 �]�U@M��=y���:~JJ���ѿ��]AG^�L�&�l�x)��&#�P4H�`�{:4R�W4�K�~Y�'&��
����-��E�B-�Kdd|bV�]".�����q̈́�7o�t�j@�8��ƖX\j7Q�;��or D�8O�+��##O��hM�y�iX�h�յ5�~My��{3�����.9���Q	�- 6�4��[y/�dy�!��\��8P�@�Š����}�#��Z��=�5��8�o׷���7N[����8
g^�~-  Mև.[%桷Q����o�B��h&	y�%�Kއ[�/�Ύw��t�x�W��,ux�0W.� `(v.�8\Y�YK�����L�L��MP����>qa�|�M���[�XUEV�p̀����$��C�9���^�� ��	�c&���'kI&Q�1b�ь���K�aـ�=f��ɮ]�Vd��!`P���Wc�F(�w'����C������������ ��4S�z�98$D�*�.���0���G����V)GQK���H�b�z�EqW�]k��W���Wj�	��#��҉��J��Jk�2���u�]������s4 d�:&%k�fqi������ϒ�F����a�ٺ[`/�g��޿j�k����(r��w@F�?=,���K$T����hI%~888X�J��5euբ3q��%%��l��G��o&�p	�Ö~��(j�U�n����X>�����,6���n5G�Ha�c��wj�S�6�1d#�;�A���׏mm�Ë^}���#���t�F�B�S�q�3k�k�pԭ�ULn@bJ��P�5nͲ���	 ����G�nl0!���=z��A~�ڵ>9P��z����{dv8O[l܌P��&M��u��x�`����<�0	xy^�|�-��ޟ?�uQϑ��o���U:�yB�D�U��^���c�]�;�������oz��������?t�?�,��;�g��)��U�_�]���f��%&͂`���[������9���I�*Y��u�^/L���%�:;ǆ%z����)�����/�t9?F�4����'����fvG3�cE�@��f�26v|�*�w|����6=����� �'�W*ڂ<l%c3��uAZeK �ꑜ\�vc�Ңrr��@�9dT���Qs���[댈�zڎ�SE�NIc�����	u?����Uz3�V�Xe�7��������,�u�E����KVcΏ�MVX�=�/p��bV�s��/Y��ZWb�?�6�("""j=0��� �G�(���_iQϽ�s˾��ư��*h��B��O��M?�g�	���:�骷p��y9��FW܊��}�骫bV}���&� T�O�~��t-鞀 ���3m�B��_Ш>���u�G6/��}n�x����kY�@�}q�AQ�1߬b�B4�G��U��g	�ɫW65rEZ����`ev��v&������H�B(���Էn��x5��f�n���4ѓ�1����vNٳ�D{�ژ�	r�cxs�&Չ���Xve�۴��ь��p�8X㇘��d�9������˶N _G�7���	�|��EN��/t�E��w��B����BW��D�9�_�N۱�a���ɓ��6y��h�4�uA^�j��?��]���gprr��U���A�PC��>���@��ʎ���Vl @�4�+)--�*�Y밠=55�4�NPP>��mIZ`�O��rCI�뒱:٢̍���$$<-��Y(hX���P��@ZD���r�P3�����;;hI�~R���oh�>�ׄ��Ԙ��.)K������H!aO��4�[��ɝ��.�i��Ȏ0J�.���_g�ޭ��.��W9��}W$k Oֻ#��n���q@Zڟ*!�#_7uth�� ��!�d� � ^3�5ϫfƵr��%A�bzh/<-g�G_�������ŵ5���̀��qAq�@@f���N ���9�}�z�3�����c���H�������Hu�3<_n�J�3���`��"U�y����v��?�g�z����!o� \���[R53���'�&���0���dy�X����]{�$��FzGW4�e�	�f���U��֡fi��HrQ%߃!�el�S2��q����m��W��LJN��y�jզ*�c��ol.p; ��m= J�C�fUKBDz#��p�ױ�����#Q���	�v<�f!qV��Om�|�@�g�-������x�&���wI������/��/�!���=CͶ���1��Y<>�`�ZT ���)�iH����P7�~�{����5�)����8��������p��������m���{��.M@#�"A�RRQQL��Ysrr2:ٝ(`�u� ��B�T�E�_�'�����%�Tq��� �P��lE'�?���f�+�M8M�}�jJy�p���wwz,yEo�+�ŋ�^!5쏑���:3�.Z�PSSS�6ke+/ c�b�;����	���w����D��c��H
F�����Z������� ��<0�5�L7�|e�߿6(Ohx�p�� f6���:o�w��W�����_��r�\''� h�KK�e���(M�Bn��T�| \��d��:��q�
.m:+�����!##3|YY9]��ff} <	
���x*��X�_�&�}3bK�#�pgie��uA���%������$��AP��f���h��m��Y�����z���O@��9n&�����cjzX�7���|� �0�zBQ�S��x�l��p�gWF��+k� �)::;����W�~��͢�Ñzw;�~����]8≇G�P��`�޹���X�˸n! ��d���#e����ȝ�QD�i�ѓgJ�;�@ ��K��Kn����P�x��L��Q���P�jy��]Ґ?}�����	$,e���2����i,�4������<�G5���/�l��C'�4�o��ʰC��)W��?h&�s�F(A����)ތ�g0���B(��h�;�����C��K���~/PѢ��g66�;�_A�x� r�x��I�7G�:�\4�;���dDoQ�ů?E������㑬,w&����
5=����$��	�rrr�1�.+�S~���Q�ªϟ?�OE�`�]����*����S�vJOpߤA=�����"�R��;�q{�I��m3�(��
z�vr�����	%,�tyg]h����CE=�m�z��)��qK����߲5�(.�-1n��F��4^�`P�ħWb
���ӧ�}��O��{�gy��U��J��m�Oᓔ����j�~��~'mmb�����^Q��Hͩ��":��MS�١� ��˲Rm]��3��((-*"wqq�+=�=��@����||o�O5U��pjN祶��	��+Ï���_�����Z|����Q�/�����P��#�ti��u�����fUs��>�� `Y��z���@u=��[�'�tٴ��w�Y��������&��yVkZ_[�Ρz����jI��Mw%ZV�J8)�r��;���ЇN�~mZ��s{2�?�.@Ҙ��'�^���>z��"��?~]]�_مu	,S�*Ć2E�:���44\����ꐗ���
�Ͽj�%���E��_���Tmʃ#�zBa��J9��0,Q��o���d�ѹY[����LZ�,����y��b��,��w�wd��˻Y�Ӯ�~N������4`�$`է���!�o�AW�����)0��I�/驩�\��r3?p�F\T��/�zlG�P>�[̌$�.$D�)wjQ<�7e����$������pk����p�R�����U�������ӋM8,�n�����0�L��c�Ǐ
��_���ܷtј���������0�;�ʤ���xܱ9��+�����B�&��I��yP����5����(�r)U�!����Y@i5x��_�/��ђ�
Q����;4"�i��ک7���uy�c����D�o���kA%�5a�x��;UBM�'"<� ��%�̔�T���< !ttu�?�3��p����YT���|�ɚ���|��D�dI��!�����E�C`�|1��.6`sE������FkO�!�W�^����S�#&{��gymb�����5��Y�������wŽ�͕��6�B.�WӤܺ1�F�����G�k�I.��{���9�ʄW�ù���t��Pt�u��x2��!����Z>UU����u�m�g��;é����!.����5�mx���L2�F���fi�(���|7MҥmI|�W\�x�w���;��{,b�5��V·PQ67��	��G;S6c�	���[��>�y�t�X�l���,��+� fzv��� �����������kff��6  K� �wU�a�jY�_�PMX0��g��p>�j��n7|��	EP�C�ߩ�0�%,ﲄ�����
���6�7Q ~�gk�@����5��bFj�W=��"�)�
B�u��r��j�A{8v��Smdl,X�[]����]w�@QGF��x��L�[Nr�v�R6Y�ѢjP)�g:"n�O7������u��@�	�Y�'������8�&F����
����&�%tS&䚏�xycg	�����E�n�|�[��E���C�m[�r���������U�MUG�s�����{��N˙�����&*f�� S�v�������\ 7�q9���p�Z���$�y���P��Z���pq��Eyf�V�N𵍛�먭�nG=q�-�t��vh��W먎�1����O�'�E�563 
�^JB�k�̍iϑL����kq��r,+�1�^7��T���21,3%"'B�)Y���oX�xciz0 ���&�/H����5SV�J�%��Ϳ�d������w��x?�"�wV�� �V8�H9��1�ͣ�g_�� Sx	&������]҅u�W�)@.Ξ�5�j���==��G(L�O�=nu�@'�y#999�%N��m�gl��������
iWO��#���� ������l�d��:[�B�K�0A�<"7����*���N#aw(��|'�cM�$>>%�CLB]�����E!S��{���;v��l��߿�DAQ`�5h,+��S/՞`��XW����kk'��O�88���~~f�l ��=��8՜A��Tv�/��'L�=V�n@�5I��r<SS��Z�౷��v���%�����o�������ʹ,�9<D�D3I$�Ny|�:񭜹z�*���eF�g�T�]>y'�n �����4:�M6K�۲�����s��<[ɞL�@XE�H˧�=^-�3��S3��6oa	�Z	��bbb,����ru�M�_������:�K�pr��nlh� ����n�c	���^Z*�9��Vlp��K���R��ŗl��g�9Rn� h���MgzS׏ �w��4x�ǀzv=����v�1n1�rg�yV~:^���y���M���M�mc��l�p>k��"����N�˙�R0���J9O0Ɍ���e�ӌ�2D�CwLQT
��CD�4��bl��
<-m���}�fҼ�hk�ov�5�-�n;�����Ņ�$<^����NM�p��~�HP�f�sՒ,fԞ>�:�u�1�:�ۣ���~���6J	�Ch�#�E��cV/���C��i��gc����6o`(�j$�sM}�%!��l�/hş�xA�%��F����i$�[�r���wGtV�&�d�����[���;&��_�b1خ�+��o��5@����5\<<�G�蛑3��t���q��)yyվ�p�]m�_�e��r�ӥ��q�ᅔU �hD�;t��`����V���	 1��X,J�<a�������O�=9�}zU�M~p'`,�N��)�ε�%�|��f��A3�� :d7t��)G�-�+#6	����>���cb�Q�}�����H�� ��T�(��*�& ;�iii��.�nGW���s뗙~��Á��g�r��,��1��X�e����6�(s��̄/_�D��t]��of��_hj�:L�n�Qh�R#��G�-X�� 5�bxѫr@�E��A����8����zujf�0;N�H�E������w���Pb�e���C�$���5냙�OLL���#���ױ<
E/�Q5��D.�ب�5�i�S��k8�.�d<w�5��@7�� :D{���m@������W�OUwRg�B�09I�⢩��u�����{�jB`�13y�L{ �S������T��_���:�a*�pt<�L��Ԇ�||j��q��`G��xQ��H��w|�]�S�A��:����yyUw��j ���7����~�Z�Y�����e򘆖V��"IQU���徝8Y�6��[��:�y�o��=Bb�W:��;��y_P�����ifg�]�G���vI��E9���AJ������>��$/'��\~�����x<k���(��!�Ϊ�#ׅ�@��H��6��i�w���ؾ������gk��.����Eޙo4,2n4�&t������jia�uLCU5�s�=ҾQ�#�pb-�=�@�{��v�r f���z�vJ��U�GDPK8�
o������@g}�EE�߇l��/^|~��^\�	,����*5����N4�>��vi3��*��G�_��X���� �h��Q�p��l^a``X���E�v�"������g���E'�Of��G��N%�h�����,�le:�o���-,,d}�3�#���FFF兠۱D!��f�5�3@��Vs��eI?��H����v��; %&͎5����S�48{�&˙���ًH(��ݚ�����|���L`�4��κ���s��@��\��s���K���=�w�Ė'���~[?<�a�zsH�Ð'�iLJ?t�)��������s���T%T��n����(��ϙ3 P-Ȫ0k}�bY�{�'~B������E0��?����W�#�+��B��So�v�=�	R�x|jj�����- G7���OO���^Ɏ��}��<��D&����}�2����$�-3�u��_�!w�Q,��ݹ���B�L�be!غ�{�L��G���E@&��&{��A��w?<�'s������z�^S[ww�wy���T�a��1[�����p����2/�;�Q��2��÷�}��C��-�G���O
��85�������졩d���)8�
(�@�_��:��W���x�۩�`!7���r��?o8���X�����&�_��Q��&Ss*��6�4,��_V��R�@�h?�$]ǚK:��ب^�V4�݉?^(=�6cf�%�|YU�/>5�o�ى�
�q\�	B|�:���m�f��m:ojGhC��Ԍ���tː�3���Y��w=
"��	���1&_~���{�i*�f�"9��b�.��CE�b���`����$�,�y��Gu���^�::8x���������&ج=�l��lsɗ"nj՟��]F�I__���F�Wn=����ɫ�C-�\�iK ��T%����͛� �8L�`�X�(O޾�U#6.�ߎ%%sP-?��������*N��݆���� ���ܟ�����s		!�փ��Kzܫ���1P̐�1i�e�����lkV+����w�D%�|�0111��E���ح�R����#T����`0��e�ſ~�89=ep���P66������v�w�($?�_��B,�k���;�ߔ�r�?�>VU�͜U�D���::�ƴ�s�v���ttU.��6���U���8?5��Rm�����J��J��\����=�=��*t.�V	��;;u~�k|��U��������I�g�y����˟g���~�:���y�}{����l_�s���6�Ѥ��T��h6�-�| ��or�qn��`0h����͡�4�ʜ��E���l2?���&����Ɉ`�O�|&�q�^[�G�]A��W�>�VB�F6��4&v���`��϶|�b
U��O�|U�K.,?�>^j�{)��}t��w��e��bs8�%��:ۻ���g>���w��o%��	?�k������=>l��Z�>n����r�#&���{g��~��_;�]Q��ͻ��P�f�4KQFaF�FLZ���%�Ʀײ�/ZL�]頏�2���ʍ���po�ǂ�XB��t-�@K��:�
�ji1W:� W�)c�������o���/*����)-5y���~�7�-�ԇ><S9��:�59��uye{���{za
o"��u����s�R�9���3W�n1����i݂��ek_�|�p�
�O%����9������>�(&���f8���p٢AʖQ9�y�Q�2&;f4���N	}�w��P^W�es)�5��l]U*S�q�ƺ�~:�S�������>2���z�ǜGk#��fk8����1����X���q��I�xߛ�{�Z����c��[��o�t྽
XS��4}S^�m�T���pLy��fR('a� ��x A��pB��1�h�ZpO�ږ^��T��o�)a�1��uwǬ����E�.Cx�0B��#5���I%/8JV��t\.%$;�ҷ�e��}@@߅�>�P*Q0��� PK   k?�X�F��^ ~% /   images/60a08d3b-0b7f-410d-b1ad-60796781a205.png�c�&A�-<m��m۶{ښ�m۶msڶu����m�x�s���o�Q���b�{�ZU�"�%`q`��� �KL�������!��L.oG�{�8+K�����;��臔��o���vSU׫�Z����e�gT���Q�J�(��	���z�1��FW�l�hYWe
/��%����lF�$�U�QV�?~���[O�[�Q���O�3ƚ���=��3��̣x�tpo��)����B0��儁�B0T ��� �� �����BB��J�������R2	@&W����?��Z�� �c!+
K-�YQx��?8���dg��	����?8L��g��������?8X`�4'�L�<��	���?81  ?�3����o� ?]t���3 ��%[�(�°�� ���_����_����_����_�������{{�gp܉y�%i��y������s��Ԭ�\u����\c-���{u{��礡�*}�K�M���}���tEA�{����=������`��]����c�VC���^��^.�]z1���6�n[k�Ս�`�է�S"ѻ��m�nZ���(I����$�w�Nz�zNDn�����>{c�	�&�띕�l'�cE$�`��Kڕ�Y�L�)�ܭ��!��BD�G��ٙ�Y�k���6%�턕���\�q�J|��F�/���]:%߅�i�4�pb߮\��|��=��@Ҋ~H�:�O�� �_������>�\h�u���#����c��kK���!�㾮~��@[\�5>x�$T�0���۹���3.�������o��}��u�S5����G��o�Џ�8����H^�H�wc���q�9L;�i��q��@g�s�%T��{mjq�����V�f��YKs� S(�t{B�nA��B4�Jݺ�|�m!Wss;��� K���JK���&jY	Cv[����E#�((��N#�6ٺF٘R�h��a�QCh����Fng�y�<\�����ե�@�*�l�-����7�J�.�>;���4uX��q�bK±������ �(W��,ʳ2Ҹ�ЈJy^�������F�z���5��vT���N7���Ca�*���Т��&@&��J���xc�`4>��8�ĵ�|�M���}t}�+�A���_M ���(���t.������m��e��d��׈�<��}��ݘI^��ʸ�
�1U3����,��4���B�c��y�gZ�y5k�<�?���d��`����ުB�89�5ٚ;��j��j�IҪ㩶*��]�,�S���?y�H�,���9n�����o�a�]�,��vm�[�k�ɡ�4.�A�c,��Yj�=�`9�����Jk|\v3�2;�d3�1��s�V��;��f���`���5����4��A�J���{�ӿFHQ�:i��m}a����������7�^ɔv�=m���,s�ai�2��<��-��Ai���~����La���D��������� h̹��&:���
�G�x�5^rv5�[�Z�0���/g> }�kh��V֌ס?[��;
/�B]-�[׫���gwa�<��1Tmz*F5�0߃�a��tዣfZ�q�ԉ8�T�u�:xk^�/c,f\>T`�����j�_3��RaK�r*�����+
�3�������W��F%,�i�� K�I�$���#O�T&:�F�|]��s�s���z���}���F�u7�HN|8�<Rz�=>ɚ%X��m�rN1��WP`( �9BD���ҥ	��X�8�d`��j;T �=n
s�w�ҙ!�� �]�<�J�۠�^�0ɡ�K%=��! �!��q3��M$�F�7<��"�"g8��{X@��)�5�ꤘ%2X9+1=�H�"w)�$��;�X+��Xc�)j=���S9H�^���bɛ�7YsX��s�$,s4�Ya�����l��l�r�d��!�tb����T̝��I~
��"��gV;]o%jU° ]e��,�'��I�'P��L�2ѧ�d����ݍcx�)��ڦ�k���6�Ü�����Fw�}Kg�@w��F��c�af��Fk2��j�W��0"�+��M���y��ƭA����_ޱ�ҿ���<�*=��&@�Kh�6�i*g����n��F@}����e��D�lb�g�u1�j���Nl�Y�bL���'�I��O��q��0��8��Ũ��N{�c��kw���2���b���j�����پ@ޡ֪:1R5��]����.F�L�7�?�E@����:��5�"��w��"�Atj�}���}��l%?���/m���L#wK���i}��k�������U��`(i�~�"��;:>�i.�<�QO��� ���������M��{�)��������=��)��w�T����#�Z��Tt��Lq��JZ�����:_uVB�;k�͇V�@	=���5��߃A|��*h�z5�PH\��A]�Q��\��c�v���X��Z詞i�C��i�v�G��5��<[�J#=ZhjvcFF���V��̣�����گ�~!��]MKo���ua��6�'��󸑈q#l�jM�y�`����8Q[�{�r���#]����j��0�ps5�̯&py�y���=��-��$y�نL��+Q<��Ů�@�W���qM)��^OX�����K�Q�����2�ʇ1�X�j]3s�:5,,�����r�'-fmA��S,��Ns�/ؘ�_�N��M����N
s�d�Eᑉ�������@�hڍ�h�)w�����leڵ�I�6d/Ժ\pI3�JULcL؟j�t-�̠��}tt�/�cia�ɣ�u�����?zq m0����b;s�3僗,i�|�I����8���,�d2Ƿ��\�Hqc
h�a)��]OA}ˮ�Ȣ��D��aD7�Iחu�jx�� ��Ϥ|1Ab��1l�������c'�]�;���N�+Z1�d�M0�cN�g�2�ʸ�Xͨ����J}�[�8z�5���:���vD�f���Xj��uml���ű�{<�����y�c-w��=�"<���U��M5��-�j���V[!D�9#<�=��n
Y������_W�βV�u7�Q6��������y��u�נq��ş��VTƐ!\F)CG�}��R*j�0��9�=�tU�j]�0N3����@����Dܱ�4q�-<�/*\��9���p�W|���	��L���^Ҧ�/$g��RU�������b�����n#u��6'h\�c��������/W�-���[S�T����=��J�[��g���IJmL��������J|筄>�*��C������=�$�}e�����A���l3D/���pm�2�@�˒\�(��d�o���W�����TY!���K!2����i8��V�?�'�f�.����&���������J�̙MF��Y�r��U�I
�S����đ$;xOr?/3����a�$! r%�X����]|����7Njw���(|,R��i�-@�u�༌��h��'�����%mF6+�&��S:8��ư*���a0^��~X�݌����κ�'&��G1�c-c@:��NT~,&M����?x�!-��\ә�u�e̲J�8&Rt��p`��8Q�b�n]�\qU-Id�[duv��V^5�jU�֎zdC%u��;��%��������$c�`U˗֧=�0���j����Ȍ�Oc�@ ��bf<@�Dg����.���W{%��0�`q���4%7	��RO�`i��Aj�l�$���%B� �-X�)���)���"��c�^c�u㊣�"
0�UF�	-ۆ���gm���֛[�niߥ�������H4�
U�& -�����p�Fef^&W�כHZ����N��$U�N�%[�y���]6R߆�r��N��rp�1>�o�����P�����O�2?V�����9Bu�˜,�;��Q��<&���/
�W�0սH���]�V2"�� �jkl� ���-{yY�I�!��񹪠�l5�X};ʈ#Ixqh�]��{����K���Ŀ�VM��ik�)�Wx$i!�l��`���yx�+I<M"ΔX�!:�=����ь+;/Pθd}v$�;Jٓ���^5CS�D��%U �����rj��k�ь�H������7@.^��N��x[��3������у�n�=��H���>���򣗿��ǿՆ3=�]�t�5�v�Ց~�HZ�(Qe��<+eY��~F��F$�b��y���^X���|��;7�XR���h߭["���P��0eA��f|:QɎo�U��o�
�����Bq�\u�>�j

�v_?���T��4X�p������������jVN��E5�>�%��g�Wm8L��N70�j`���}��.���;�(ԉe��5�^�)��	B��6�Nۍ�;�D)�<n����z�^��"�`� ��I^M��q�'�����T�ixq�'�\f�9n�0�ݔHE��Dμ,9�LBy�F	������,��a*��cMM�ʖ��О����Me�F�����8�PO�NQ{�A]>_,�����q�1б9��=��M$c������y��yX�K�XPl5g[����}C'�}�z�;��R��D��b4��B(��C���1!:�ٞ<RL�b�+ �����g�3��
��f?�W�燈
����:z�[}�(�O#K�T�I��^����5#t�	�i�U�y��he^���\t4�P�����f���qa�Aꊵ�%���>�ߦn_4�%|�e�-YLH�@e�h�,A�3z�=�`��eÿ7��P�+��EOڦ��V����i�Θƕ����p�{�eB�?��J���A�^\hq�����Ε�E���Ȣk��NYi��͇�b�舼HB��N"�Ob������t�}/V��+7�R������l ��"F\�B���JU��*���r�W㎑��T�D�P7�M;Li���H�	 ��F�nlL����Җ��t�$,������(f)� :�$!�YCceE��
��!m#1�:��2�q��"6���-�	Tʒ��N�.��7����J���a�yC�+ ��$�U�Bzϟ< 46�
ߏ� �Iw�����ǃI�b���_�m����=���o�Al�F$7����ܐP�N�*�yc:��w�������=�Ut��L����&f�B:?����U�B����?<����RMo�t0㨑���n�w���hB�1E�)�>��a�8�:B���Bm`8~>�?�^�)���(�0��������r��k����S���NW��K����~?/�o�M%V��~��N6l��y}�|I2�ٶ녤�)��݁z!8f��8��`��HG����+���C��0Ɵ�%P�{�A	zWI���q�xG�����$�Z�C(1�E��>T����+�L=�3�$:�ZF��yq�%�pQ�^Vm�"�D���t�����&(^�m�"���4\XⓉ�F�i���.V��(�����%�?T��ww�gc;%�`�w�/��3S.�����*R����a��a�_�r[��x���#OX�p����t��v�:4���u��W0�F��IU�^�rwج)N��4��C��m+�Z��U���C`�GZ�N^2�D3�)@﨧 �m(	ˬ.%�&�^7"�V�9���¦�����C?��f<���1|w���@Z��Sv�
(F�%DN�䒬��j�4�6M�ﱐ��տ�����M8��d�����W�
3�_�"M��1w/�� y8��J����aq�HQTq��ɓ�H��g�¡�͉�Oǚg<8��Y����L�#�B�P�(�����DUh�k;��4%ҳ%� 	ó��M�� u;���G/N�1������?� %;��J��c��;YK���=�J��p͛��!��V�~<�*[�O�����
_��=H����/��{2��$5�yd�Qz��
y��5Q&n�N�ΰ���Bc�����d��V~@�����>�|����2V�k������*#1�(��K�_���v��ԛBʱG��{����2&��z�������oz��qf�҄��P,�`��1��Gxt��Q*��?�J��*־�B��S L"��I|9y6N9�������[��78����@pD�.�-�
)ؙ^��i1A�%�ܧx|\*���3~�v�L���>�!B��G (=$E,h��~~��dD�9Q�2���D�� �;L���nYR�Md3�D�#+8�n,7F:(�Y��I��!�˝R3����ϓ�r������j�����r�?L��梵"�ˌ4b�聹���I Z�1��H�պ��eYiY{��{��h.p;�����ﷃ��T=8FQ''a&�n�e0�,Ck���b�[B��c�ם��췭�p=�.Zs�O�t0��,<�mJG�>~�|�5k"5[b�X�D��M/tR�Ħ\�Wb"��L��o�d^Jv'��MJ9���V��s?�����u�Q�6@�H�����lL>�ȶ�q����j0�S;̻a�t��M�7Y�[`p�|�Sv~W%x������J�����5��ZrIƋ-��0���S9&e�y<O���l��D>���`�JM�r�2��_���kVP��	^���M��ى�a{�nv�s#|��=ad�Q876�%P*u��������!g;Cw|��ؖ|�ļy���u���Tʈ�4�X��=)vϖ�Ռc 2Ѝ��L��y,)�qG<�A�����!�D~o�8����#��|�?,1
��ei\!&l4va�P�a���r�󁲨�D��'}Y�߿����r��S\�ӝ���r��H��:�Rz�4�t��?����w��f�J�z���ō��|�ZÓ�^�����i�6!?�BmI�d#@n.��n7�x��W��~�10)@q�ݣ��a2�H���n	�������-6�hM9�tC2%�dR��sh)2K�M1��;���QXZ��~uYۏ �������C��='�q�I�Њ,���J.= �] �Ϗ޽�8:BT%�X	R�ic����!�R��t,��R�y�a���]��T{��g#j����~��e?;�Ni���a�8��`E�E�����G�)��k��{s��ٕ�����~�J'���0��4;y*c�ջ�_~��S8�D���/b��x���R�
='k�k �9W@��L�865���(_�3'������$�0�����	��,<	̆����N�q$k2Z�0ngA�U��l|��MnεR�ı�f36�Y17�
S�����9�n���Tz6#0�-�}(�i�jjH��ˉ�K^-�<QQ-�R���D���VLH�JW�DN���
�O���?Z�U9<��l�v�W�+6%����`�ֆ��[�U����X�^XW1z��Ɖ�D������ ��dJ�y���ƱC٫u�0�������_�I:u�1}gxC�����]n�\"@ɶ��SN�UQ^7��fn^jG1s��}��*&b�	��כ!xt��l�Ê��3�� ����6sK�ң-p�z�ч�H;>律�eZ򸔶Y�֌\���e7�����y��b�����t=�u8~�������X��0fYT����Ѫ�W���������@���` ��,s�a�V�ftR?�q������̞?�{H`Ø2�n�9������Z7T�}IS�{H��F���n��,��~|U,����@�棊k�(jϵ#,@��*~�ք4�8 ��T�MZ�2��f!.�A� "0ه�NR�~��/&_� �i\x�K���
yV8H�2���ޯ����b��߽+����aXĳ���cT0p�����nSIJ7nDx��W��M�]s��v�ؒ�.���G�N�����,U!��Yss�ǭӖ�D��-�4�v]*'�UMĞ�^�o���4h��+��^�Nn��^g�� i�˭�sc)=�}�
��	��Q��L��m�@?��Y8=������E������%������y���y;��<cM��n���(�QL�1F��K&~��6ؙ��!D'����tE�9&�4dOיYz}������_;��ӛ�J;���naj����8� �V�a�����u��?dA�'Ù�\�uX�>]�9��Ű��gc�}ZI]�(�(d��F��{��']i}�MB#q�����-�,��Y�2�]F*e�B��(���j��L�9�Dv�U3��[�B���l���*;b�b���k����ʂm�� ���0!�.Z��f���?���z������%�Y,��\�A�1yt���fo�F�#+E���c�I���y,�0�F�Q\��o�|�E2�sH?�|٠���p� ��SO�9�{"�х,�;{�·��E��ęK��%����kT�JU�ݏ�u�Mg}o�}#C�v�_��_�3��&��_�������Q��n�x!�+ӟ�p��u|	?���n�q�z_M�z���q�Ǎ����7�"���}]gz���5��TRQ.Ө=��י6�s ��2����8��Ke���g��2 ՜Oz�9#����;�ҫ���ޗ��%
Y�-\��A4����T[��)OMR?���>z���f��c�;� �t���H6#,T�/T�7�o8�]�y����t����8b>x4�dQ�ɰ�h�+�Zrj}�/�D�`L7�H���+aj��A�j�5w5��P1���E���-9x_#e��k6�3�!����n�tD�{܁����~�ݍ&���3��q�\?��^�wm������(�z�Q���
��ד�M�ש!��� �/A�ƾ�ɤ&~����C�	�(3�̪I��%s���4.�� ��$\3&�)Z��F�8HY�l�^4��13���5���R}]���"���/�Њ���Z<�yw�K�hHPy��2�HN�\�ш��[�:�>ȵҏȼ��Ԫ:�L�u$�����E�S�]h ��51D�{��#W)�Vqא��{S�L[_z����!�*éV�B9{z����4|C������,�'�����&���Iy�'CZ�۵n��&�Z��*���sQ�0Kʽ�&�Ï^\�hVp;����Q�ԅ!<�[�++H�ߒ��{�Z����%�ȟ�m���gI\c��Ӹw�����*h*�_'�'��N���d����T�@fm	�c�l�
i��D��$PoG�)2�\С
X�D�PZ��j��l�*
2�F<�ͩQy��Y'�E9LW��P�eN��WL�0{\�i����C����lB���̻<��	�۵l�����X��0]�0����0����CG�R�Cw%v��c)P�=�ݻ�p7H}�3���_`/��/�<R?ag�	�hG"78��?���o%퇋.��>5���o�	����S~1G�9!��;K	��;F8���B84�b K�q�by��ie4 �����'5�&6��õx��^��Ȥ�$H�);f,߯��%�q�׷G2�\Ɏ���f	SB����m:m�j``��S���]E'8�N���l���>fK�LR��iŎM�a˓(�e�ŀ�y���΁���c���s~N�g���E�Rʋ��/n\�LDEc�_��v���$�Q ��P��YI���	�]���`�LF�Os�X_��[�u}�NE�ϕ����ߺ.΀�0@��A������ΟW�tD��tA74y�W��+��f�-\ѽS��+oD��	��z˹�ʙ�<���~��7����-a�z�(�2�z�;��v�&F��߅�~m�K[ʳ����2�ɵd��R�系y�L~��ܩ~� aN[T�J�����vk����<Z��L�͸��ͳ@��&9��WR.�P^���E���@Q����̓bt���'�
�k0�u�o!ի������!���g�u�������ym],qV�����UU�������z?�Vi�8<`��N֢��D�I��,��k��B����t/���^�I���\G�h(�(y~o�d�Z����$�]�1�1�x�@�9K�Ҥ#]A�e�@1E�Q3�pd��t��'y��.��&]��gS��~:v�j"@��"'~��Ŗ^s���.�j�!}m���M��`<�_�k@�N�Cj��)m�m#�{��w��V�q�(w��)�3ԉ����G��l@ѭ2��ů�0�@i�����
��ʧ�.��!ݓ򸰅�<������.9%!��k����Ga|иQr,|���z*d�j�әj"!�Id9Y����j��܌��e2�PN����	lQ�.[:ԫ�_RX�R:���D�yS���2�N��C�&���%�!�n�6�>�}o��FiK�-+�A��]`2���=pdE��5�����)��2z��HJf�;�J閪��.���/���t�O�H�b��9��BE�G��������L4����]�}�W�$uldU0�?��z���s��������J
�َ42w_�K����*��#K��W���u�{�V���t��o5m�����r~o��00	�p���g�ɤ�� �ypn�L�/��R2[s�'m/��Ǒ����f\-���>Dp�-��R��.b�>����uc+�PѴ�1dܙ\6��k'��^�O�Y2�V�gT��Ǒ�6��z�]Z�7���\&/`܄��H�I��m�]*��������1YNzMl��s����6V��~�:5;�\�����q3��A2���;��/��̰#У1I P��(�[��?����b�Hçc�dUs���n�:,�㟎.]>UqK�t+�$���Ё'��E2
3k!']�~��u�gz��������k;�cg�㧩����UҞ[��[��\S�]�p�[�<�����杠�W�b%	#�	������pN���	\�4z|I��~�ْ���f6�$j���Ƹ|T����:9�]���c^b�w?�t�O�,��@�����/ɝ�uC�}N��O��&2��Ժ�8F�G�Ȝf
�^r
m����aD��'�Xq�+������ΰ���� h���Ǽ)�n���X\�{��@�?6���+��<��c25}��^�a	!zR���^����F�B��BNnв�~����������K1?kا/\7>@pN(��ĵs�����Y\�n��_DaA�]Rኹ}�	�<�YidT3��)�9i.�ȇ��1R!焹A�`%�lNN��
�p��@eÐ��:�b�N�K�v��#�����#�^��>��I��ɭ�Z�$ZR�<�2n݋�����T�dC�������$TA�,)eu��dv��|�jX=1K�73��J��1?�B��qC]Z�sh�`�33e�j,Vcu)͘�ei\�N�]���W��o}��C��d�Ii��{�[���C��x�A����|d�Ncj�u����	M�1��W�%��d�������a�����<!��i�F�Ⱦс�ʤ�d�����q�T���q�Ob�1�^�5i3w	��Fg�t��
M�����d�������B���"<Ѷ	�;5S=����������0�۹	��{q)�x�g���]=(޽����>� ҵ/r�aD���0m�'R+�wy��m7�>;�ۉcƁ���p��6&R4և�kk_��s�����a���1w@Qz�,q�!������<Ϲ��>"��T�`���(1�!̒�H���>,��y��4?$�ƽ�FR˛:�r؍2�t�>�:�]�.'x�:�F���sch��xYJ�������\� ��1��Nx%�f��*��%�P��Z�П��Uμx-g�����m�a�
S�L@c�;��P�-2[Y�l��P�����D��#�	��]�������H��+��F[Z��W���p2����G���=2���u�v���q��cx��M$	�%aT�z�ǵte���Ɩ	{����/(B��:_(�Ú����3�\$���Of(�#�\���/;P[�-U���ނ���n|�f�+;!�
�#��-���	��g���X,��E�� 7��ҙ���0UV�C��H��W
Qn�D%�_$d=Z�*/��<�̽�BqpC0��@C���׿��}D"�+gNH�Rʊ���a�;�'[�����������//׾� ۼT�Lk���G�Mfd��٫�D���B�Nx{��T.����JUc,�7�*;�����J��9��y���l�;�6��2!�(�^I����ņ�v?U~7��㙙�Z�V3W�k��o�ȹӧ��^#1�"�<�?\a��>æ��� ��U�	�P(�����{�aQzϱ�q�pV?�o���$\��e:���Q;��iA��0Ҷ-L��E�
	�?k�d�uk����l������f�,��ef��v�%n��i�Dbn�`�G ޹{V����/^2#:��0Hq��$�I	�� [9d�R�ʀ�e#��o��v�A�x:a���M��i��Y{�jY	)0�R-�W�����Z��ętr\��D �~����A���F�d����̍��� υaｏ[�F�ҷ���}���p�r'x,��q��^ꮊ���������Ma70�`���}�8��	:A�$��V��y�>��lWj9��䟌Z�p��PI9��_��#�$���cb�1&��s(��,��� ��]ךX�$�|��l!�� ��U0�,u��ƚK7�a(�ͪ��iO\IjH�]��z�C
�1���3p�JsN�qf�<��E����D��v̄G��Q��#��?�L��Z`6{�ZJ���D�̫����QOz{�u�� ����w:����y��&��Gi�]OT������l�h,��^��cǫ5�ݱ%V.�I�5��ɳ$��Lx�1�N(����N  p���"i����s��&�i/�(vu�����c����灴/4z��=F��Ԯ�1:b���������q����d�Pσ>_��N$8x����pg�x�����b
�tgޅ�ִ�8�ck�R��Y����{$}ؓ�\���%�L��fS����$�Ql"M��_�j���^��ik���}��Q��Ĩ�~��8T�?��a�
��6��'J�/L���=X��s���oQ�����I�õ��2��~��'h�;Kn��0f����LU^S��F9g#�Y�J	�$�
��o0K��v��W���?fp���񧧖�"�~�����6տ�!�Nl4R�Wc�i,BF��J�#2�i�<�f'�2X�t9o����ܿ�Vr_��+�ׇ�]�6���|������^�D�73Q�6�]u�'�����Sa*�O=�;Ҍ�hӊ��'��Ǌ���l���E���N��'ֳ�?�P���b�r�x���<����?F񼶋�P��F f����(5��f�~Z</l��%�~t؏�=LVpJ��_أ�(4���
�'`�k����W��.H��󽍊p�ey��ҕ��G�0�2gl������3I%��fN�=eQ]����;�P��� ��W㏃����&`��t��Ҭ���{2��!&1�6�C=���Q��M���b������\��?�|�1�ch7D<+��#XI�N
ժ���OY>��$3��5��{q���Ƨ�?�Fy=��Â$�>��LFtФٽdI�9�G�h�zŦ&K���P����@/�{q�;
~T��J���럅p7��E5b��)Ak�,(S��*�3�@�N�·��#���1�[��W�)��L'�_R�z���(�����:.�q����4��e�9Y��双��4ZH��]�s
�DNR>�<R��GT�Z�n�y����v/I9������!�~��{��q��T>wE�[��"��i�ˀw�|��O���*�����3Ξ�nV�c��1`fp�o���zu�d6�@�2w��,7tS��o�#JO�����JA �T~#C��}F�
&��xӼ�f���๣�x�p�,����.���%��O/���������}g7�0z)l���V����@�W����5��@�L<�@ "Γ�4��<�wVU7:�����1����v�N4E6��6�=,#ϋ���-X��*���y?����?��8=Ͱ`A*:�.wtc#�@:N/A�3�:��ך�l�됒F�Lv��Ką�7����M�9��w�}��*�����F�9��@��y�#s��|�a 5�/���={	�7���}�O.���H�]�IA�?r�{r<'F����+������+5�&�0~屻�9Ͱ����q����́�U+�(��3]첌�#̏0�H{���iI#��l����#�KZI��>Z���6����VaK5�j<�3��\��JC���y�h�-~S�׃���13�\�na��gĘ���GI0��<��ޘi����`s����G'e�	a��BX�2��xp�Q�Vb��/d5� �%� �5�X�<��]Oea�C���0�YKA4A�Qk���´{?�mn�L�`�zQ�em��Y�-�ʹ2Z�P%Rj�E���Z�7	a?N�ӛ��k��R�����}Ok�9`59�M�:�wK���z|�&�ZթF�)EP����k�{V5��Q��P�m�2)����fy�А1�T��(�'�&;w���!����/�}D�n��q�jY����&��?�6�5ڎۤ�=��7���������h,�j�zYqH��ն�m&K�۷{`�]�];���s�NA�m��O��Ф��v,��\���~)%^��G^��Wv�:�8!v���7`x9�Х�_nߍ��i���c�w�,m3��ce˃5��0^,R~ݍ�0ɌLv��nȽ��5�si�|��/�Y�.�
F<u%���_��O���^B��p9�z�O=���f&�*��搬��ߟoM!�hk�����NH�������>�VM�����9������m|�����V�.�|�썯f�=�Z�Q�H~2��%C�ɵm�7_���Q��E��&�|wC�[w��x3��78��NeV�o��UT<����y�� F���(o��}���Y�� ����G���yϥl6F�&����[���~�}�����)��4��ɲݦ�܀�������y���-�(䛞U�6�A[9��,�_��ѹat�����Ć���~���&#:_��5��ו����~���|O�O#3WJ��'��Ǥ�~���������z��M��^�� J�C㧷"'DXn�͙����D�⃘�`c�|[t�鮢����W��vqF4ks�N�xp�4 �v^6�x�4P8��R�	Ğ�d
��<� �㾌�~Э��N��J�˚�������߆;�������)���ۥ�3*I���f��D1���~SHB���m�����rW��f9I���^�E�ٺI��L*�-1͹����h?	&�j�����p������U�K��Nx�o�Hc\u"e�+�Q8���bՌ����WbA]J�T[bl��؝��V��Cc�8��i�Jb��e���D��ө9�Vrѯ.��N3X{�{���5C��Hu<g!�ځ;,���n�_yՔ_�|ٺ%K����ݝ�D`�Zpj�"�d�3Ĳ�Q����}�K��z�
�d��@>�x(���/]_�3kf�M�Yʿ�'�v,Ֆ�0n���fA|'�m'!7o֬���"�	��Ce����q���Wt݃��D6�ZT<��P���ƺJڈ�:I;ѿ$$���	�Z0HƜg#�h@z�ê�9u>yX����݃�X���ĉ��z����i��?}h�����%���!�?����n}�L��em�6���9*�[�h�r2�.ES�e��i�������������àu)H���{�{bN��J�{���I�W�ڄ�Ԛ=�W0�V���2#�9^��5j���ՎbWl�^̡p��;_�F�.ݽ�C�Wg�������<�"��6�W7��7mf`�4�����+/#p��N�Ws��;�����C7��F*ޓB!�{�{+�Q ��U�s��}�zԌ�d�nE'��Up+z,�8|,9�����~'��j �υ��ߨ+šѺO8��㏕!j��H��y��Da�I��ղ4�O�ⰷJU�6?���YC]�*��rm�P�դZ���-�8mA���9����Q�����N�,�����M��)�,1J����枘����ж�;Y<A�p�>�d��kñr���X%9�X#�9�:�� ��Y�����A�l�V=-�1�Lu9#����j�̜�Ҥ�	I�Z�E&>���2қ��g W��	��E����`(�7�����ǂԂ���2
ء!` �������Rg��X��Apaj���,�3t�Ugi�(�%0����b�L�����lXB2�{�E�F���V@���Ʃ���s�~9^v���ge��n����GF3X,�x�EW`!�qpq�a�_e&3y��`�a�9K<G9�O��\[�O��aq�jwQ�)t���''���\�����ҳݒ1��K����2�t��7�soIݵ<��q����f0n��DU?;�;`1Ʀ
��g6D�_#)fCX�31+�HHژ�r$sOb�ѻ�����m��M��Ν;�O,�<~�Ġ���	���<5�,��M/G+�0���x\~�Y8f�z\w�'��El���o��.�@¶߾�N�x�͈<_�Lz�׬�/]y���-v�����0���H(>l����g���߾K��{���Uo��~���}�������f���fg���g8b�4�t���ވ�}�.lX�
�����7�J��8���YZ��G�YY)��v�}�9ߺ�Hl\�F8�KԘ�ל�F�ĺ�	��z�3:%�W����sx��'�<z0Щ��3��سg�<��b�K	�?��3��O��r�/lj�|�w>���~�<x��_�>uí8ԏa��F���SO�����k�N\����ݹC�x��1|>�v�ǿ�8����g��Y���o����:x���?�^����]�ƞ�v���x��'������~��n�ޔ�/s}��'�+���|�2���G��+O���	�^=�����{��U�i��9gzӨK�,ɽ�ml�������M���@BB�	l�lI�}7��f� B�&@��fc�1ƽ7Y��FҌ���޽�3b������y����ɚ3g~����]�Q�%�|^H�:-�#��!�Z��iHY��|S�To���y_��kV���Ϡ�|���-��*���d�t�}������P5r����o�p'��Fp��&,�8n��;��"X�V�Y^f����
+�sE���kم�l_Y��D�Xli"L�r�wz��Lf���z&����.Z����ǘ��K:ގ�_�(֝��qB'��!ӌza�NW��Y��f��� �����RZ�#����t�N&+LZNq�^��lIt������IC�t�%jE{L�Z:9�he�fN��o�*������=�����ɡ"r�:�]q%��Sd����i^X�Y�. w钠":\�ԄeoN�2�a��FK��:�"�5R��ENm����w	�T����MB5���J�0�a<8��NL���5h���Lc�v	k��������xRsKt��O�������{o����'��cu�4z��.����*q����+��Ϲqr��f*Z�!Δ�r)T�,x�,�ZC�Q��᪋a��&<����`�^Y���}��b�E����x�g��<,��?^�E�F,9"ĸhu�X�V�F0v�X̘yrE���������CRЙ�r�5W���A������o��=,r�"���/?�)jk��=���}ｽ3�L�?����6���y`A�&G�=����i�����t2�\6�sfMGu�BV��� �UB����E����<�9�`�G����G�p�t���P�ů�%nj���p:��To�؃'NI�������{'�,�@��ϼ�
�{���%�nU	%��$<��9�g��w�.��M���CG� Mݿ�1��n�����D���o��;�އ�H�eᒕ��߽����ؾu��%�[Z�Ʈݻ�Υ��g��\[�*]�ȽG�1j�$�i��1�|��N����כ"��톷���
���� �PTP0�r��T�u՜so���V�?����S?�8[�?�E}ʆ�=���X�\R��)�CX��J�"zu����q��Z���X%��PM^�[��|� �N�=�8�b��s����#�)ƜN�8��y�Q��BN��1���;��P��0�����r�7�d�H���c���D
W��7�n����vyd���uK�]fMU�tU�QTUE��=tQ70f���Ǣ�~�t�������Q��#�lS���5|&�'�d��ԩ��#􈎙u0���q�uW!f��r ?��	�g�j�<�|���gYp�RN!���$�kw��r�A�<�č�+^��~9�~��h�D�%j���f>�l"&�,<��ŝ<Cp���~��"�����`�d��ak>�tہ�i��@�W�����w��T�Ġg�oVY��Y����a��6�����4ԁ� �x��H���C1Є��3�D�,9�QH'PC���BPI!ֶ�ZW���&���?�'�i��q���+q麵B�ڲy3�}�iq:T��(J���YsQ�F,�����6�Cs+���ro���c$]��������������
���/Ha�`�~����F��Ef5�������:�#Cq��g��ޝ`�����]����:�t���K2>,�+��h�c���=R�9%s-u��%0��� 8\8)���9�o�-{�[�)w�� �:���nq���#���q�4lH�FN���e�N��#�Ƣ������e���K��0�k�\xf����}-�P�������]*|�d2!k��σH�B^Kmu56���=�b�h�	�b��k��o߆ζ<��C��D�QUE{{���3��4�4�5��5� �ʨ �p�{�R=D������\���Nq6��T�MY�7�J�|A����P�Q�_pyLmjxkż����k֞��Ϡ�|���-��*�N���?l?zo��Y�!��zK�+fs�`�;���|n�kn���j4����j-[:k��2f	�D�P�����C�ЗH	���s�Q�bV�D�����i�a���X]���@	�]@T��5+q��%�z�d��;����=���^x4�O�(����.��oF�����F`a~ȃ��n&��������U~��yg���ƬY�����DNC�s (����fxCQĒi<vB$n���g'�WUY���zTE�bG�`���$�Qw?�h�P�/p�go������޴����>�ߝÂu�D���`�)r�%?������g���G�y�Rg�t��e�EX�4P�fQH��m5���V�iN2>�tb n�&8E(�gWM�huʹ8���rdCb��0z�kP=$s%���D�$5:���Jhޠ���`@K6JYG+h*3k����.���^�4�D?����G���y�V֣�e:*Z��Q�5dţ�+�*�ETX�(��'Ӌ�/�Mc���G��]�v	����E˗aݚ���<���F<������(�E��Be��f�Ask�e�~�������e(>"�ѓ'��;E�84��U�_�/}�&�����6���,����ʛǎ����;L?�����7���>�u���������1S-���2bB3D6�r���TUTI����$뜒��B����]Hm,^2��%N��ӝ07�c���� ݽ����vV
tZ�a��"Q(b UĖ�w�`['t�����C
��;��E��*�ٗ6���^�P.C����V�D����p.[��7OX���r�<*�kO$q�T;^xe��P,��nw[>u�5���[����V��&�c�0H���� �9�N#?Ǽ���]��G��@�1H*s~�Gr>�O�@F���s%�**`�*`��h�r�k�h��{}��Ew�ݡ�A���O=[�?���JM���'�����T
�jd�}��K�g�#㶐AX/b|ԏ�c�x�4z�@�񅉬i�?����m�{������-�h�!��~B?hN3b���Ch���%�=�9���HX��Un_��J,��"K��!<��O�����L�D[�z��?w&r�aѲ����j9A!���fRq�vu">4 ����K��}��ޔ��NP^�Lw�S�AT�/�����}�>�GPUY#�+���9Wv�-c+q���w��T����ر{v��/�h���?w:���PUFNxq~��;���z�� b�"�a�YϺ�ɂnG*G�!-e�nV|����ď�ϸM:��ؤi5Ṭ��l�|^:s��g���F��Lhvn3��WCe��]�y��r7L��׉ML8u��,r�o����ny`��P���M���p�=I!_U7�G��钊\I!�	��r	��i��Bƣ婧���1���a)^�ťO؛��j�P�) j�P�C�Ƶ�\���F<�أؽs��a���X�p!���غy6<��X���_	���'N��hU�܏�r�O!���UȽ��݅;w���#�rzk׬��?�iT��������}�"����6\0w.����=��/����F\�n�0�����@�J"7�֜rB��x=�*k����rK�x��4��*����u>A��,F�>�L�h���X� G䪿?&��ށ~q�㪪�ik��&�"Y��O����p�T'2Y]d��zfA_�`>txꅗ��/!�+���4k����^(߆fC$F6VWaά�Ҡ�9�]�rG�F��v큩�DV��}1������m�����ىcGc0F�?0D�ANd2H�����I�M]c����׏�2���0<?�44�#*:Q1�?3�����
'�M�[/��a���-��wnX��38~�>�c\���c\�ѧ<ؗ\p��Ï���)yƑ���`f�b#�g4(uV���O�����eB�Q]q� F2C�4:9I��s2��A�]'�x:�I�"�<xLǞ��LN��vl 5I�j�z1&����$ƅ]H'�8x�(zf�a���Q�,_�5+�BQ�7�AHX������9�be'�Ab�#�!�Mr����,���THΨ�S�|a����EK�p����O�76,.pt��7g.�/Y�1uaT�m�+�c�y}�Vlݶ]N'����s8���(i��Ǔ��珠e�j��Z&�(�8�;0�p�l�eF�ݬ�;Mg���P���T!��A��!�PB1�Afd�)�7Qu�z.+���v%�ȑyP�$��q�#����J���g�L�p�{�tS&�ݭ�I3�E�P`�ғ��z�FQU7VH�����/�\!�*�.[�W1PȦQ�D���
V����x�/0Z��.=��_CT͢�D��H���W����>����'�;�ĥ�^���_��h�m}�>��8��\���{�Xܲx�%���������j�,⇎�}2�E��ǪUk��}�h�����_��		�|���V,9ܪ�=۷����H,�	��0e�DL�:E8D[�Mϴ::�ь&N�c����PQY-�^�:��A�0�i5L�Ks;���X�3����0M)�,`D��پ}���ѭ���J�SN躢a ��ɞ!:ى��AIX�D������?Y����~?�'���7e�%7�_��S�,�Xz!̝�Gy]=��A����5�p�Wa��C����pY\���W_���N��yv��M
��Ѐ�)C�1�>yʱr-�`���W^�����+�u�wleG�8��Ş?3�#&@2{��Ί	M BѦ>=
��G�<�_\�xv�l��w�;��f��}ָ����j�!"6�)��S���>zZ����O~���n��v���*|�m~����������������^�7Ϫ��˥�Jb��r�Y~�sE�å(N���誡j.�NQ�MRU�4-�_S�E��66���2�!�����.�}����n;�`�;8�@�%I8�$r�!�=~��~!y4�!���䴕Bi`�O�    IDATnBn��!�6�,��4j?��D
cU���i�L�"Ra����p�������!�s��.��c�q����ĺ��a깍�I0-�S.[�W]�^��ښJ�'<�xNa��=�P�@o�L晑a�S	�q�L[R�>�������&�=��؉��*r��L�HG�i9�j��`�ܹX��<DB"�Fwg��S�#g`���xs�V)PD)l=��\�/��9)���=��cf!�D00R�)tɗ�q�]��:+';܉�UH�#�*Ip2�pR4a��H,���{�g���m�S
�����y��n	ވ=�]��0���|_���A�tg/N��B�PR�8��"U�pE��6�[݂D����m�2�uc00�>E^����8�F^�Iң�hV<yg���� Ǧ}/��:43�J5�pi ��qx�n�j�L�>� �>�x�k*֮]��W�R��۷�'����n!��ܙ3����!�+Z��pR�@�4�<�[�����ڍD&#�ʵ���+7�"<����2�'����n��.��F:��/<�ꫣ�p�"L�<	�Ԉ��b*�u���Z��E��	��j��C>�BE$��alE*�[�de \1p\��'*&����;���$�7�|G�F?a}�>�Gh5�3�,��{�u��~����-�{�X-�c^� ~ON�����ψV��҅q��_�����_���C��2����_��O���>&k����Iⳟ��x�mx��mx��W���.����&��p��!'�<��N�I�|/�H��bd�K�}������_����?����#	Y���G$����c�*�a=N`�mf�#��")J�P<�e7��:V��U�v1ƶ�0) �
�r'������.��R�R�kd&2�RM��ض�3u�oۦ϶,1T�=�/-�E�#�ضB�'���i�b+�7䱫hrt��!��2.b��ؖ�33bZV�JB��4id�g�n�4��@e�g�ԣٶM�k�H~ar���ʪ�_�|՛ʨn�jӇ��_�5�����w�.�o���<�	y͍R.�tWl�k=�\�����{@�WE1�Ɯ�TAEA����Rѐ�U�KOvN�sy���s�aA�t�����9Ne�D�Ew������c��r�\�r!�\@O� �~n�젻���ft�W]�O^{%<�%?�Z��p"��RI�@�{K'���8�\*%�6~�I?sb3�5´g:T�4�u�t�t���K���q�&�sY?�&N��Y�P�(�����Ϫ"!1���ڛ�M�M.-����u��I�Ł�>�Io-�v%���N/Y2�iӄ�(�3[^��b�ϱYٚDf�e:4�eA�Q�g�I�PHA522��Q�_+�.���
��f�>����-Ho�@@��Lc�a��p�x::{Dڕ/�r��!��j��c;���"l_�0�'L��hM�=#��2e�r��zA������*����/5�:�#�������t��mfQ��������b�h�YЏ:T6T���K.��K�ja�]x��a�.ULe8I�۝�� _��w�%ާ�������C�HrX�e���/IA?r�$~�?���aY�pu�~��x�5h��F�߇-ol�O���2a<V]�\��b��B�+%��z�싄`���67cض0\b=��X[���_�z��DX�ɒ�o�
��@>�@�S@M�D������=�f�k$�V���"����X[��������w'/^�T.�?<�8�x�%1.r3���Ur��S��|�L�Њ���_a˖�dUG�C�&O��������ڀ{|>�G�z�MIA��۷c��;��?���Ml�'�6K��hA��6`�f�I��gY��Phnnƴi�俖�)�\ѕ'^Aϲ��;�0��Kh/�A6@l�)�$����&�ֶL䳭�KE��Ȱ���~(�OS��(M�(�es�c�4�CjӤ6��DI��
�wHŶmL)����߻�����S?�ǚ�8#���@g�����ɼ�j�_K��S��2��`�]N��|����y��
�R�d����,^��<�����	�.��{c=��?���s�1�e�;��ѥ�^Oj���ƈH�/u��,�L^��Rr0wKZ�n��Ձjɸf9�@�(�6���i˟�	I��7���5+�r�D�&���s�8���7�\n|��u������ؒY-w7Me��l-s��{:ň$�A.3���A1fa!��:'@��9���J{uU�͞��l	}�:b)�k�FW<���C��	&OC��f'����,栔2���{����[b��ж����'�{w�!�w
���o"��$�HU�ʀ�5'�Ҕ�kѰ	��KN�^锲Q�L#��_�|I|��^,
�<���O"���J�E�\E4�<SBu�#�{�ӹ�����G��P��O���޽����+f5��uV+��0�b�;u.����pQ��	��"����T*�\��b�M�O���4E"\��%Aq�H1�t8��iP�����it�6� ��>���q����d�+�x���q`���I���˱|�Eb����x���Pb��W��N��E}�
���#A9��@�_������<~t�FGo��^�_��b�k�^����M�|^����Z\�x֯Z!.ov�����P[Ō)�
���1��E4��5oh�[����j$m�bI�|��0�T��0�B�h%��)8�a��N7@�����uؼy3�;&�S6)�zǯ�+y�jq�k��y\�����ez}��������� � Ò�GC$3�L����^���?ñcGPQE�Δ����_s�~�e����;�����!��>���o݁�{>���AG�I�Y4��bxx�O�;� ����A"�W<y���ɓ'K��i�D��L���9�g&8�3���q ���Uz�]/�4��~�Z&�9_��I��W��Sty��*�������0�r��� ɯ���k%ʁ���p!�Y,[A��#_q�F� ����/8���K���A����Jb���ճ�_9#�Љ���ICt���ߋJC7�+�Juuu�\ż�W��<����ق~����l;�@���cw�ˠ�ف�@?|�0���h��E�զ��Q7�IH��Q}�iA*^�Mc;0稳�]�7gA��V���;P*R�ŉ_rVS}%�Y�
���0�������ǻ��a,��!�q���q�� ��G������g3)t��Ʉ�4�B6���^�ӽy=�y��h�7���f:�H��_(iq����'���m��P��&4M�*:^��y8eFP�,�V�p��~���k�VѲ8o�$��w�XC_��#��N���-jU����9���g�p\\�6Âfڰ����D�����C������̍�m�l�����D\%4��W_�ƚ��GN�af��$�51�I��� v�ڃ��~��fښJ�l&�y�4LĲ+nD�Ĺ8�9����K[�Z.��Ǝm��l86�\&+�0.��rj�m��]|�P���CL%�CD���U|h�㷳�1�b'B
׬_���*��p��iNX\,X�u����ְc�{x{��%�	��$I���eŴ��E���ũxpH�N��Q5&N��@8��'��
P?�	�]q���s�^���5$�<�w���~U�d��XD����"dFޗ�>�qY}��p~����?X>J\eq�XU�A�%_@�{s�F�,JV�%e�cqW�f٭���;Sg1��&�t�(�5�Opt�4\�Tj��l����IKA�?�@�O=�'<��ϲC��=3�m$�ru��2_�鋈����bϞ]�Q 2�󥦱���w1q�d<��+����II�v�W��;������{ݧ;�~����ޮn9Kx���;zt�鐯���,���;�<)�3gΔ�{�|��Q`���Bow�!A��PJ7��z�Xѩ�?'SK��T��+��G�S(�3�~�?a��rBʫ��d8#d,K9�/�>Z|�Ў�5}��?Z�G��I+�ܣ͆c�����kykW�˿1:(�^�N�-�l�Cuu�?�xݕ�Uf#�u�������e��{�>�ے�b>��e8E[lT�*)B$�xH��	ML��<IX�	)��N�'���t����9����#��9]BFʓ4w�d�MѠ�Ua\�z9�/����:Ԏ?��8�vR��׏��W_��]y)BAgGFs�<}H���4�4:N�@6Im�c�2�G����.�h�Bݑdҙ��i�!6��-E"�c�qtg�ľ�$t��z�:�|��Qt�Ǡ�xTQ/��h����l}�m��$G(|�9Sp�w� ��}��z�����1�Qa��3m�΂a����?gK��Z�"n���
�L�l+�-�3#��	Z���+3��8����ڐ[lO[��KCP�P/{�hE�L����;O���6�ܹSX��&	��u�.M�}g-X���~#�����Ɓ�8oE�QUS/����^Y�p-�Y�nɣv��z��L�
dKh�������#Ì�C Y�K�(�N b���W��	��{�ǎɮ�&$uuu�2q�|�C��"���//�$I&���H��\�h�S)�$��th��qط�����'Oy޾#���1Y�� �45���OV�K�%:w���
p��sq�%k0n\�H���aly�M�8tL����$5OC^/I����Hg
N���<74�s9�d����Ti���:1�l�~��M�󹌳kW��o�C!��6�KS��L.���OfD���%ɭ2��_��'�����_�Sz�#I!�It�i9�����i,���J,:�<��8�ή���ux|!�����`!�~}�����vQ�p־l�J���;����x핗p��$|>����8Nwtȵ%��Q�rC��1��4��
L�0��������ڊ3f|�r%{ʴ�Q�4�N���cIJ��*�v����%��Rn�X�e�X��G�/���T;z\tBv
7���\���]��_~�	Y���:S����#$��G�=:@�)���Y�N����韟/񛐞�Ӹ�B�3��� �]>O���^2�|�T��Pw��������}%���Գ��ޯ:�W<����!W�)ǂ�NC�逕!$Z�����^v��,��.�P�V�RQ�Y�'�>����s� ,2�� J4C���F�����Jٖ�=$Z��g�J�eTq(#쩙y�T��~�ܸv)B*��c�=���vҳ8�1V����S�_�H�C�c�LH�]7?؄�(���f�e
����Y�HX�ϓL�8p#!}uu�h�4CYG{�+��u���1��pE�0n�t���b0�mK�_)��:�J����
��HQFR��]<�q�W�99=���~��y��Л�`�*�9�t�`+�kf/L(�$'��5�OZ�r�Z%��RPHg��@Ԅ�/������.j)�b�ji����֩@˘��6�e�T4�oE��(�ߌ3-$#سk�n�*P��+����`��w����Ϣf�d�|��w����w�3i"o�����3�в�	j�}nI���5cZ�-����a����0�MN`�g�N]GP����FNKA_�|�L�ԡ�vw;:e۔C"a���l��Ģ2���I���ǝ��
#�ȑ#覿Ak+��J��x����	��2c�Ȭں���3��:|��]`A��k�;/�"��>V��W_u)&Mh�5L<6�����{D�x���.�F��V�IeE�悃p�u�t��m���ɓ�y~k���\������e�p�왨G5N�^�p$�>G#���R�Xhy�3D��s]��C7���
47�
��?0������_�P&�咩���/���~�8nn��z���WA��l^X���0�~����fY���B��`ι��7��#������KP�h8$Ll�O�A8N����Y�)aljj�ezMpBw\$Gu�IP��������r�w�c'1�A��@:�"æ�d������|�T�g�c;��9i�-����6˰��`�|�U9ٗضe��Ə��ùmw�s�˜�)��=��RT�qp~/��9�sMO�;�B�#���zsU"��i�\�[��h��UQEQ��)٪�����f�4���j����+�V�-3k�vFQ�MՎ�m�p�������|�-�gp�~q����v��w�S �lݓǡK(
cŇPU�Lؔڠ�E��O&��Zq��5 )x�����6 g�7�.�p���WDd�*�A'x�9�[�z��;d~�H���lTE��?sn��j���<^ߴϼ�'���4PK����?���ť���;�����P1w�m'0<�+���� ���T�C��¸+���0�B}�X�4�` U@oZGwJ��ǻp�t)�OU�Սp��r@�UE�H6�6w1���w��wߓI���QV+���/��E�����_��&.X���$�}
y�N���E�߅�l*��<�)���D����	�C�z)/��!��
P�d���UL �6�,)���B�:�\L�>���K#���yOW����ߏt2��,CLJ8AVTFp�����/���0Tp�+m�=����'t���G!�ICO��.8]�௭C�䩈�������5�9l�ZEy���R
z�� ��)��8�X��CR��G�m�ӑ�)�e	i�
�{��j0	I+��)S��h���yc���oű�m8z���ol~L�]��p���gr�@�5�S$(�u���8��=��o�?n/Z��.��i�����q�A��ݜ��=7s�����*�O�%r6N�=�xj��x��WQ���㕢�1��vI�77~+W��_F]�r.6���X�]������b#��ĐH!��G$�j���B��'�ņ�oIY�^�mG��&D"dA����ԉP[�Ͻ+T)��O���;�G�RP$�4_���K.ĝ�~￻o��g��{ER�P6~�=]r���2�:i�PCP���'s��X��ܱ��������k�D��]�܇�6�Y���fJc��s�r����r��n��"��
9��rY.��$�A�R�TW*r�����۔��\!�eJy����|���jyhZ
�]d�����2�7�j�*���+䙒�N������JAQ�Ǚ���(�F7H��C1UM�U��䲔\｢�����ۥ�*
�=�bۺ�cX��[~����uK��V�T��P�2�8k֬rf������-�gpv��Gv��݈;�@���'�*0�a0��,��4jT�bk���uk/����-{�����3�^I����? ]7���"yE�C��ss�r���b�`�yЋ����'�ǹc#(�ǎ�����|p��c���x!��Q__-ӫ8?QϬnB�B��GۑC�F��X_7�ٔ@N� =:�-898�I��@�Â>�1$A�'�c��n�>Ս|�Fk_�@��b!Z� �Q�blU�n݌�^~Mt*�ˋP8,��Wʤ��]��7���Ϡ}DR�byQ,�ݎ��S�mF���f�#EB�:�\z:	�S����'�g� Wt��k�8R}'�Wr���{ %R���kK����2a<f�:G?Nq���:,���!�ZFjX�\>/�.�H��)}"�+����A�θ�_
`Ў�m ��N�\��H�%5.�_��ʆzē#�'G`�e�h�!	�9��D�e";�����L�#�ep��s��������^;$LJ-�)��o��Ж�S�oI��%LKW�Q�;�����'�v�4B�j��w0����7svȴ��p{c9��b�_ ���
�����
��W�^���cdB$��?+��}!c���ZT��y��2��><��l�����eOd�(���=��u�bŊB���'z��bk,d8�_��T��|��O:cI���Rl�II��9LWw/y�9�?��D�M%�"+4%;�����V�Z�L^;_��?4Ml��4m'NuwC�VIF9:'��˖�k_�	[�|�����z0��ɑ8N�>-
�����|n��%�ٶ�l����D��Yܥ�){+0S����a    IDAT�H"��Ј4-�n.�ߖ�<ׇ<lF{��H�/��P p*Rzy��	�7+^oN��E��4m�+j��E#@��U)s��*2"�TL��ִ����y�4m�[�<���(F��t��-��T��Ƣ��a4ɯŢ���G�P�ߟ�N�X�ܱ�,?��H�Π���Գ�.��<~���v��C��g:z��V&/D_(4,�M*��$�`����aͅs$��{��c �AF���qbH�K��N����+�S���#wU.qEz54FC����Xw�T�����G����&�n�mc��X�|9���厐����TzD`NZ�=�����)�<�8����a%IU�*i�B�����2Z�	Sg"gi�Π'UľS��}��;�H�`�5� �U!q?��S��/��'�{�Ǐ��`�E���$���1���'^�[;��O�7��@�ˠ/�!a/�lUi�Zd�#󉇻��^��k��
y�tI�3K���J�����p�aԄ�Pj̽<'x�:\.9���\~�40���F�����>'T�MPG�v����O��Z��M%Q�5t��}'q*n¨h�Q9'b9�7r%rԝ�B���Kw3Mȗ��JJ��/:��B���W5%�FA
0�b�b�� w�š6�G-\��\!em��z�;���9(S�8)�L�����0PV����.\�X��h1:
�����ʦ7�Xd����2�\ԏ�G�|�$
|?�)�4Sb1��dq!�b*AP�(i`��ɺ�6}�H�$�@�a*$Q�`�!*��ȑ�F��m	<��׋ �����T�N��?3�M��l�ĜHU���LG�����2	�	U2�K���)lޢ!�⃂�1�����8t�E���C����T>j����;�~�*|�kQ�{`2���_h����ko�ݻp��&w�<�Y�\����-�˖����Y���#�=����C&t�%d��v�3,�|M,ޔ����?��F��"ɤ�{���E��+K�z�$I���^6IT�D@�S|3�n�UG�O�<�7�.�p�+V��|���W�lA?�[�_Ot^����aA/X
�t��J	:�A�ξ �-y!���<",��<�_p.]v��o۶�<�$���L�[�т.$�t��&�#�|�a������^�J4&�Y:|��J��gN�g��c#��bρ����I�U>EÒ��n��rp�����]3̀����[N�8&�*�}��v	l'{3U�hNQb���%�� Y�6�� f�slo�=��J�xW?�;������31��E�Ei�:gR#�n9���&l�����W�*ڨmj��|�sX�t�h���8�_?�Nf\���Z$�
�a��#_ɨ�4�i�D]��r�:�E6;��E�8���*d�R��5#2Rй;��@m���g����#o�{���Bɏ'y�h���	��A�9�	���n��.\,�(�U�9r�nG79o��f�#]()	����ʝ$m`�?n�vv޴e�I�R��g���B 
,[G��ÕbA?�1U
�?[|^|�1"!�]Xܜ69�S�Q̋+Y��I��N�;��kW�СC2�������uؼe+,ՅYs�c��h�8�>� �R,|l��.a��g�`Q��F�z�@�:F�q��I� )����;%}>Ņh(,���a����>d��m�y��ׇ������Le��29��-�Ow�	�Mu�������G�@�N1���D]4*M��|��4Z]����(���>��������Di�b$�4\o���9�;{&�ϙ��Q̑���'O��ٳgKQu��x�/�!�L����e�l����;��{o�M�H`o���j�@��Wd�1�g�Rٲ��2_��ѦZ�m�C%�3j���g�fc��;��0��CE�W�R�rCJ��.ٽ`�컫p���X����>����+p�������]�<�K
zMބh?�]=0Sԡ+�ݨ���2��[Pt!`�`�0�i,�O�)�ȶ�v��c�d�BH�L�d�x�~��`���1�ӱ1��@�K�D^㶋�[%�D���5�cɜI�@:[�#�<�7_{�]s�2��x�C�	�0*�k �C1�uj���I!�����G�Z�W��������*��%��hh�4�@CL�J��O����B}�84�kFMu5�!f����QSS%����a<���xi�fX� .X�\��ڪ
��}��x�խH����ϣ;��w0C�m��S塨r�dc:���:�W�D��<)��3��(iT��h�j���0��ѓ@nF>�1іҦ��;���:'�aU�B�����Xt����x������ȉS�u�$��&��X`�Ltf��ϻ`{+$ ����t6#�~ʥ� {���1��#����ȋG�>gȄf���z`$N�*PĲ�*�3�<��ǎ|��.�R*zp���"�3i�ļ{j�iV�*8����u��}�I;�aԗg��Id�cs.�c۶m۶m۶m�8�m;9�s�ɉ�}ޭ�O�#��ꪞ����X�O�t�ѯ�^��������p��f)H�N����&�� |��U/4��sF�^�
š�9��.w�y�_��������cs����]?d�1ȉET��R�f��~"/��[��Qױ���h�_ܖ��!m�i_-ZA'�9<��+���;-�&/��Z��~�y%5�f5Q��^g���_L(�]��ve)�aU���ȅ��j0
��p66�N���&s���	�{ǔL���M�V�_��@�+�@B<#_�J�G�;;K1��3/^4��-��≫J��jec�b���`��� ���B'�yk {o�V0����0d��HSؖ���0�c����~�\�~��7����/��� ���?����Q��ðzK)������V$u9�����J�pV%T���X�j�r�d�1V�sF��&3�{���;�9�L,{U��H���ܺGU�I�����J�r���!3l���-���9�`;�q���@���[��ȱ3*Sq9��`)_�d�1��L��M�8����X�2G*�$�x��5�єZ���Z։u���#@Xw;�r���3�^����x�#�����̉��v��w5t�����a��۵�u�~H��}�vù��ڟ���l�E���x���*P�M�V:I�@YNex�[�d�V�2��0},a����$�
?��)3�I8����T&i�c�I�
k�Q��i*xM�4�Z4MJϽ�����O�l;����z���,����� �n�;�b�#1�8D88�����8e����U�e�Im����~ $4nөh{*8�~��n�|>p���Φ�wO+�G?},�Xg�p<I�(MY-���Dҡj
N��1�=��)�����lX�ÕƵX��<1��LQ!�2{~�3ba���ݠ���.�\��.3sZ��Sl��eE�8�mm�+�}�g�w�|�O�Qo�*��?G��_ð���?(3��#��g����1eD����+�����b7e	�,Y���]�Ӛ�'�_��K++�!7a�H� [�>�~���dy���
zsmjM��o~��x����o�<.g�]��;�Ҫ�H3剖� �m�^�ԫ��Jn:�ĉ�7l��*Á���n��	J�wj��	�WE�O�ֶ�X)a����L���[q@�xϻ�
���)1fY\ib	�	����0OU����ɸ��f����\^/b��aP������cبg�G�Ƿ�H!Ġ�%�ϒ�ǁ�������O��>�.%=~�wЫf\3����5 �C�٘z��k{�f0ۉ���[͟tx�q*�%�Ls���Ł~?�"�KJ1�E�M��H�{��]�����.�կ]w��j������v^6�b��'5:�.7��v8^n�(�M�R:Ǘ����E��PF�G#(����eT�*ˊ\��H�GlR�'��4�a�7��|cf��( �0�[E����#���z���:� ��v�<$�mH��G����+
y5R�l��_��6ݑD+0u lt��眽VW�$��i��kWxL$��11�)û6�s�!�"y����ˤ�X��Z��lj�V	&6�`��`�u@�1��p�=����Rd)���� RY��A֦�u��ơ$�n'��'�C�g�
�~:��C/�M�����VωE�4Q��p��Q�U.��H���0jձ5w##%�M.g��΍�#]��ndy�N%�RDԚ\_wT��btT(�C�q%���G��4i�{E\'�� 1�����UMCz����!��|���2^��ZNxos�p֩Xج���5�I��yT����҉�X1&�/���ꅢ�z`G�͸G��}��z�����q�X�+��Yv����q<���o�&�v����a��l�5
� ��kY��zX��~����:�׵Fh�l�,�W�4yA�Tn����y����U��f6��ф���ӫt*}��}�mwl���?�c�̞�o�ʨQ3�췩ѯ5��b�-��I�7�3���B~O�5� ���W�/I8D�<|�:?Yp�pZ%dhb�R!��)v(��ΏKۓ�w�i" �s�Г0׼/��,?R�0�� �B��SS��O��ϧ��*�;��ς�����0Cˮd�B�r�dU�,e؀Jĩ��T�A�(�R�-bQ�7� ��.�+m윸x��!��C��m��6ހe�s��f�3��j�k����ݦ�#�����8K��F4XkI�M!&{0��|VL:&���hh����$1�;:zH^��˹����P#i8
>o���l()vr˱�n��4�s��k��;i�.@TYMά&,=Ґ]�X�*�y^����$BCz}�Ox=\�D�f�.��:��F�c-�]Q��B|��'TPm'�1�����k��g���/י�
]�S���?R�r���\��!7~|P�睲
���&�\����l������eeĕ���8Tѱ?�4?�$8KF���2�B3Yq�z�����=��B)iÜA��,1[��X�Rx��������/}k?B]<p�tUT'������h_ �d"�ąe�
�}�0��V�(%u��K�e��'W����8e�Q	#.��jI��(JY+�i�E(ц��>����������)T;r	��0��d%��͵SH�B�A(/�H�t����W�E�2L!I�ݥ`>�e�9�D0=���5�t�i�U*Z_��1��b.Ȇg�,S�PԚ�*���cP`�r�H���o.1|��気�K���@�:]������� �H�v�_���n�5>�鴜
|���7�X�nzn��M� 
�+���qMÑ�>��:2�=�Lf�����>���h�ۂ��@+�7O=z�~ ��������4q���v��"�:-%T�c�g����Oa@T�FPc�tLi4�5�Ba��ދz��Ì�E8&yK�+�;#�|�{�E���(���/X$"~��^�{��}��;������Z�\ �����z��rL	�V���˘(TI\8��F���voX�.:���Hp���^lU�GK�pN��B>"� ~���/T�◼�=�h��&����ȩ���O1�����V���17��q�]��`ψ��A��߼�����qbK605!?��-�'���/���`�;_k|�6=)T�Uݚ��;چd,�h?$�R�W��$Ґ��Č�N5��|믫<	7";<����h��t:�2n��aZՀa>@���P�p�m����~�뗙�A�@G�j�|��2���ru���_s����&���1�����ɩ+c�D�E�KH�'���Xo�W�(3q��B6]�u0����ꕅ�%��=�O��^����.="\	I@Dg� @B��DE�v	�<��܀�%��Agov%�S8Z����l/veB�Ij�SK�M�$� [�Tc�}���c䊶m���\A���޺C
8c�G1G١:i��>���捿J��2�@5�ۇ#
ύ�9�2�##*-z\os��ȖY�ч�5�#o�굘g76��g�i�A�I���Ŋd��G����Ӂ��Vćh�����bI���Z!;6s2B�P#��;4�x<>�JF��������l��Ǜ��yLiՔq,;`�,/J�ۊ���a�� �g���܃`\����h�&�|�n����$�B��m\��#������s��S&�8`9g:�A�`:��=y	���A�c��y����?���d�O+
���}�?����0Z� �	�@��v��qNe��1 ��p����yW�Ht��
�t�!��ώ�D��ѱ�"��fn����H<�����KU4z�{D��w��j�I��Q���_�����
'�~�<�$-��<3a��P�bԡca�`��fx���\��b>}G��x�w���O3�L���������[7��s�3�0/�Z��фj(ó8��4���4�rzU��B˘-����n��_q������:��n�w+�x~�m��D&!�,��4�l$a��
�Ғ<�����♏�"ƅ"�W�!"&+�|=}1Ph���,������g*L��5���M�����=�,p�:1�iU����"U�Gєt���*?����y�s��=��ѝ�0�Y&��lt(�B�0� k%����H)'��3����(���\��9���أ��`{�+����eȋ�ڹf[��D~A�e2)Κ� #��������h� �t� #���^*f��B�*=_�4�t�R6�Ϛ=@���d�뭣4}��_���V`&��;&����^�:�׈`�I����[
���*�$����a����NJ�Y�d�g#~��A(�	���{�A?�k�8u-������Z����~c̹1|է+_
H�P2㊷ǲQ��'#�Q�'kw��,|×��4�@��0��x��(�#��A�3����A��̩�~�vz�7���*y,���H�i��ĹX��'f��.=܀�vD.��#�zA�0d��Ey��J��&M�-��"-��ѵ�m��717��ߩɈs�Z3�0䓞����7tƓ�d���Fͷ{���$��$h����}ǛM@����K��x(y={&�FP���C'1]������.t�nt���kɧfR��@|6��Jyvc/�4�<����~�AΟ��\W��o��U�Ƴ��ov�p=�)'�I��ߚ����Ȏ�Sά:���*��J��D�8�wN��Ԋ�������)�^\�J�6\�8�"�

���Nsj����� �ld(&��ǌ7����c�oXߋw�k�"�x��c�^�k�=;n�
��f������}taLO�E�[�D�zݎ��L���5j�8w���s*�;M����iR�ë�7K����xJ���1�7���~��$fˮ�%�����]�d��al!���� OM�&*�)I��<�h�{h ȑa���t��>"暺�o�$ѕ��Y������*�U�T�7�h�A���~�Uz_~�0�0�h21�h\t����*�1�[���,����!�=�۶���<���ib���C��z�8l��$n5كC��/n�B1�Z�YB �W����*�۳�������A��P4��Y�����0������4,d���Q;lZ�J|�C�"��l�8,��F���N 3����8��h����L[i	�0��ǔ]����`N̩�/�����TkE3�㜱��f���S���l�I���N��� �$�aL�x�U����b|Br��M;tT���_9�L�?�jm3xo�+�M�k������s�,�S'�\.-�z����65�����XJ�d9����z��x�ꐔS���{�XXx%]�\!Sv���P�k�
}@#�-.H,�q��	+S�If\8�-����gE��"���v�6Q��z�$[V0>Z;�G�T[%A�L��Z�^�9�:HPbeISf�/ӱ^/����딚ғ�R(h�3:8���N_}����䁗T=�n�ծO���J1#���C��,x��cq�>[z�NKݒ�h��LAX���s��`�E
�+R��G�\�����ˣ�,�'^��i1�FJ����E����̹��]G#��s���|\p���n��;�_�[wk1)�k�9�!�KLy�[h���#�z:�|
�t�5.���ߴ?F
'l~O��4����O����Ov2A��W��2
^<ܤ������[�;����9���-���=�(���Y��J�֭�����4z��A'7^�L���|���Q�+����F
�2%m}=Q��'��k��G��ܯ�գB:��z�k��k��q�e���cn��v}�*��m�L �e�c����xk���?�)����n���%$)ʕʢs��b�/E��A��R��@�7��!z� ����`L໣9t��<�l���r��9	�1�ΠӈX��jÙ�	�f��`���35|���|�*���LJ�.�xc���� f�����WQ���v/I��~�GFo�gŎ��^���ùj���p���u�7�.��L4�Ț~�"�!,�0���V$FDכVl��_��@>.�7��e�ꝇT�TV�T��9� ��O#yI9t��}#�L�8�Ȭ�ѾF���;0��\Tfh�l|B	OS�؞m�:t虴АR��i�֝XWI����̊�ӊx���WxGGB�v�\:mZ���C��Y炕%#��sA&���0�7,�Ue�汮�}���Ц�?�X6K��#�]���z$p p�l �X�����B���r��Kq#��dî�r+ȸ��D�O���H��W&�~�J��M�%�$�m�Z��'���x�m�]Uqsr��&��ms��W�XL�U�{��&)�d����c��=������V��%ೢ��K�/d��ۀe>�;o_���������'�`��0SIGE'p�&[YNW)ή��Ľ�ɚ�^i>r�T�6Q���/"|�q���B</�{��Ե�١c>8��]R�Xo>,�z�*�s�8🺻�3w���@���v�����N��k�'xqk��r$l�ߏ7〔�)�=;�7������u e�j����W�.���� 3�������;K���$��#A��@O�F�]��V�:h�v:ǔ��]p(s���]i���!�F�*3�c��x�.��N���8�{nR��ݓ����J���S��*l�������E<����5�ʜ�m���{i)�������ϐovE@���o��	�Qr9Bn�\`# $˲(��X�EU>�w�ʦ����t�\p���W�ܾ8�����w)��7�Cgg[�h��"$%���˂���\�� Ο�}vG�7[�9_�y�.�C��q��>��� �)�2� �\H�)l��C!�U�q�6�m_�>���������.�^ه������d7��2DB*u��:{�4G��^Ӵ]L��&8|�����D��$���� z_0:P,D�9g��d%���UlCL��}!�O��bq���&�I+ �g �U��Sj��aE%�<�X�"_��L���9j�a����t0o����}ͷq���~!	�]��PF%�;��Ԡv���#�'�ҥJ7D���`��g�!� ���Z�jD�c�`rU�*��e�F=���F=Rq��ɧڜ?�TQ�P�3"�m�p�)�x|�|@�3��8���f*�7�t�%�4N�~��ժ�bQ��NB7I�WT��*J�?ш��BZ���������quzr~DF&f�M�����#r��<��z�r��`F�)�+� g��]��y\3�u��GE?/�����o}+=�������G�������Wo+�Y��᎙=�ykh�w���8��R)G ���`G5qd�8������/�Z��92`M{y��&��.��0���jRDS�-Ρ<�b<+N�{ӊf�9�J�ؐ��~��Dq���\e���}0���� ���M���7��S�x����V�|�GK�����I���d#:F�Lf�`����;e��b��RI����s��@����r��cz��<�']�۲tV���c��`@Zg����Ek���8'θ��a��o˂@�R�f>�(q���3e�G^����3�F�/���.�}[ZȽ��P�筁������No�;���B4�j�B����'�0`�W'΄�x�<���$'�4N��8����nx�"��+�h�Ө����z����A��=�,��졺���qY�R�
wVZ��T<σީ;�H7G��������OW�j������f�Z�A��@P���B���e�{��5މ�'MT��[Smb�K���gт��������_A��Ͽ���;9�\�P9�0�d^�R��FH�*��	PU$,���mEg&��q&���������*���D��GtPȄ�d	tt��/�m�͎�r}:y}�~dh��l��)3��?*Ӧ��: c�Y��R-�@R㰪Wv���'�G�j�.�O�̦�V�Ff�0vM�2܍� ��^�R-�c�u~��K�{1�6�hf���~�9D!�)� �p��Sh���5rk[�����ww/'����_ͲOqD01�1�8v�[+�"[��,�"ћ��B��)�P�i�^�@D�5c,0�p%���՛�˾I����$5L�Cʏ(�	�Q��ў���Rr�H��^(����'�p��1y�EHP�ǋ�^����7��+�e���F���o^Jr�BL)���l�63$\��\�e5��V����|A�-�N�]�PhvF.>(--�^������n4����<��$ƛ�TrxBv�\�bxMn�7�c�&t#�1�?��[S�
<���_��=H��j���Gbqoe3�@���p���#),V(EU��2��v["(�&Ξ��~1�n��Px�S�?~��D����
��de�:���`��"�N�*~RWP�_E����䶤Ϸ���F�1��!�M�A�������^;�K�AR�e]���)r-!r�ߣ�5��4d��=���B~� ��"(����C<(%�h�e)*WK�����Φ�fx���<=�jV2�Mp[��0: 7�_(W�@�={�51у)Ӣ�Ӌ��ŕvݴ#`�������ט��p�rUvS�4�~a���C�
�'��C )d��F�?�;�9��ﺽ2���j�0�����g�� (6M%79�	L�3#���Jl�C;�b�&>���M���3�7ſ���o�|O�B�����x\n�;���.����(��%Y���u����.g�}F7�����%nֲgI!����q�������|��	4.a�V.Ŗ�� Xbeɍ��J�s�t E�YԞ�;�F�;$��F�R$���k0���f��+@v5�[gA�U��7�:AA=��a0'/lBA���2�$�jz�:��O�a3 ^��b>X%�37��~�!!&GS�:w���n���$3��$�J$/&1z��13���e��;�@�k�N�$4#G�-��W�e�DOm��t���������z.� ����ꠁw�	��o-�ajM�	|Q�f9a��j���Kb��A\��Ԩ�&�ť�a���R�P����K�tOA�}פ�w��6:�><(D��w?�L����E�-1�d��g�;�R�sJ�i5.�)6߆�p-epF��yL��Cś�$*2>=Qt������a�iQ�j6��T@���9�]I���a���Ȼ����v��}N���a�r�v�o�k���ʹ�I�8w�x���N��x[�tڹL��8Xh��\d�7*�K7��s���a��a�����=VH�,o��{G[�K���:�9�M`�����������D���0�d-5��ʖg�%�v���`M����%t�J:
����j�:~��c��%xp{7��ɻqh�9Y��<>ng�h5�ɠ�R�7=I��n+27�{��?60>��h��B<_wp9���#����7Ŧ�:`	�Gp�ͤ���"3"Fj3��=���\�g�{���oRΜ� �lj5!���k�]M�NF�uN���2Ѐ ۻ�/�Khjг���7vє��t��W4��������r~���V�	��e���ǔc�0��W���� �l�0=�pѕ+��N�.��ϜB����³��/�?�V�?~��F����'�^��/Ώ4���e\�m���/��C��YEҹr����8��I�"Y���d���i�^�H�E�5� .��,V��rx�D�Aw�6��J��\����򼞖:��T�LX�V�0]U�	�o0�-m�<�]С.��4������A���~_�s�y�I+8�5�͏�����ؠ�&s3�"d0%E����\%j\)�9#W�҉kb��-R9��?`^��rm��m����ԅ�ҍ&O����5��t�,t̀�o��X�R���j�N"x(��
s�'S�4$E�b������m�K���ђEj�q��A2��������e�FA�}.�<�i	��c�����_ұ�p9c��C�T�>K5����Ŵ�Y�d5��)$�8/��> ��*��Ū��Ǡ���k":�ߦ{ZR@QL����$��.���L�$��"�&1�w^�1}HF��޷+O�!�W��K��a�<�A��^����*���(:���.��v2�y9Z��J��>Y={[;Q��Z�/���Ʃn�� ,Ua���_Ju���b��j�<������_&��&e�Yo�5�{�⾮�������O�@"d�[�� �O��O��Q��z�U�TO�v*$��eם��nb*���8��G�|v�{���ly&��@��3r�bQ4���U��D��iu{3�ث=/�Ǯ���e��%�Ą��ڙ1RܻcG3���dD�-T*��rPC�Dv�� bi((����R ��m��T۔YK3@,�a �ڝ��� 򶻁�P�3����4Qx�כ}�� ���;�.Z5Ϣ�
k�垼�ቦΰ��V������ﾠ����q������P�F���`�=]��3�{�鴆��f$(�9�8�V{29KV:�ɇ��ѣ����dp���qI1<ű�zi� ���
����Sz���R�5���������T<k��)�dK���=-���=�.�9�~�;k/XA/��8��R��bs�.��L����Dh� ���dnf�����7�`j'�O����4\�I�N��������!��-;<"����y͝v��(gY������a�6d$d��"i����2LI%g���2e^��بK�J;Txd�h]?a��}?�Fr�-��s�̔+_���J��L<��|	푱qlpy>3$��;d�Dj)i3������{�^3���$�M���Id�݅J�E*���Cs�qC_$BQ�T�Ǉ�&�����Ψ�d��H\1�J�̓h	o�\K�[.��aԍ�{șfp]C"��ޯ���M�i�`0K[�3\_�HG$MS�n����ym�
\n�sA�XU����qa��,����;�NY���<kg���c�w�!,�L�!�t�bj��ձ���y=��������,�0����f���~7B�+����Y�K�D��6��EH�/1O�1�H�6e����nN9R�C�0��0ٿ���:`o:��|��3�N'�&4��D���ì�Q��uF�,I�4�v
����Z/����.�����n���2��6A':_����	�oQ��6��Ua#H����@��s�"�{������e�*��md�Y�V����ӌ��!T!!�����2�������=�3W�%�-;�m.;V�!����l���-�QQ*��]��hS�%�"Ѡ��R�ƣ�&���#��p�ਗ਼��̒+�YE;�TD[r�o����z���Ov~gD	�����*昳���7�ʮG*;'P���$ ?w�5g��B�A� LġS%�d�qK��9�=f��K���鼽(��AF�^t>���и��3����D^���kc/
IE,k?�-�+��Q	�!x[[ÿ�xM�� �F1�y|�h>�jK�en�u;pA@v>+{szM���߲Qc�B*�$�cR��"k(��U*��ƒ�6
a$�i���3n3c�S7���S�?�uf�m��2C�����N����0ȡk�h3k�1n�#���L���βg@U�:�2@ƴ�H�j�.N���T���r�\R���gm���k�B�)�J���3!�l�V����lJ����zu>�$����4��Ǖ0���%�L�S/� ��8"Ԗ�lC���tUʐИ<�x0�f�p�M���%=0m҃�'m$a09W!n����պ_l��+�s1�^Y@���/����z��]�򠠍,=���Z�����!n�-ǩ0P�+�]Bjo4;	�sD"���B�+��7e�>�:�����@�R�B^�����mDz~��[�W�?�ֵ�\��	������+x HJ���OK�2���5�җ*��c{�'۴�Z)�)���I?Ջ]�f��=�K	�,�xL�	.gZ�O��`�%y������,v�%�Q��"����=��֭���d��N�@�����?��Z8B�A��y��p�u�yr[ηV���h���U�/��U�s�F���]+�w��Bg��S|�lR�I}� ���j`������}8?�>��5_.��=�P|�
���ǭ^{2���H3��i�i�<V��`��3�o�+p��K��ѭ;|�����#�։��`8�F+�a�)���"S������m�	Osf;!�Eͽ���y:Pl����gY���#�N��a"�B���T7�e���Y�����d��j��<U�;3x�a�:*.:�����$Xd3y:�� 赗��v0/C��<�����{���'1 D�iƸ�Y^���m���J�3�kN��b9& �6���L������!_����x��w쵑������ ���C��Y�'�d0EJ�~8�#�ab3�;@xm�C��eKf4�2��Y��Ȱ�������ơ�(e�s"�xh���z;���_N�r�r�l�����A|��ܚb1B"]Dw�&J�U�R������d,g/Sd���ݤ�
)���M�BƟn�@[[mr�����#�P;5���H)�{�I	�h�1D�J��w�� ��\����i���-ܳ+GYG3k��_�XٳFF��^�@�;�!��(]����ױ�c�&�����M�C�x�7�=s��~����pI�/�1�>Eiz�/��.�dDC�|��H�|��s��],wm�{|�������5b��TՖ#�fҥ<�8Ӛ@���4A'�@�;�Q��:�BKt�7ku�
������m��:_�f p"wiy�a޹�Q�߱~
2���d{q��}:�sܩ�@�������GK,�qᖺ�R��+���&nQL��;�Bs���(2
A)�@n��́`MuZB-��S=B�X�W:y��~�����̒Xx���w]��-GT���'��"�LEL�I^nOކ�FE�b"����{�1��[�
D'�R��Y!�_�&��]O�9z�o���>�K��Z��
���Qm��PM���س��D D��)�$�X����[�JTk3�gA�?z|_�V�j?��k@U7�߫�^5c��2*ػ�]Ԟ���i2e#Nk,��jj �9�����X�J�ԾT�xi1�6[�LG �"C���7��8�::��?���W��wۚ��=&ڗ��B�l!��o�q
��c7�AK�TEX!�uz�I�k9��sKM����b 3�V\ѬIP5����&=q	,O�}4�~���پ�L��0���I�eq��!���
x\9Xy���)Vf�;̼��[�\ѵ�o=��|O9/g]P�l:�+���-�]��r�B�^�[>f�^\!`��	Nl49�#,L��G��XWL$Kb<����E�H ��_�t1��䄠?����ȩΩ?
Y��-��u>�?���K�i�	
=o���H��N Wf��I䲇�J����d��_�
��q���ۭ/;�w���1?7��>��j"�8�(,�a9�P���Z쥏�0Ȯ�n���BO�ױf��J����k{���pOEBt��	> � �k��b�5�����rز{U�� �v%4� ��?��ow� O{/u�t�.�Q|�E�F�U>�s������<�#�(-�����Pȱ���y]}>����<+ -���9�����B1�\6�&h�CÜ��״䕃��}�'B�1Y�Q7�Sm�3������������<��P�{G�{�^A�h�?s�q�Nd�c��Bg�Ba������+5�y�4��;��6.C�we-{�J�N�NW!��C��1�?�����!ֶ�;$��B�ˎ�ZN�BK.՚Z��o(o�(�{/^'�ej^&�����ߊ��+>Qv%���]N�[[���k�$�~��`�E�r��rx���W�D��F/F��� ��*ʁI&���fB��tfra��ʀ/*�HV�$�d�T56usu��-|`�x�B_@P?��^�zl2O�#��X���M�y�t����@�&<�*�wPѩ���I3y��j����/k�j l�oi)q�j�i*!�\B��t9��XH����UD(�lց�<XYh�Kn�� �� +C����	F4�l��\�c���mJ��Y�m8r���O	����s����i�><'�S��nbR�a��Nl���LZ1=F(f�J�p3�i+u�$2�uU������H,Y�Lcd�ݟ�)5����[�����]2�;݀W��g�2<xuZ��!�k�j�S���Rlß'�%X�נ�be��AP����H�I�d�d���}�+�9TX���;�(�tW��hzԒ�aE��"e��S�C$�����UH�U���̾���}õB�� �ۘu\�7�!X�l���w%�vA�Cd��ہС�L�,��N�/.��,�&�3F�gC?��W�U�٧�-����C�D£	*2e�D���dE3�m�����l��r�[�=�	=�
�$B��d����Vi�,)_�D�
�8D'/_:�ƶ"r����W�
9�R��<��oK����٪�h��)G"gV���:@=�����D�����@j"��^���-� t6�ϘS�9���th�̜���y�D�����i����8����:@I���WO���5��s�R�nC��f)`�y�PȨo_���(�}}���L��
�� ���'uιo�@Nvƴ�����;�
�\8�Aj�<����'����F���Lͣ����at����\ʷG�&���'x�S&9Pֲ�VZ�0/i�ɂ#|SbJO��M�P+���OV�ˣ
���&񑛭
�ې�o5\ֺ�&2B��|!T����V��W9H�&�ʊ�	5��xo1�W���_υx��j=Mj�[c��b ����񾲭�@t�J�:���=��s�s}/��n�K,b�ˣE�3oY5�H��*5O͓&�GP�����`VFw�m��x�^�l��[[᯷�g��!�b�榗�����~�i�Dg�0��
��vF�ۉE3	1��r��Wt��A�[��lm��9�:����<m爐�%2.,~|(����C!�_�����K_s�}�g�~�{K[N��Wfq�Wu��,�B�8"�7��)C.��1!�u�V�nhՎ	e1� ��_��JK�(�aU��-
�\�n��IgO���K����8��!O�>x���v�Tt�*2�puHy`�[R����Q��Lí8� /\�nk�L{;���th��j�(*GQ]n()�9!�X���Op�P������VSk+}�,�^�]��c�w�M��|ӻ��Uzt,�\�h�X��Rv�����D�X��վ�s��ِ���y�u��.�@<%�'C�[t.���ۿB�}1���'��R_�J�G���g3{a��|7sYV
?�=if0����+Q�W�r����>�9�_}-*���#���� M�LUS�z]aKMZ��'�s[�.%��P.�F�.u�'��� �?��iu���0�K���86!(��%�������@���aq��5����_��9����� ��q5���\��Tk(��a�]��R�a�x7/w!KL�סG>D�|�z�F3�����Iv����5�<��˛�d_����Xz����$#�`',��v�a���������Cf4;E3�u���_�s�^^�J��AW&ceA�o	��@Vn���N�zĥ)���p��5cxݼ<�N���a7�b"n�ȟ�[���T��d3��V3��=i��2�J$6[��x(�y1����b<ͼ��`/[�����	����F�ѣ�C�lX)�u*��3{�����OJ4��ܲ�gN��3� OF��A�:������+g�W���Jʉ�"b���Y3�"�i^�z���B5�T�2�Kg��r��%�ѿ�n�c��:B�lE&u������^?�k���u�ޱITE�{j��\���sn.�q.�����Z]�1���q��
��Z;�FZ�����pN��gB������1$��$"��7�*,,��LL�)Q�&D@�O:�4������I���*��N������/�N�ڴ!E�U� z��.o7��n���{���6�'����<v�_K��"Pa�t�sw�#!�'B"��o���=����Qş\�B7\� #!%��ͺ�yZ�}�TCJ���*��������Ś�w���n��0�ƌ"���hZ`�g�n]�1Zً� 2@Ϳ!Lᮻ����i]�x��"�b	�ѐ� �����P���J�fs�^Es�b:���!L��H�ݹ��U���SR�*.t��{D&�,���w���ۄ��}���3b5���Ǭ^���,���#�����x�7��g���-���j���@s{L�V��%<��8�K��E��­�#t��S����g�s����Ivr���@����$ � b,/V�msN�]>!��rn���ա�Ӱ�<�˫ &xx8f�jl8a-v�vIX������=bi[tu8VM�s0o�804��3L�=��m0�-��*��3�p�x�,�}�5��t
�BF�:&�J��[��J��^�*����;t���K��}h")n�Z�L����8����b�z���I�58Ї�濈);ᎶV���Ҍ�x3c����@�]�h�C@�^U1�ҙ���ah|
Ū���:���S�Dxm�>|����?2&�"g��j_���=@���p�B�g.p�P�M���UG���b��N)b�s�t�
���:!��(&�6�~�\�ABa_&瑞K�P�F�Q�T���1x���b�����D?���Zx�����1�A���l�\5p�kR$s��L�LF�����%��`�ν��N
y���|�|\��ؿk~���br|XH��t1��`$�Z�����w�u�[�
�>�ߋm�����zT��tXר�_@�G�:t�D�2J3 ����YE"ڶb��;��<gu��i�g���{�n�ں�]�n�=�{\��V��f8;�lW*N	 !�EUQ�&GJ� �얢q��(��slk�
��'�w�H������ѸT����
Gc������p$R
�eEA^U���ᢠy�����IV{�L]��C��h4�S�`/_�f�Xoj��C�7��ť�͈7���n����i	l (�{Y�مmm2�f&�D�A�g�:V^�{v����T�M����C)�s�Zq�'?�ŋ�0�*໷���GE�B�4ڢz
"����p�2����@���B{w�Ə~rz�䆥����}L�Ag{�����C�P�!��� 9����0��Ɛ��D&9)�f�u2����Ѩ����-�h#��Z�����lݵ;�`�!��%+�c��p��5��Դ���^xv�;��G��=�U�ף���<�/|�s�Jg=��Ճ���?b�	b8�#�����	֎+Ɉ�[ǧ5�m٥�ؽ
�.���;� ���.�d��|&]󐚚�SLCsK�TGx-�0���L�����Z��K�@Sm��9�l߹�CP�l�B0ކ�M'�&6�jyOG8ބh��'UI�b|m�\^�?��HS�:�őpzzRFŚL&���l�[�ל�t��sYذk��tJ�� �n���bp��cpם?�H_,Cp>�3d���������?K�Nv}"��e��x�\�Z��p��ٌ�s�vpzc�L�d����TO?�
�3ƚc��'���X⟿����d6"G��sK�Hb�eNb�#Iy�[�1v��	���ŊE�qԑ�p��eHD#`������s�M.�X�JE�k���9�����siijB0���Z)�S5?���06��+��D��1?*s
e�<�(���,j���Ɂ�W��td3M�֑��{�����{.��,]Ȇ��y�gKY��(z�'�e�aǇs�[q�'>��}{�y�s���_`U�u����Aȯ�<u?H�f�J[��g�ĳ��=���{}���+�z�	n��sOK[݊Jz$ccl�4��/,^2�G._��9�;�6�y_�_�'{��q���V&&o*��� �Y0o�bW�1J�뤗x�Z�w-� ���c1�ڻhm���'Ȯ=�T� �X��#���b������ő�/�Y
A��)�&,��lـiyJUɻ�K��bUEJӴ]3�����d&�P��JWU7����S(UdU0��ab6��d
��Ķ��Ѐ��f�54 ��HOO®�D�26=)�HǼy蚻 �d	�>�	�v�ʛ7K1�FH�0����,^؉�T�����qh E��F��=���W3��۸W�݈h���8~��o�ē� ��B�t�M��{ߍ�]r":w�����`b �t!���v��A}����9�e'M�KuxP�A��D���V���L=��ux�����&B�1w�B�8�H,[~$ҳE��JQ�EG4���|
��D#-��E0d��K�������Q|��M�]��ނ���R�"�'`�d5�'�1)>�J��IH��	�r��Q4#QX����&��tK%)��R��,,ݓC������m	440Ζ:�u��:͊��0�&T��kN��DWF2%�KI�$.�YV�8|E�1����b�d����1"ҥ{�G����r-,���R�QA53�F5�37�D<����1��z�`�:ο�\t�C���Ǎ7�(q���t4�#(�2r%�`%S7z1��}��H�.�-�H5�}�E��׈������ַo���_첳&�G��%L�*E��T�f�2�jmlD.�0<���Xu�2���@(`!���`o���19=%�w�P�#��~��5�g�	��Ʒ���s碥��'ϩfRYI�-}o����:����B�"�Zl��0'42����L<�	�˘[�]��֯GCЂ�9���`�����#�$�������(Uv�t���ڄ�|��:t�?�0f&'�Z%ӟ�)�q>�3U�?o�s��'����s��$��X�q�r���	��q���}��/����H����y�x.�`����ɤ�k����B���<��;^0蹮뙦�ض�+���4%Q�>n������R0�����C��,����r٭V�^�\�J���6��p�u�.�a;�y���Y��z}��?��_�=�3���^���n��k72y�B.�4�;b�H&�$�P��PZE�g�:�Pzc�X��ؖ�E8��2�<�G����yA���#���QP�!���8���V� �.R,�Le�E�P��k��+JF�6�)�~M�vUu����s`NSM+h���.yPg�U�h\a��X�7�У�5�kh�E��L#���`a�I����)��]#x�׏`۫��
a��h�����]���19[�w~xv�CA!�A���s�x�g�ӎ��8�{q������aL�z������p��ލ��!^��������u`r|#�����Ĩ �ej�[J\c��E�5��Ѧv,9�hNe�?��k�#�y�E�BQQil��EK�hl�]�	Y�@SX���f������'�A(G��<hkV/���%D��x�7����,Զ#�F�����$|nd9Kg*^�����E�/Iq:�r�%��]��UG��r��6�"���,���[ _� ���FIb$l"H_]�م 	J�=�#G	���Km���ds�$�����������U��f��˵4qdaư�������:p8�$�Й�?�ߑ�=��Dfi�L?����Л���'�c�p/�F��\r	N;�t455���ø��w�� _:�#�<�c<��Ν��|��RIư��v�D6_��������O?�}��rO8؃��t�/�cgN_����&�y5�:?[����U&�����S6�!E4��������ߏ��)�R�E�?6�	�r&�R��n����Ӧ��{sk���r5���%L�\�,d�щI���+��ۋ"���DUg<�*�e���_63�y/)��Q�<�]���ZcQs�G�Ν���:G�Z�"���3x�� ����:�Js����/��{�~�:�So��D@ 'q��[?�*�����L��3g���;��=�1�)�0>6,	w��,Je2]h=@)�U��u����`U�,��p'�էzڬ�i����zj
򊢑�T�H���UU��N�'}���ӓ� oq��<�Vu%��L+��3)�
*�Br���dш�SQ\�S���+��+@՝YQ�"��k�4����t��tWU5�UUWqU�S=#`8:���y�g{��UOS]�0T�qGQ5��tUU�S�?2�UOU]SS��C��V����N�=�寿�Ou���~cϖ-�#�� f�mU0H�����f<$i_rA�&B�8��L��t�(щFE�]R4�*r�����czjV�@�1�,C��܈<P��jZ��MS����Lð�U��+���̀NtvU��c{Mw�V��\�6BΑ�ˌ��>:`E�2��@g�7s�Ɛ�|�5��TG1!�ף�b�����7H*S���0|�^޺���¦�c�d5���|��X���6�s���g9����uKu1�1�+.9g�\�`^yy��o���d�fɈ���y2>pٻ��E�#J�M����,�]`rl��C�*�F29N�	�3��C��u3
6�:��:�x�j�O�1�*bہ~�������xV�=�B�398�����Y<O>�0~����XaM�Xҁ���WikƎ�,���O ��x��-L�\8eߕK�e� ���<�M��:�G�V>IG������IJ�a�Cr��oW(��������FBF~L�BR�����F��BO��!��!>��"�T�^�+�aྖ O;X���9�"�UN8�61'nl��z}��F�N�%}��c-��(>˽�D��@oin@�;,�2��e�]"z"�(���Ȉ��$X��6��4����6'KQ���JF�@0$������4%	��s����8��o��/>	��L�T#�͏�+YNUw�\ilQl�<�x��Ւ��A<� �={�K�#v�U0�.����rGNFX�����>��пf��W�+��}���X�h��^4_:�?�?<�<���B�[͐��k�9�v��E��Y�ܫ�C�����z����`�����W �`�k����-ؼ����F��y�����؀�_� �����)�Й��뇯����|~>bU3��s��³���9� ��׿���uu�)j<49���A�L�a�ף/�S��AYq�æ� o���Q��7���'uҝH�j�"�h���|ԭy��!�����ǩ=��&�G��7�g����{*���������/݀JF5�<rU�J�'�h����O��&i�c��~��(���;+�h��*�gW�
4����`$�s~K���c������������Ɂ�U	(����(�aswkS���T�&�w!!��K�*���Xf�g����v\�m[�z��#rAҕ�*?T�/	��hd�u�x"}�Z}���X8{^ūTX�U�R�ī��Z�R�غ�T���f�F����u�eG�˕9%�m/�'j�Aa�W�iJD�"DJ�x�S��q.�G�Ñ8��FT*L�
�Nt4��x�l��g7m��/�(���W���?��X��c�6�}���Y䊁]3�Ґ��9�ኋϏݷ    IDAT�y'�؟vp[_�&���Ff�xg�v>��K���EA��o<��}1d��tzr��)LO�H��ڲ[����E]c;�J�cŮ��h�jN��g`/���D(��F4�[���bp����YS3h
��>�֐���0���S�]�S�҅����B�	l��[w=�Ē�1�b&��fK�/����H ������jv]�;9����7��E��rEAnfF��
��-D��C�,*d��ޓ9��X@�$e���Z3M�vu��O�\�l*�b&dsŢH4�H�^:���s�CS��
�~�N[�E^�����DI6{�Cg�O}�.D2�c�7 ���R|�cnRv����g?����\��EcWF@�Fb�z�O�
�Z���H%��q������IWb�S�֢>]I)�c�C"Y$����_ݎ������dJ�I?G�ײ3������ɉ�RaIcPE@�|��}�2Sȧe����`|�/Dx�p�`0��X9G�5��:��YB��' J��q*	G�9��&�r�j,]�LCW�B��Ŧ-��34,[�ܩ�'���h�;i��v�����,�7��U&�XX�Չ36��ǯG�0�i��x~Ӌ��NF0�͋�4�t�J�8����������:�p���>��d�^'�����s�N0'g��v6E+W�ĥ�^*^��{C~��rF��K����B�iX���{�3A�N0
I�����|Y���~�|��W����e��/Af�L�����:��gD��R���WD_���'���_��u��ڏ�F�<�yD�1�Wy�ձp�}��X�,e����tq	����"۶�X,�y��E�-^�����֥�����w�穓��t�-[��
�:HXS9��o�@$�ZU���Z�U��aY�;G�⻄|6��|Aؽ�&��,MMxCq�70()���V�o�q�Y��=k�m�5l�vtL���ׁ���Xv����;�g�����nr6�D˰$x��� �J�&����{^uh���� O��w���H4�Y&Y.!U,A	�p�p?y�w��M��Gએ~�V/��T	���`w�0ʺ)��\t�KG\wqŻ����>^a�����;�C2�F ��)d8������ۅ�H�8��tۢ8 c����^w��F*9��� :=�i_K9�}�0���t���Y��)�p{������Ζ`�0k�X��,\�#�(���h�RJ�+a"��QI����=�b� �������g�ښ��'��}	V�j����8(�b�N�w	c2a# ���?��x3�����(�{����ζ
�P�W�K��	�^}�����Kg��#n���h��Q�¥�`��~�d��k�J��Դ�3X�67#���P,��I���-�U���bɟ�h���:F��@�M?��G���������$?�E�I��u�	�q�������~���>��r=�]�V����ͦX���yH���]�m�()����9�)��AV�
1��m�b��y�6��׏�N��D<e���Z��R��aP4�4�X<_���vw��<�Jb��ػ�51c�{�b����y�F=��'���_�{�����eI_���{Ir��*,�倇�ŋ�bŲ�X�d)�+��9��^܂��u2���L*��7�%����rO���̐�2�uG�ĥ睋���I�Mrf۷oG�P��,[��Q�6���=�p�D3��K7|�vn�c��J����Ȑ�k�ȝ�'���Q&)5�F��q����(1��:��������&73)J�ёdӳr������|��k��Wp�o�_���e�.�Rb����g᜘�FZlykV����Vi��������7�豈��Ss ���_�_/4�Tc���oj?�͏�{W|����od��r��UP���˼>��.^��e��<�)����{�YY�������i�3C�*("
*�"(*��5n�M_Kb�M�����w�&�d�YMb�����FT�X����vz{����}��M��>���]�9��8�9�y��������W����+t����l�t����-`Y��UU��`M�@��ػ��3c*���̃������)zl�+�4���Etjk[��F��Əo��7m����}��q��eqFl���7��W^��{��9�cb�D�Q���[(���Pա�Zf��_nj�|Z�nt=N?�C1����*j�!�9X�0�������PF�q��1�ꗾ�Y'OE{W��������!��b�P@��B��r�R\y���iӛ�ͯn������ޖ�s6�ⲋ1��NA�C:	۠�4*)t���z`/�z:��ٮ�;5��U�׍��z0,
���r�+�i\�M��}Gz���Պ��z���0P�b��騨�L���p�rC]�PGmȅ�_��O<��T�A9�SO9����SY��w��'�D�SqhЍ����c�jt̍���Nb�Tc�r̉�W���oC{���[|�\�  �\^���ɓ�����Eo&)�b�M����S�&ϓ�
b�̙��m�]B�@w��� �̚�@$�he�f���8��g>*ٱŬV$HS�K�K�
ȘdJ��˫�N_�B�>�FX���l�3�{���G�kK�:�P�w�f�<�9{d�<��M�
�|=G����)�4ǈYgS� ����Ҳ<����7�����s�7��B'�+��B*��SdJ�B���UQ��tf7�LJT�];wHَt&��ЩY��+Lb(�-��|UQ
sa>�4ދ<t��9�[���x-�L���� !U
��w�uk��j��*#��@i���t`Y�d�!��柆���]܊E	�Db���hg�-ǭ���+��a̟�Y��m���y�|�U<���2y"��nz�L%�>����0�-��9��^��@8���[�I�Ƞ��P6����8�v��H�)�e@����{��@#�C�
�\�0�x<��P��	�,�>��@o���]B�ʜ��s;��Dͩޝ �jY�2'�%�����Ȁ�������.�s//�S���k�SL���/��/��,�C�'L���N���ƫ�!�c(��z,�*� �r�tiGf�9t�xX2C�[�n�{z�^��yfS�1s*Q�+OiQ�f<�(e�������R]�xL����[�MZ��S�}c�ֳ8;=�����3O��Ic\�(L7���������C)K��!��J$Ԟ������<�k�_1�q=�э�{
m�ە���/	�̙���~��c��V��d�RF�,3�|w�,]��\|>�B@k[V�w/^��"�u�р������a\C�@q&%%�n��VZ[�!U�Ii��N��
���<U�L;�7��!���\ȖJh߂q�bOG���������NI�
W">��x5�A�X���u� �l|�q�:���^��V���Ӹ�s���x��ź�r�R(�{ �B֠�iZ" �@�9��x���4�_Ӫ��g�t����������lsZł�Ҩ؅Tц�|�L��C[{��u`h��-�%��#�I�\ġ�#���1���9��M���#T�@4^�L.�=��L�lcv-�|��#�Ts�>l��}�l��:UH�����G�����zq��y��]����6�@>�@0��
i�������L�O��m�usF�k[��z��϶4K�8��� �P�����Ѱ�l>7�9��{�����\���p������M�%�U���7"90�Q ����k���ť����L�h�P�2o�sH0��Э�����9�"9�Ԭy��g`�)��SZ��cضk��G�1�Ϊ�C?��IT���:���O��c��Z�D�[;
�lZ�5���5��r��N��u�~h;,-���n����ǿ��W^�㏮�!ۀ�$IP��~M`���TL� ?�N���̙#A&F|��x^0������VtiC&=$?Q�(o�Nmn�!u��ۦo\1��>�;�x�m/���˅`��
(�)N�\��x��<e�)w��ѶeY��zʔ�s��n��/��'t����d�v{K��E��-��ssR�v��.7���[yDx��kܝ?)�V*�	d4��3y���r��bҘj���u�[}��.��:I#��y��a-[�0��v�#��M���<���;�?Э
�P���*�lǚ���ά&8����ȪH��.�ev��+�缍�������`y��L�2��0���\ϡ`0����ڧ�U%n͛��Gn��ֱ?�N=N7��O��:��3����AM���DA7g[�B�ص{�2Ա��E6�#lf�e7�n?��wb�O��g@-ARe����;�x�8؉�x��/x�����~(��K�1m|#��5��do��
��?n4�R�j�\|�r�5�T4�m�6�E��E�������I--�8r�v�@6=�ޞtvAe"��.}�CD�S�6_@�"f�:��G�WV�a�d�f�x�@;^��>�ڱyO�p����?K7=��L8m����"��|���Iu1x=�u���1k6��~��ܵ���9���hΒ̚����J�#���d@7Y�َ���4 :F�ѲG�*t���/D���͉Ʀ�4�����I�V0[��� ���5o�X�[9�d�� "�L��s�����F�q��{4*��g����&y�2���S��0
�70�\j�{�� �5�(����x�U�"R�;��u R�����G�Ⱥ�ع�=�.�m���7�R������L���;l�"8��wn4���y!(��x�P��ѐ�芛Â��2
�5�<�o�r�%TD#��L�����a˾={̇��g��0�F�Jɡ�W^L��Ӵ�
�J�l�3���y��=�ɌI�B�F~|?��7u*�_~!j��0��bǮ�X���8�э�/����U�۞�&A�S�6H�tc�qS1{�T�زEI�ܹs��������� �B�9Lׄ����x��������!.3<���uŘ�r͘4�}r�A�Q8<<+g�v�<[ܙq-ٺ�9��cp��tҦ����P��D���P�Ȥ������'�_c�T��x���+�b��"���/�w�}>��[pәKKT,��e��������A��0����t���<4-
=�r�].���w��`._�K�>�_���|���)�U
J"7�Y�����^����r���f_�A���\|%𿋡b�q^�q3?��O����\.�K�+���b�#�HTl��f͚��qJ>j&�gYV�\.|�Y��F$����kk�%D�J��-�Ƌyeڬ�C�e�k����|����j�	s3��h�1�ݮ�H4������'��izw���<���m\� �L������'��C����)�0.E���Ԧz̜<�����ěooݨ���PX�>Z�(@�A��o��Ͼ��������k��y�N����r��vV0����Jp���x���[_�"fO+������~s�o�& �z���q��2�����<��ֻ2Q�SO=ɡ~l~�U�����S�"rzy33l�fWEaO�4�
����E��	h�@O� 5��;�!oy0jtb�
4�L����~��W�Rcjxp�x��W�Y���4�d|�_A���2��mk��ύ�λ])��?��PF��D�+�k j+1�o�Х,g]8�{Q�7(i��ۼk	V/�B�}�J`<?d�B4w1/��2��6���O�qߡ6�IAu��gFkf�(fD�Q��OT|�t
��_�ĥQ��U�x?���]T���
�l ]2�ଲD��n/�
�9T��u�'�w�,��D<���<�w����,��h<>�4%�"�V�"�-QJ�r-u��Ix3�%����<��R��Ov��CO�#�8���n7�� u�C�Xm"�p���[��Q�����G{k��9�lYMF(r�5�n��6�c�s[�@�D���}�a�5���z���S7�������}�bL�z�
�'3xr�F<��u����G�� ���[��1��Eb�R�Sƍ�_\z1fLl��n�FUV��.C Fw� SY�j=�G7<�}��3]!����oa�����uH�R��Tģ��3�`"��ɴ��ڡ��p�������u����r��M�N �2&@�
��d���$@x*�~�+;s���,\x��>{�9������s��M��匿���[�Vy6O����wo�_>����k��	�P�`Е��F"n&'��~���u�G�$ŗ��J+�͖B�ѣGg�\|�#�sв��&˲j��.���A�Pqd[D-<��ɜ�Ʉ��'nl1���l�'�/��+
�xX�:����Ʉ�������r���w<����GN���6u&F��ǺG��m����0�*�yӦ�)@yD��=G0��a�G!�.c�	���^��xCQܿ���}r3�Buu%���pq��?��Wز{/� ����b%°
J.9�\�b9*�^�^��<n��ϥ:F���3�c��H'��"o�7��>�V-X�s�lD��޵]b=l����e��%d�-l�	
#ҹ�F��͓��'���C�xo�~� :?��q3N�ĉ�Ma7 QW�%4#]]�_��F<��E"D+�������H� ����~y��cp�+П�)���:����F�����*�쿢t��SD:"�m�m��f�D���AG����5y �!L��|zy��`
��3�I
t_k��nݖ�|0���-	.`!�hs�y�A�׎nh���42ɔ�c�ٮ5q�T蚡���Nl ��Lx)ܤ�ƌ��V��J}��AxS����yb/����xs��ꜱk���ɑ�11 S����`G�ي�d:�$�&3;�w��1�F���b�s9Gv��,�A
CR\X%T�"�:a<.Xv"~����oذA{��'��<Ї�
^{ɘ� f�������M�vb�sv
%�R^Ke�}��������ƍk�i���q3�Wҽm�.�{�)iػ�Q$�U$8�Cm����X��� S碥�`Œ%x��xd�,Y��\~�|�m��uZ���[p��G��k���fPʥ1q�X|����;����Y���
�2����@RI��1akB|��a۽j<2t6�Q�xJv�Ώ�M`����SɻE����=���Bn�I�n�Բ%?���{�������q�@	Xb��,���q��j��������S��bF�Kkn�
�lV\.�sy� ��(kCC�����Om5�H4q1nL�x�g55���r�����0��v�����G1��Q�؀G���@q<pbn7f��G}ȏH9�@.)�MS����HW��f4���k���3�U��z�}+ї��[����Ѹd�r\|�
��~�7bӖmH�3�� �
"��yz1c�x|�3��)3&Hʵ�Hn��/����;������s��@&c�p�%�v�?���jk�P*%����f3�K��c�|^�)�o��l�K%*��<IV�Gzq��[-g��&MB��	�=�& ��"Q��&!�� ���;��3/>��׋E�/�g��ETWT��}mx��Mx`���LĴ�K��W��7��'*eU�E���0k)�� 7f�Fm�!��rh�fo��X}H,øjLAA��>;a��lZf6� �ǌy����#1^x\t�c`�d&��Y�#.x�DF��F�F	.��(�P(��������d�C��M��H���d�J��4p �|�,8U��ۈw����x������#�1����)���`N���{�d�ܝ�.@�g4����sg��i˳������E�2Dl{������؆:�cA�uaժUɲ��t�S��:I�G<�&Y�)ˈ�62�k�^*i�Y��bQ8����A�(�H\�������k��󓝓Ó_��Ͽ"H�JHSl(N��J$b�+�!�|�>�Ic���%�%1    IDAT��#���/�9�,�=�އ?l|��:	���'6��'�@>���K˘1���k���7��c� K�|����
���C_:]�Bh�V�H��T�V��1lq�eI�5V���);�2����Y�E�#w�T�1m���/Z���d�c����O9�G@����(� �4�p��a�=;�k�}����U�X��4$y�񊫚��N��U�9'�<l�3��T��r :��&���Q�o�\��c����u��k֬���y
|!L?�4�o�����杬.)�R��>DC<�ۅ����	I$vtvbTC=&�LB���x=�?Ё'�ۈ���gL6�2�嗬��_���>�����7�نQ���-7�n�
4	{]hU�e�-�K�C,�`d��w��]w݁�^}�Ǐǉ�/�n�G�ML��lA����#�)scc:4�gfl�>��`
٬9)PJ/�lx�D�{i��/��[�}����_>ge,¨��鐩�U�cy�����Hsh�>����0q�U�/��6n�gv�7�N_��7������E��wupSpeD@W���J��F::+\��T�}бu-/���8w�h����d��.[����f�a��9�|>l�@6o�*H�߶�ͻ�RcP��@0���f8^��<H{{��3��Z�&�1CޔSj�����&F)�(w:ą���Ё\����8�������ؾ�]��%���/�"�I}T37խ�d0�;���9��T۴!v@�?�IwP���i��@^C��]e���vs��C��Bèj|�k_��`$��֭[�~�z�~�'9�e`w��K�2GQ+��X��Hٞ�ˡ|X �t�5Y����"����d2=̷�C�rV�S&MV�y�$X� �پ���d�n�%�8.	`�� �R �&�W��sh���ݿ�z�t`���p��xr����[8i�\|��_�c�ã�=�r� �q���/{�o�3O=���>������p@g��������8A�i�;47'2��Y'���E
�d%�C��(�x�^���L�Lmn�cɢy��+�9�s���~p>���"Ά[}�
q���&5e�N0�x��K3��N�����h,�D�b�Zԑ���AI>�Y����E�R�"�jjb�p�"��r�Wo�2��5k���q�	'��	-�r�jikSa�T�"��2�ڰ�B�!/�bQ��ǐ$"��q���0vK��W6��w��W�&��XB��E����^�O_~����O���V9wѽ������-������0�:��.Z��.T;��?���yS���&rD��r�Q"��%��lZ�C� �M�6Ѱ�JZ_�(^TH�"��5�a��4��~��H��/R3(2�G�uOjL0ĠQ�!��������Ԣi3���y�c�S���ݵwܽ�x��hx�cƂ��W&=/��0NtJ�\��(��jrC�]�$Vbkҗ)3*MF��2m[K ��n4�ϔ�#&E���Jr�#(.�ϖ{	��q�isP�y�0FQ"j�S��'p�97�D�	Z3�'R�ҮE�K�Q���A�3Yd�E䨾H�2����$|���n���B����>�:v:��=Չ����m[��T�
�`Q���@I�F\1����p�.Y�9�N@?:�0�XӺ7]��S�s��D���̐�sg��� ���������cL�3'�;-c2���u4����'�%�.A��y���Ιh�#�yGV�1'$�R����;�4̟w�\����;�ġ�^�]>$y�Qh+���-�3iDxn��K.8��x"�|�E�|�=ģ��{��W�q�yK1a�4�~�J���K���$��n���ϣ��<����3��h�γ��8�������J�IlF��#G#+vg$���l+Y��!��~d9ZF᳅y.�"�Ǵ	��,]��;7\z�1���r��o|���=�5,k��R�+��� De��ug)��5��Ψ��J"C���HD��5��Ͷ�tǍ���1�yX{|�e��áu�"�k]��!dď���2�֕�W�=�uA'͚����X��!�>����u���R7
��P�
,��`K"a�J���7�M۶aO[;�$����� .[����Rt��'?�w���(�������h+�B,��U@fh sO>_��_aڔ�6U�8ҍg�z�vlGWg��F#<� m��GU�r9*b�Ԏg;qp0)P/(g��T�bW�����k��uM����`�������
�-�ߍh�U��d	�\!�'͝�N>	����"�:�����G�@�G)6��)�2o	�\���!�f������ˀ��L��
����Ht%#�SH?\��	f-:+�}�	�4 ;v$�Wv�V�c[*(*ZI���1�0�d����űX�Jl{��.��C�>?Y��r
�4?a�@�q�]nDb�H��[1���h}t�7j��m��"�DDv�v@���b�}+b�>t
"=������ۆ��	�i7v;լ�QP�/*�P܈��������3��S�a�y!��s´�MK�@8��G)VS�`lM%.\zF�T��"����b��U ,@ӿ��93�olX�x�H���5Q���eF
L��ȪөH�t'`��Gt�[�ǖW���!NN��#�PĘ1�b����(��x�g���1D�"��X)^QID�m�+�s�<�8,[�cG��L��ؑ+�TK6�˛��}>$����'�����W�p�܆��q䈸��f�̀.�Y�&�a���m�Ff|�5r����D�禺�O,&,yZ S��	T(�`4&�'A��S�5�Z6�7n���O�G�I�a_@w[7hVy��,��~�%��;�<�\V&��@Z���9q�M��BI�v�����M����R�4_ἆԕxt}$Vqm8n=�u[���i�ܻr������j�r�\L7>�Fm���кe��Vu>9�X���ۍ�X�dJ���(����H�\,!)��#q����������\���/���#�ɏ�m;�����*y#=XB��;��L�B�Ι����4&��� �EOgrh�� �=�����i�h"��HG�t.k�_��{�v�@GW�Z��:&�;���*���
��\�qM:P��'@v,�D��>{��0fL#r��$3���� �?B>���r�[��A�����@���"6�d����@-:Љr�C��;�^��c @#�'��Q��g�h�kt�*.�9;�y;�c�ߍ�������ce�Z$##������i��u���&"�ّB�04y��$��W^J�4���:�ݽ�F��4^Q%×!�w�hj��Ra�2ү�Uq�a���R�ba��/�!��`�mV?.Z�P�O?�4���*�^c��@]b�$r{,a�88�o�6�P�VS(�F���ٶ�.#5�$�=���ۭ^�ws��g�0nTV,;�rR�aӦW��'�ʛ�?�ωng �n:�g�[�<������I�@R&�����s{�H6�[�m��|W{�����?u��8�a�X����1K0*760a6�"U��nW��ô�͘;�D�kl��2i�e���=�x��W�����%�A��4�T�o�~-B76<�8�C�8��*�z���O���w��Z�l��:�`��p*x~V7�>s�{��%-�bQ)u
g�Aݱ�e��8��a�ئU�,:��_�₶c9�?y�W���~�r�~��������!�#�\EJ!��QE~�JR1^م��Bf"�
�Ɖ����8˔t��*?�HT]
����ͭ��z��U:��G+��B������J���Pϖ�R���_f��C��B���?j^Z(�c��ayi�b�=%���C������UW�ܳ��H?n��/��[�d�`y�P�����B��LZ��46b�f,Zx&f�h���`�pڂ|F���S�L6�h�����uH����W����oDGO?2���	?���x˘F|�keg��>?��o��>c��Ϧ%����P�ǥ�m��m�č_�f=^|�yͩ��0�.*F#?j*�.8��*d-$��`��:�)�� K�W�L�Σ�ҏ`�*����0��l�ٹ�GU�4;/4� �~�����:YA���
���g�$V( Q3
Mcǈ��74����L�(@:�NP��
�����u����ƶw�#�4z�x�\��9I�2I藈}c+����.r apD.�J!W
aw�@+�=�p��EH��x衇��[o{aS�����ǘ�H��6����i,#���P�Eɉ�(h�@I�3oKb�:��1�T�D�D�a1��� 0�*#򢹩+�,FuE�j*p�-�������7=�^{.`�ڑg��� ��T'��xe����hw'�i��7�AS�XIpMXx�(ߙ�(L��j˓����?a±8��s��~�G:A��`6w8��[N2���|�P5˱1/��-F �.C�<�Q�\,
Ll�Ƿ���엟�i���[(ds��7c����&W�� 8�|t�r��xu>�w�IikR��e�L�(�LgO�o�c0O�Bz.H|{���5lM,�qu�k/9��뮻r�1uN��L���؏'��X�u�p�����\w����@�dR)Q�B1Ӯ��Z�DU3{��ll�FR�*����D㱧����{�rWoz{��+Z���?=����ŋ�%��o��"`���P�T[�\jBNP���sI��$�he�(C�Ŕd���/~N�����q�/~����G��`�O	X%6��鐳��܍ ��&��'b�ɳ�2�N�d.=�Y6�j)4��N�]��%3wRq�3%W�n`�~��X��'�F oh�������W^)	�(�ר('�%�Ea'I��mZ�l�%i{J.7���,w��a���B����{�� �SN��9��"ח�tAܒ_/	WV�,V�)lb�;�?�!�`=l�IFXw�#v48/�4e2F�T���{v�Q5Lq�g�,�(E�т**I����h:;._�nъ֡�q��������:�t�EJ�vuM�(lL��}�e�)J�e��[�LF�tPV~���[D�M>zZnk�ۍK�.De�b8�;U��2`'�v���@�ކ�RL���W6o�V�s��ڵ�茈.�L>D�_��Fl8
sT|d�� �"~fN�����#1�~���	��d�*�Օ�
�蚙�l����Q}n�=r��1<�?j̡���"��(Ζ������G�&�4WPB�U��D�s��h1�;a���Zۻp��u�r�}�fSE��V�Ҋ�#[y��gGM"A����.�d�2����>�)�����|�kx������4"c�k`��q</��`���p737��p�H�@����@�f���X��x����X^�銒�h|��F�9�ȥ�.��'�X����З�}����5��ٴT��r��T:�G8�;����e��enP�Bg�/��0�(���h�ʊ�o�#�7�e�x����\���֞�)�X/[&0�ͷܪ��\5
p�t�,·�<t�o�RU���(RN��ʄ .�O��ݻ��7ߌ}�`9jy�e��3�/ZizX���K�Y�-��[H�x0���M��D$��cc;|�b ����P��HI�Ja���5�g&^�k�a��P�"G=�&��>W.)9 (V�tAf�����N�B�5�����C]��]h;�*�;*�5��!���/o�p֋l�DL�>yГ䬕Jml�䴆�� vln�1H`�����/8w�&��f7�$F ����
�4{z��عs'ҬDT���ٓ6�Cnv���2��&���i���R�Q&rÚ���k&PU55��UEɪ�IR�`:UB���}]4#veZ��<4�!��#D��� �={ɶ���MMP�ۛ�6�}�KcG ��{���WT3�BN�}��c�B?so���L� {���n��*C2�e�a<�=L|��(XB��z���hB~K��λ�(�����W�c�e���"h��?�mz܇��hƙ+���؟� /.�F+%X�|�t�,�P�L*�\'ϙ��Δ��`*��W���{������4�����ҩPz���x������C�VTޥ�"�>�,��4��*��o]��p ���<��>Y��O@^Kr���C�N�v�+��8]���w^窚Z̜u"b�8^y�ui�Q#$�;�@�� ��CS鯀�H ������_���e�4
=�3��c?���Բ��r���f��|�D��#�L*@�
%xUu�FU��+��U�ݗԖd��	�ܸ�p��x"�p"�ڱ\�{�}��k��PO_.X�T���w݉�~�'��_	,���p��}
TV �Ɂ�C��g0d@��g?�3��}����_�
{����Q���ۍ�N|pK�&�����jq�<L��buA�5/���*o�B��!�B��%�y�?g���6���eEQ(���eQ�gP�H NA�b�P�R����t�Nz���@erW)�B9iA�с��������U�Bt�t�1s�����F_�@"�l�5^T���.L�4�d@7�E�]���OfѺ�3��<\�q,��@]�����66��4%��Q&4�a<���Ji�\]i�q�-��oٮdG�G�.�J�2-N������/��	��
�酳�%4[ �U���m-�ʣ��C�{/�ø���2�y�G���on����n���z����Q�!ړޟѮ�r8c�.WJm���1)ە���S��8fq��D��zq��31���%��J'�j��!	�BODcJ¨H&�R;qt*t�k��U����?'�+A1C�!+t�b7�8D���jA�,4ȇ�����.?_ݬ������¶�Pd27
�pހmdB� �|)�=���?o^��Y�a��=I|��r�rUA?����FM<���n�}w�)ʫS���ý���y�<8���9պpv�ݡ�)��c�ǃ��-�Ԩ�i+��}���a E�֩�0���](�5�����E+�}�[-9t,��'���
|\}������>BpQ�]�H�Id���d����R�B�3�`����5si'�����������kB�ʏ�`�%��ɗ����w���7����atn��V�Eqv�j��Z��b+x)L��nWЪbt�[�
d 3-/&(�g�RW]�/}�*�u���u �y�Mؽ��r��o�p5�V��;~?fN��)�-<��!5��UsKҺ(��r�ގ	+"�M��t?�?+��[��m�5*`���g4���Xzp �.:�|4ԎB�>�T�(#S�IZ��Q@������]�1_+U�x��k�SO`���x�V�b��Q����gcg'�)�$,����ڑ&@���6�x����+�ذB����l��B)�e��eT��
HЈ#�U�5��	oKi:����u�4���
*x1��}k�����Ӡ�y�,�a��G��)������V���ͩ?���ʗ�y	˄=��G�� ��CX��4��}�Ql����j��:I?����w�}��3:(wG�L���ƙtx��K��v���-ɣ��2P�Q	 �-c�)����׃Uk�"�Ί9n�I�*��Vg~nRTs'�Έ馔�=0�ć���4�Ǧ��-w��i�J
��%섒�@�sV�3f���.�i�����ޕغc��:��NU5�mI���>m�!aql���̹�}���tdu�)��y��o\��ύ[�ŝ�ޢ�A0���(�6��t25�G;8�$��Ȁ�}�8�<---UW+������7(g���/5�GQ��AZ�R��xȏ���'��h问�$��Ys��#�wŀ�����N�,ݼ������ ��Sz�i��Kژ�B���S؂hTrv�AUe�a=������>�Hl8��_=�����p{w6��Dq��'��������(9���H�S���K�8�ԤA���{�=J:�d�ake3�s�\?�
��Wb�s�}�n����p��S:�g��i�=��(�/�Xp�l��gR\�d��R ׏�m���Jf1����$�}�}�Y�x��M`��    IDATV�ou@`9�ċ���q����~�����-d��P�aa�l ��<������(	7�<�� �~��r#n��o��6��Ig��fF7�ڊ�"�����qX�s�ɪ�����[�@��G]�+��QМs�9�f^#�,QV����TjH����� ��d���c!,s�,E��/�k(`�����pK�y��4�/J����U��\&P-[ŏ7I�0%�cf���g2:�]�$������NDsmX��Tɗ>��cx���$�$r��5�	x���-�JT?���<�k0B#f��-+5^W��;ռ�O&v@'���+��x	�t�o�q�'bтS��v�׬8��2n�8��&`1����8���9�-�W��	��o'_\K>�3o��
�>f���89-t�)
�p�p�EHe^�з�٧�c�8�_]���:�J��K���J0�_6�A�a^v-gR����/������l����7��c���&z��Fw:#��&��:�S�t��������CWHR(;�zp���@T#4�Љ�	D�U��E��h؏	�MO\v�y_��B����Ŝ����ikc>\||g��s\b�AnpH�S18R�w�xY��{:h�C�${v�C��?ؖ������TW_��|�����}ܴ��%k�}��T��	gϟ������U��o\�ק�)og�h1կ��<Č�)*9tbW*��iV�W��墁�|�@qm�j��4u I�E�[~��\��u���a��(fy��N�Q-������`�M3`PN�I����s�e�Aq4U��Ťj��{�wlU�`����~T�][�����R] ���c����b��|���p\y�j��Jln���0y�!��i�� �M��]c�Y+�iG��>�q}�`E�I����7y��c 2�6�9�_un�Τt �
F�, )^�	�3�Q����t.͔I�S�-�.
z��U.����<m@���#4�#��[�<����.�� {¦W����K�($�K:���F���R��b�,9�h@�W�(��\uL�]r�v�6\)��h������JmԶ���V�$�m^�T��/���9;G�T�Fh�[*#�"�VaO�O9^}TE��]x��1�L)���!�Z�i-s]�7���FiȦ��V;#'��}�k��`��F�s����M��dZ�sR	�#����SN���ːg�Ofp��jlF�G�U�l��cǋ�Ö�UPeWM"F#�-[�EH�w����~��4׏��~{�oU@O��45�!���{��
R���fF8&g���;:#!�>��H~�;�O׷��!(�"M �;��?ǁfA�0����+.Z�I�����?����Bgr�e�wf�����':\>#�69��<Y��,���Q��Qh��7�F���:pU��04��`0x����Xu������G�]����h�j�K�EK��vT5����Y�l0��:d�a �o�Q�T�Mf�4���)��/�D���ӗ�sc��ݸ闿ā�#(؈ $�����b��6����ۘ2�QB-=�]�3=�ۨ.�l�TDe����jX���Wm�B���Ͼ`}Cx�ŗ��WQr�D�	�8hl2����&�8}&O����z� ح{>?�V7����b��.�_�^Kv\&��GSC5����~��{�D�LA��3��=��~�F��c` ��b��^��VVa�L�l_j��C�-�+�2�ܭ�����DMu�#Y�e�D��݇U���96G�s��,[��\�R�t�����/Ic;��H��E=�~�����:���)$C�9㌥�J?�L�M���y�UB�S@�ЏEg���Q�j������S�tUK��;
�\���M`+�oS�t�m$���fP卒��\��Ίր2M�%끸'�y}2C�ra��i8u��h��T����@Wo���رc�ET�3p(���,�K����n'��'7�A{׮X��N� J���̀�
z��\�w�Xtι:�:zp��q��C:��r\'�8	/����Ά�9D}%��g	��m̨�6��rI�PD���g>u	��;���B&+� ����׶Q�����݇�'5��p�ޜ䒉 �"���,�k����;�+�M C�OE �@�0�eDCA�k�{���/��w/]�	(���?����<�*��p�\��:,	9"V��TiӉBV�T
6��$&Sb+�3uJ0�hOU��踶+sV-���eK>:TYY������.�ːH?�����O=s����1�p�-\(������M�GP1ϲB��"�h{V%6�S��2xئ���x�C�h&#�.Al�H_���p����v����c���H�JB�˺��*����<���oc��1H��r�������k�d�I~0�[	��_�`����M˹:�vJ��7ΎC*W�����}>�
� D�쎔�{�����	>\���Z���#��!��c 9���`O�BHY�5$]�$��/8}���/!�g �{�?��V=u�[f`0�̘�C< 9�h��U #�.�K+�0�i�g�̄�?��"�_@jXe�s�S����T��R�j.I�h�۲�vP7զi~��eW3���h��4fh�P�� ���c6m[31[����� 2�!���ǘߡ����;��LA����Z� ��&�9��B0ƺu���/Is?�*�	��5�ks���|P����٣�/5M>A�
%�Njh�j��73�q��,�k"år�PXHl��Wb��P�qA}E+�-BeԏH4��k���56ae>~L�֋�
�𷅦l.����0E��DܩL���n�S�:kʄ�Ii�>
�8�a2U(�������`�
?�D$3y�ؽ��?�d��~?�Y�Х�j�}A%�R��Ed���#5>��ˢ$oά)�͏bz@3��h���uصe6��	=ݦ���@2�[:{��<0��r��Hl���ذה�g��b��gG^���
ǐ*{Q$�$^����/�yL�#W,?�k߼b�'�2!�������y˚��u7\������Wc(OҘ��,��4�E�BV��[��pe�ꪂ�̛$-r1sK��e��M��m����Ne]�:��E4�G���ɗ<�ؓw�����Z��Є_��7���"�lA�Q��T�P5��׌��s�6R
SL:|�G�Ă�H�М0����/p����ލ���غc���Q�c��
��dd1~t��{��Թ���%|���Љ!�8;�^f��Є�������̲�p�xH�&4�Q���@�N���g�����C�����ۃH<�T&��&��s��@/"����@��T�!��q�'���}L�0Y��5�ᗷ߇��G��N<�T�hi�K����q�����loC��C�>Үk@���#2��"�#&�ҫ&Q��0E�2tT�3ֱ�К�����x0�2]����j/ۉ��L�F��M��k���T����<��Nu6+{�r��֪�.vD���,�D�-_Qmw4
��o��m+��~-a�f��E�1�Y�o���.>�������=癰���c�),�7`UQ�HC��0G;T�^�����ma�08������XGa�OU��+��)���7��_��"��qM��J٦K��&@a�S����Ng�i�;k��V��RQҭ9�����#��xh�+����*��^xu3�z�%dK�Gg4$����W@��(M��)�faْs��Q��1���>6oقW�xKl����F��o]:����?��íH�Z|��Нn��=�ǌL(��� ߇��#��|/���Ǧ��@�"G�\�����s�%bQL3v�e.���~",�"������)�X��02��'�[��1֛��l��7L�VSc���il��m��|���6�ժ��S���m�U߮ihX,�֧_���G�:�?�L�C��c����}��%Z&���&��Ty��H��"a��Q��t ��@'y�����FT�Dg
9N_���q�Y����?�����-[��DbHfs�ry�����T�����a��&��y�{h��UA�y��o�fD����j�n���B�2ި2Ղ�l$�1R٢�*J��9Y��Rbe�֠]M����Ul2�WEOb_� d
E��r�|�,
�=pg�(���f�kւ����
��_�-Г*�޵��ֻWJ���!_��MI���"����UW�;��:N9q�@_W;z�:��d�	T����V��>L�Ѵ΍ǳ#$B�3Ρ�BG\�4��@� ejߛ�ο��8Jg㕲U��Mht�f�|������n��*��R5o���j��񨭭�� ѐ���=aF	LD)��dD�
�EdP(h�����2i2��o�ܸ�۱}�.̓��L�z�#*7*�q-�W!��~�&Y4�1>���	 &!�GNv�.�I�䜞t/���@V1	���-sVvn�nx��VF�l�Y;�5���x���]�V:_g}}�*Y�_���d����3�|)^�m�q$H��q�;Q��#'6v�2ęQ��z߅��bW]u5�2��z���@�Lp�}���Fb�0�����N���_������w�����v7ti�>y�4%	��]�7�zK����WD���|K]ĝ�ٵ[	#���`b�؝1��T�|�|N��0)T#�P����p~sߔX�ڢa�pv(���n@{�[�4�G7��Ԋ�_����?c8?�l�g}R+��k�u���4l�f�DMf�h:���
��B�R����5�e0g���� �Y�p��D|�6�yvte�E�
G�*+�����~�˕��o����v�C���6���Dp�Yu��r�]8x�hw4`��Q	c��F�WU��*�ʊ���aF͹���vlyw��=����iQ�ҍ����b�g�����[w����?5ҫ�=~Y��1�y~���⸖z�{��|@olj.s]��E��"�ő��զee�Ά�2�p��yz<�U�j��o n>�TB.��:M0x K���A"Q�
����@uM��JbסvQuRi�VU���^dzÝ�C�h|��i�6�׍QU�[�Л,ྵ��m�=��l�;(^; � ���F8�ŕ�_�Y3�"3������B�d3�G|��!�i�$�������g������ʖ�EX���(�8�؄87�ô!M���x8Hb��L��WMN��]q��ʕ������ĉE3ce���.A��H��3ӌA��nW.��uf��pD��\C��<����H���& :����r	9J���$D����B�I�H�}��~�Y#f�	=�=����p�
��M��bG�W�3�<�u���O?�D�C7������E�u 꺪�B�H�?5ҳ�_�i���(%Mg�-V�*FV�κ1	�5�]�_{��,itvvwh�Ν���.A*�Eo�߿
�Z� M�B��1��s�B8�Ò�a/[�����xu�F�s��1�K�|,�pι�a���^��5k��SQ៾�=vu�;oGG��&�|O�Pp0�����ï���<���k��И�h�y�~���!w�SBE���<~L���]x�w�v����?jP�#���*��)�b��r�4E�� �@q�ɘ�ֱj2��r*���X(�#�C���r^K�5	��ʊ 1�R���j��G_�|ݱX�����-������v���։w<�������@(�s�<K4�{V=��{wAwU� ��נetN�:�AxQ��|U
����{��p��_j����0�e��=�%Ҥ���]�`��}��O�}��Q$�k�YQ40�'��q-������V#�*`��{�����#���U��,j�YU]�`$���v����$6�����fEUQU�z��Z������j�լ#��Vt�TF��I�j��������=c&L���O=��+��[6���!DQt邋���"�j��ѿ��'�A�Pw=�(n��^ds%xQX^�{Z&P��c -d0��U�0�AXl3RKߦ����C�2�r���榊g�.��)u�Y���iģ1d�Ic�)]u�0��
�� ��94g����wj�3��{j�
�PԚ�1L�D����y83�:�8���f��V1eS�2>�G��,q�)�ɠJ��4u�A� �)⃝.���URC�mZ����|_|{Ӆ ��t;L���� %�4��%���`l�31ȳ�chM��k&h\�bY/g"������e+���I"��w��k�����A����Y#'�be=\��o���9�l��7ߣ��{B�V�L����b߅#G�����QSU��˗�q�Xq��x{�<�8�R�yQ�%��	�Pr�A�2Y�R�?��՟�4.8�~�x@~�<;B%֥�n4���+����[���M�2�?��ߢ�p�����j**��^z���V��������t�x~r�q�9Xg�}V�\J3KՏ�,G/�LL9��Խ>섊��X(���x��3���/^uL�<�����%��S��J��ryo0�Ulҭ�	�ff�l�x��Jf��(��Kڸl�2�+Ѝ1�D@J�������?�%JV6������#��FUߞH$z?�\��)w�_{��Ξ94X4�IM�~����x'�saLu5�O��Z�����NreMx\�3���%	_Z;����a��6@3F�����u�_�3�8�v���~�3�uv�*���h^�%d0@�Z���o�M�����z�}��i�9��98���
D~ 5��D"ر�}���ftvucڴi������3<���[��]K�V���A�Q��XR��--�v��Ȕ\x���}�$!���i'�B}]5�|e�l��o��Tw�ԍ���V����*�1��?��?�yl#�Ҹ�5�������G���<���`/�Her��/fR��LU.G[���1ԩ��*5JJ�$�+9���
�H�+#54�Ì{��5C!��niӜ�l���řa���Y�.�[	y�D��(��� �UK�A�	���e:^�Τ`n˚:�.'�u�V8f�b��
"���v.-�1�nͿ�E��|�غ �jTUj�~fN����C�z��n�k�ܩ�Xȫ 	Y��C���ۃ��J�W������]��d=��>������DW^q)FU�T�Sw�ƍ�1�e��"�5r���I�������v����t��2�qP;�:��sY��%���s�ۉ�BA��t����l~yW E&��!؝�&�^�����Ԓ8��yxx�j<��3��1�PD���ⲫ��Ɨ7	�j�yv�:¿���w��\����k8��LW�N��`��
i�***�v���Y#)n��Q������a���Ad'��I���-�����y�Q���'�rBSӮ�O>�`Y�<[�L	z<�@0X�ZV�*��V.�+���b�X�M�>�<�޽��u��E+�J}��3��Z�g�.�\���G=�?��Yl?q�RNVy,��/�c	�VnhZ6���T,��M!*oj���.}b,�����J�$�D� �B���V�g�l`����v<�����ʊR+e��x�#�؏��wFkk�|�k����&ݾz�m;w���BXr�B����;nE��E��FCES�1���<�e�C��B��A�:�VQV��fИ��7��}�r�z͛��Vkӄ믿'�|v�ދ��t���!M���-n�'	$b��!��6�÷��k476��Oc�wc���9��8g��X�h�(f�n_(���lݶ���SK�������k����Z6�Ndu�IŬ����v�̖�$K�_��N��]k����׍E���-S�1�*�J_��6�<���F����b��C(2�����?�L�<�I�v�Z�v�j�(Qz�&0pc0�ٳ%!����N��8L�e�����b3�b焭qU�ܞe�*%uǌ�X@�&6L�x����T�FMO��~#d9�x���}��,���S9ҿG%������,�"V��x���垔g    IDAT�
�z'&��}��K#�@��JE�)�>��;q �����w@iU��>{��O/��������b�-5����5�$�H,�nb�4*�b�X@�Bg���a�a�������y��G�����s�]�k�`������۞B���]RE��y�W.\>�W�vn��iJ�<��$~	�\��yNN��-�A6�D2�dM�����^R��z)tw��C��T�=>��Z�n��vД���S���5�ׯ�_|!v�L������"缜`��^��3������:΋�_:�6�˩ڥ��5��$�Y�Ι(��}�GcԨQ�۲u��*�[a��0�0u7x�a�!���Jv$tw�a8�����҄�[���a�[h��������"�J�kЯ��2�����桷�K�:�3Ύ������Ҧ���jdQ������ĉ�����(E%��b�hkE��K�q.��8&��3U�����;ef:��?��Q�m3t^	��>.����l��U�������m�uWg�0V����y2��̮D0��4�24�+�v�Ҧ�$���%�.�	k�@���i��`�i���뜅V@T�LC3�O�д��mY���c]k��k.�Kgvm�0�r�\.��i:Bb�&|,�ïi�ç�t�<���Y�4[��pm����K4��&�gzF���M#�P�ġ����Y+{�t��I�U<"�6sF���9{"���-"J�pp�qDҎ���OVdv���=�G"�{�**)))i��}·k�=����l<,�ḣ�Fee9y�a�)�aY�3Ę!1��RZ�F*.��h �hȇ��x�n�������93w�B������O���Y�H$�^�y��1��ЀY<�u[�"�7�	ѴFɰ���b��5�<W^r1���f����Ob��/HK��RGuN=�DT�W�As	���@sS�|�����\��x�u{�W�Q1X1�e�Ͳm�\��N�G�%������� �w@����v��5�p1]����pz0�؇P.!}ܘ�5�>�X��LjF��3n�����ځg�/�3���0ui�"1���yaEps��,���=�"�KOm�e�
J({l'sL�6u����%�L�R���&�~8㤃��iS�J&`���ր�n��17x-���R���7��lEyc%$�A��w����,�∞��	Z�m����E�[���6�rv	i9w8]�U8�v�Qos��Ə���" �(�?�uX�s3O��QQ�:i��'�S��p,U2����Y���}�Q����B��X��lؼ	o@u&^B����n� ���Z���X'$V�P�X��.{m-��I'���8�պ��Z%��G���RE�:��	����r翥�u{D��Qi���c̘18ᤓ��&��h�j,\�zҔ�l��v&�x�!- G�"�n��l�%1���q��	"+��6���Һ�~�%�|o��[����׀�/8F.�������c����}G֍m$r��,�뗊���P+��|0�M�&	�I���8Z�L4�ס�ez;;��ա �������񹴠����.�si�����VӴ[�����q:K��ϭ���SG���*W�u�ʟ\�F;&EѴ��v3Kp
��i	ZT:h.���2��k$ ,���0E��%5���tR~[����d��f!N�xڹU�a�[�fY���
��ʦdȧ��T:����"��k5��O=��!�����5����]�p��D��b�hZV�:hv��)d),b��]Vfuٴ2;ɑ;M�6<+xի��P#�	��v�d�F�	7BM�n������G***�|Ӏ���#�=��-�MG�TTb�ԩ�����O=�D�K*�~6h ��J%�R���$�'{;QH%p���<��Tz�n����`�^��/��PI� ���/�cƏAs�n��������^d5*n)�*�y,��0z� ��������ü��Jk<�u����9g�)Jn�
������r��Z477��w��ʕK���թ��p ���"�v�Ft��a��&��8&d�%�菋~y)�k�=��K?B��`��}`y#h��������FU�#�t_{��Q�(�s�[n�#�?
-�]x�ٹ�3�$�
|��iHAg>Ѹ6��g��l�wɺ�O��'�3��m�/��d,�D���-�!�B7�BAy���eB�dk����q����d�1���r���t�����l�Ma�׎0������W{{;֬Y#Aݮ �>��%sx;��9�T"�}6k�`$���dN���͖I�x>��%Sq	�S'O��~v�h
�����������9kW�B��Cy׉��k�I��H�G0����c9{w���X��g�硇����PL�dQ0�g2e�RR�F\:<���XC�Ǐ�;�L�J˱y�,�}�{�d��900q� ۾Va�"�<��Qb��D�M@�J�Xe��lI9M�S"�*� ˒�E��A8��cPʄ��k6n�K�.Ķ�f��k�5���D�#^C&��R(&��v{1j�PĸoZ�q�̼�W>߸��V�Sq�|^Kkg�ｽH@�<n�p B@����f7��*�Hd�2h3	U�zX<S�L��'�ܗ����E�)�Dw'v6ԣqg��x��M>�E�砤���˨�@y�l>�0��0Ѳ��b�ʄ
 �^
߰�PS_ ��G8���}��{[X'Ipl&��O�õ�"�'��ѕ�ja�(�3>��1Gw_k�!8�=/Y ��t���"���x?<t�o�N���7�S�M@O��շݞ��8�	讒�H���� � �tf��*]f�4��gs�E�p��#\�p6G.:�q�����/�Q��4
�ኃꗇ�����N�t�����K���k��<A�����຺���,YzӮ����EE�!#F!	bK�F�8 ��f��O'���@�s6�,u�s���P�e��I��轇����,��Rx��̙��2d���
�5jv45J@����&Le@�]�]Fc�µ���+�9�y�̟�����^N?�d��9�Jd��ʍ�b��TU�ټa� v��}���c��w_�#A��h9��3J� �W�Z�)L�
����H�?�կPZ�)X��3���E��
��r���*�r[��0Ni($]�]�[ehji�̙�cʤ�hj��3������"����H�2�\�¡�ɔ��hn�.����~��f%���J�Pn�lZP��D��{B���YQB��`8x`\p�y���Bg'��������0P+����>��T���P�� �Ug�&�kn<T=#0������R�%y�dS�͈ϋ%,�	��YPm�B^��ec�j�N=n�4	zs>��W֣'w,�8�I�򩌈��u�����-�3&�aQc��X�G�rҕ;��<�IN��Pk7l�]�=�-t�=]�ٲ)2k�e�"uR,8D=>��>}F�!A���������JB��B�Cږ�jw��8����,&/��i��O&��)�RbF8�'x�����Gtx�z�	iS�|�i(��',�@8�����>]��ޔ ��=� ��7�=A�#����%y��teq	��7F�X($����.��>���^��]I��P�-��A����~z6<���^~I��4��1h��;�@�U�ܟ�=:σ�6�f�>u�T��}�+<e$HĻ���;���)׃�9�pBe��L�B�y�$�я�-!A����^���S%�6Ŗ��_m����8].�F��ęS)eAIHm�c����c�+�]�3�;�t�����H���:���=5�sb/ğuk���\��O����&�wuun�t3R����u|ЊBpEB��;�,`�&��5���`��L�2J E��	դ��~��B��E�7�d��MZm��Ղ�,�쉘�K�J�)*-��p�d����*J�-�Ǔ��rnò����Q��r��K�t�h�IE�;{���\ii����*Q�_͓��qC��njZI+���eW:;Z����\*��m[�=q�X���*�H��ԑ�==����R*�*q���b؈��7�{�z�nF\g��]$����Cpݕ�c@Y� e�{�I�0�9x=n�M?��p��	��'�%�\�R.嗼f�:	 }�駂�6|�,Y�SO=E8�V?9�'X��475a���,�/� ���W\�Hq9�9+�X����0\��+��J����Q󣚊XL:�n̛�6�n�TR���L�v �ۻ����xf�K(h~���Ո'�R!��F��I��[I����W-9i/����|6%�o�`�?��{)-p��H0�X4"mP�
C� Ǝ���
�%���;%\����HeS���r6P~����i�:��ٝ�:+h~�SI9�y�L^3Y���Կ����M0�I%d7�];`92��z'B��{V�ٌ y�g�y~��|���ADJЩ5о�U*�P,*ɂ�pc�u�\V���@6��{���qD��{�	O ��_�ŝ��/���@�:!A�"����N^as ~K���c���i``�j	轝�ݸu۶���CF�HP�3i�
��*v�;ǾU]w��M���O^g�`,$k%�JP�|y��Я� ��d�3oP:��֬����
u��4����+�/lASg�`g�+�-9�LNJA�r��8��K$��Q�y>|.���_;w�E'Q����%���bޜ�����R�#�6j���K���^�N�Й ��I�e�QGɵqdp��D�����Q_�=�]��9��N����3Rb V�{���-S�>��=��Mry�aE�����}�ם�쟓ɞ*�{|�Dё�0�^P|K2?��(>*M<U�����S_��i�9�<�/��c{����t��#��7p�ߌ�g����z[[�iÚk����z!�v<p�B�Ƣp�ª�p���M	F�2R0��5�OI�!*4� md�y���y*��N�7-��!�}	��)�#��������(�a�a�2����,²,�e*��C��eOIR^�ggWo� ��P$6Y����p�HDd+������CMn��a.�g������hC2�#3]Vzu۶b�1�p��ɂ��4l�ۉ{y=����j���]�{�MM�1���ہ�N�dry]����:��.(`��!���W``e9
���!�B�s�p�9g�ܳ"�T?� ��%���:s��߿��m۶aٲeX�bF�!V����.��}�6�]��.�/�A*'�pv��ፅ����k�G���ك��})�To(�Pq��ˠS4ۋ�υ�̺sB�z~�|�n��ъ��p���`ځ�E��R�?�,���a�-t2	��&%��e!��9��l(v��U�u��K�7f�b`�fR�M���U ���)��L�-Ev���T�C1��������l(N{өȝ��ܔ����'��~~-���Z�Lj�Zg�)��W�rε����K!>o����00��l��AQ9��)���>\��}�iiɜ_��8���8�����"Gl7w���iI2���ݠ��������[�l؄{xuMͰ�~؞��|l�ӷ^�"%�<����D|��`~ȡpY	|L�֮]��u���	� ���Gu�B}�!a���g뜇�<��DbR!�Q��M��A��L&QZQ�	�M��I�#��".B{w/��=u�MHK$�އ�����B $�(�|zy3� .���U��;jk���w��ܬ�ؚ)��G��>�&�X�k�-D>��^ȡ8��W^.	��/�CcC��BP&�k��`��u�JY�/g���1��y��-�#�8���lH�L��۶[����MH�Ta%tJVߺ=�)h����s�.�׭���]���rӲ"ܒ��2��(ύ�)���k�I�FRQd��̂�h+�Q���Q弝�qM�voX����ENȲ4�n��?Km�L�-��!(�/��˙˺�1�F�����LK3��0�����M�Q��>~��t�"&�$n�S�x<��4m[���5��6iR����nm�׾��l{���| !ZQ�`I	�pHf��t^�E��Nu��p$c�H}(x���2��R	"!p��N��Hđ���Y����v+�j�nq��f�.�W�&�����j��`@��\Ф�$��t[G�Y0̀7��'V�̲	^#���h��Q��dE����3Y�ti�ɶ)6?�~�;��Iĳ>�b���
\�:{�{�X\u͕6|8�66��Y�`��z���{E��C�=
�p^o9�?���ү
f&�g�|���0�g��T�t�qp�榛��yd�E�r�9o�X��;w�a���Ǎ:ۼ�sp�`͚/�a������&��>������QYV��/�C�GK[V~���qTT� �JK^(f9�"�Zs��R<��|��|�Le*��p�UWb����d1g�x��9Х�ld����)�J���(Y�$��f�S*sN{���H�K��Zpʿ��4@�[k7���U6� �Fv�	i?;��÷v@q�N�vP�N�v��#z�*�T]�=��Q�r���MQ%�ZQM�oW��т��6:���2�ǊJ�y�Z�����*��j� 2/h�c�U@?묳�ڽ�`fΜ���)AJ�`�������RĊ�����]�TF>�6͍ϙ�&&O��[o�Y�/�o�]�>��uBCd�/�>�W2���#�jf�.>�>3���(��0�F��uDPc>��Ν��ݲA�k��4>>V�|�C������Z�1�UCuJAm+��d2%�C�1��s�߀	xeUUEcbm���	o���lCGOBU䚎4��4�;^�Е���N�d��Z����ǩ'���|�^})��ؼ~&o�G�˯�kw����Q%���Jqݕ���>w�shiޥ:%�r�L��d��t�QG��k��8����5��ѣG��0��j�nd*����$���q ŕ��(5K&L V>�;I�G�iKYI��~��]���\�R�0�LM�knWZ7��t3�r�!��b@d����偙�iB'��a.]�X:e�]Y未�g`64��HD-�U���mr� U��S���z.M�cZ�W�,��[^����4S���[]����B;���l�x��\�e�5���4���-]�
�����)���E�<��i�5)���ΓY���w|���H��8JE�R��c�]L��Q��7]��ek�++"��\ �A� r�i��A�5EʤR�����ġO��p����! ���Y���8�c�ˡ��¦%�'@����YK����T6/ �ްr��%:9y�tw�jA�$��
���SX�* ��C����ՓD^���g����ې���F���������:�u�=��ԂY4���H4")�8���_~9���|&�'y�����Y�1�y���H�I'���h��u�#�L���D�m�[[Ű�}�!B]Y���r�)شq=6�nŏO?o��6��=6lF���='�_]�K�؆���5���*��%e(.+U ���P�	�Ҋj<��l��b���T��n��&M@GG7{�,xm�:/\����G�A�;
M9@4�彳a��l�̟	�#���7u�)CJ#��pHd\I1�qr���q9;|o�;hmU�b^?Q	3r2Gf@T�?U�;�׃�׳m'��d�:�l~��w��
���2W�t҉"��v�2>���F��J(���ji�s��������e���C��`�F���&�!I �;�<�0Hϟ;O>��T�b"�*U*tVn�8��&�-LΛτбT��-M�2�9�&��WZ��V�������)�PҞh�bk8��r쎘� ޽�4�^e�%�<iF���%ݙt�ͻ����(�<��#��׆#=A������ad��g����`]B���`����INEh�`J���%x����p�pyarv*���X��
�J�RUb�N�
n�;e����K0���x�������L8) +-����흽�5k���$V��ƺki    IDAT�A!��SO>���-v��8�\�*!T��3fp��JJX11
";���9�~:3�qE���0u�)��n���p{�#½��b��S�E��0v�_'��;---���~���d�q��`�d�=�h�x�jkk�N;�4�&�/��������2?��ϟ�-)/�x,~zS�/��Db�r�ܩ�}>�3b���wwk	�ߘ4i����;��,�7��h����(�O,�C4D J�J@n4W�x!S���V� 3zn�lAx���Fa�H�L�L1D�$s7���%�b�*���:�p8*R�\������V5;:[�%��`�k7u>L+g�i�f�Ե<�5t�O��B݉d�^
g��ЙL��'"화���'<�|2e�E�R�1�	���
PT$��	�;�Ů�<����Í�x�pC�ÕW_%}�:�y�}�ڼ&y� j�;*9�YDH�)nk�]y������?| o�����p�Y?��M��Ŷr�7)*t|�8k�I���{K��شo��>����k$ƌ��^Y�����=��x�RL=`�$-�<,~�-��A���KQSS-�F&��sC �f��A��z���Jm;�W��^Ɗ/7HW�����G��C?���,�,d�(��M�䓎ǉ�����,�Q:hmm��ի��G(FSK�m���u���1h`�Ċ$�`�~��e�s$S�Z�HDsTe��	��^8U�C��U�ܿߨGOh1�"��42p����.�g[S��s�=U˘���<b�0Y/\�<.�f��S������2��q#�ҁ����	tg�n�4S�V�9��Q�Y���9�\	�D�ϟ3�?��|._�\���9д�����R��+�s���A[�n�fwL|�X���0v�h�}�_%�X�~f��0�ַ�Щ�ǖ;Uveg(1���\^݂���Y:GY�%�؇ �CEA.@����v4�ډ�����	��	��CaA�;ʓ?��(PC�
(lII��4:��("E1��B�l�р�?X��+>AO��`���!=V�uO��̈U+�(pZ�[7�Tɥ���p��b�����d|ǟ����lŊ�p�?��{�W�#���EE�y���4<��3ؾ}R��4G��7.�O��T$�ǒ{R��N�%פ��V��bj8�K%�2n�cKY^� ��W  ��53����aH�߯���çM������]�e��"��?�/W�;�W��z��Y�D��"��W�@�
��y���HQmDf��P�U*�3�ϋ4�z�1�^tf�HqH.?ò�I`��-RaWWWJ���aiq�-?�����˰^�'����B>gX���d4M��|�P X�y}I��N�������Ƴ�h:��o����k�I�ҥ��)�Zp����+���ʜII$Dy,��`%� ��� ��!ԓX$ �n�����!v�w�E��źMpB�.�M|�ޣp��cȰ��khĝ�ރ��M�{٭���b"^�������+~��������x�{��{�J׀��Yg��)S&���L����7���A6�4G0������Ak[^|�e|���(��d�ֲk�Tt����6m�EGO7F�5�&���g�v��44���m;���*���£����M�X���J�Ĝ���k+Яf .��
8@�C�����&.n�9����QbG�&��H��$���~�J����]�m�6x���%�J��"]�^4�!����ŋeM:U3AQ�9�+�P eG��b$���ȿН����P�\�W�kڑ^��u�/�E�Due)�;�XIH::;%a�ޥ8��ot��qsu�I'���}\�� �&��.46�BW<�O>	^x�����<��#�<MK��|
]�aܸ�1jo��J���*����Vn���(mtyO�o��&������w���ݴM�� ��������J��@"
�\Y
Ͱϩ�%ly4�}ǎ���#�+�>������CX
l��tL�Ȋ���X]��:BZ�<w�cr�y�t�olƊU���U_ Y�XPG�ֱ��Iׄ�"^�rfNa ��)}v�X��f!�?���8�Ѓ�M�ѺK���1�tO�<�Yُ>��=����+����?� bJsf?#,��}��?:?��1�	�r�݉\�}j{v�� *�-moUC�&�"I�Ig>?�K��!㸂��ՕU��=쐋o�䂥���o�
|g��X;�S���������@��*��mn�RBiDA��NXU�uG���pHq�@	�����(��@YU��T��,V}�
��<t
q��Voiii�K����O��v��Jh~oҫ{zM�0�:
>���x
���Y(T[�w�(��C�0�V���lon.�r��ɋ��wm����D&L��`����Rԝ�,��>��è**�j�2Ei8��[��h$$��H,��t[wucѻK�~�VQ��>�|<�\{5��m[q�=��ng3,z&ۚ�4�җ:��fa���7�����Cp�=��޻��[ ���G�C�.2�-�ͨ�Z'�0�I ����!?<�L��B[�R�M�"�@	OJ��V���W�k9�->��1�L�2E���>��c���"��^Ç�\��=�M��5���!D�*p���kd�1p�`\~��Կ��A���G�����1�)7�yu�~�Q�77�e�vq�"�_��G:!�����ͧ��]q�=n�C��5��$Ǘc0��k�/�;�T�ܠ�>p�c4���sg���7�j���I�d�c�p*z%����N���*.�H��N�?�Y�֓�t	l"]�`'��9JP`8O�I>f�{�[�D�N:g�u�t�-Z$	��i	��ǧ�.I�l�W���-uy����wuK"FJGG�z{���F���w��D�����-3��v�hsM,����9&O�\�QĈ�P&%����f���8���1z�Q2~���fL|��f%��Y
�V'^��P��!M�	�Ǉ`$���$�U��h�=�&�d�t������e���W����by���gG��>v>Thr=
�^���f���8`�>���I()�٦'
�����:�7�d�R���;p�J]�C��-	��۷#�I���r�'�*l��˨�/�8��a~}$�W����-`D?��H��\����b��+�����1��n��yߘs����>�;��U˪׼���`.RV��Q�F�����%Ȋ]fIv�ʇ �, f���
�3����(��@%�M- ��a۶�qSa�΍+������ҿ�J"_VVk��ھ쏾����]rWCc��hQ)~0y�<��zi�
�|//�a��A?jJK$���M���X!��H��زc'�\���:�t��

�/n*��\y͕0h ��m�̻�B}S����!
��]�]f��7~͕�.-A���x�A���"�p�9��i8�����SW�����֊�ݻ1a����e���KlݺUtTۙ��
b|�L��ٱ]�j�F�����l���6m�(�/B�s���c`8������{�ǧ�7�t�$`�����a.|��ǰd��Ȼ��z/���� �]�����ʋ"p�\^��X+AeU��� ����d$����fr��͒��>򯽶���� �����\�m-�?�+Ou�rw���{��v+�g^��3�r,��w��Sqc8��s��л:;���s�lk�vii�$Q�,�th&����_�e��i �bӖ�x�ɧQ[�MLR�>�8㬳侾��k��p��k�M�h�b̀b�O&%�PI��\��%���S�`���"D-���Jʊ�Y��3�qK,�W�dk'2�pkF�|2��P�� =�W�%P]:��!�G0f�0b�`�2���i1�!��IN٤�v4�M�]�P��C\�&zz"��{����iܵ��_�߈T�@F�ч,t��2F�EǜHo~�`t��.|g1�QI2'ڢF�J��aQ$ Y]ΨgO!�(H�i'b�)������;��z������/e����N�MQ�s��}b�j�������
~��q.�T�d�Pd�C�TPO �4m�G@�S�G����ACꎜ~�������������3�N:O�~���:��n�R�����b���C��HeR2g@���p��А" �뇷�H{[2���-������\6�����z$e�g��!8p�Y0��>�������Jj�}c�W��9����y���v��O��aڴ�$X��֛,�����6(LB���A�4*���ij�E�@�];w7�v[Z:���)~��vy��		�������� l�߁�n�M�ۑg'�(�lF�/��)&1y�x���ע4F��=p�p��}������/���H���M�dn�͚�?Q���mG�Th$�M� #5oS�*�����S����R�϶>�H�J��?���J˰�>�`��&H5��4�~a���!C�������0i���|�'���������P}8h�~ܯ�+���LIp�K��d���|���f�|ح���AU��3��U��觟�@mm�lxk׮�;�ߒ��qr�FC�5��U8g�k���:��s�T[�(����ug��l�{&<~��Pm
��1r���d|�w����W]�Oպrɸ�1��WS#U:�T�͟���!�+�H�4���=W���_ģ�>*��2�^z)2�<��[-*��c��A��xO�`Ex��m�Ub��� >]�����63o�E����F���;���T��38Ɍ ���`Q�����g�H�`@�8��X�O�נ	����#�c@���BI4" L�]�N�әn�ư�!
�<��czI�'�7��U_/��l�BW<%fEL�]���Kd�+�!� �Jث�|�j��-�v�B��}�D ''��2s:����Ҵ*�-ubw|l�r�_Q�Yw܎H ��_{Y���m��h�k���ۇt��[ۯ$S�8�{�4�Zs���5�[ �*&�	�"e�yH���~$H����)Ϯ�۔�6hp��xޭ�<��
�[���n�Z�ݴ�xK���[��Fp�ǤA3T���jV.Zo�Tb�Uz ���$g~����%�Y1qa;�?[^Y����u]���_:j�5����������䃇����GcE8蠃�޶��!Y>�Cl�+S�����~��p�/3�T>�L���z�.@W4'α)j"�	���W_-�i�w܉�������X�&��y(	��x�x�5(�2X.���˗,U<cR�tR���w�Q�޵�<Ҕ ����P� [��M����\Z���m�*�7�U�Y4���R�ũ2��}^E���'� �L:+ݦ��r������e��~����K�߾���ю'�~��ǹ�n�A��h #�����$���x�	��t&/k�1�)���@6��xw����n�رc��]�trye��f�NŬ�y���
���+��Ӫ�d�ϗ3�t*lg#�u����e÷�ڬ���/�N��lmo&�ހOT��\?�3���S��˵����g����{�����%KQ��Q�;+���;N(�<����㩧��4�ᨑ#qÍ7b�ز�5���豣����\��	$9?��?�0V|�J�#�8���FD�c�Z߄?��l�k �zt��gUb�����L�h�� 	�5QL3�U�iH���K�qV�4�2��z�HEᐤ�?ҫ��S�ƀw�[�A:Z;;д�Y@�������Ѡ��U~���ǅ��S�ױ�U`@%ZD��AD�t�ĕ���m+��/X	�Y	� _A$�	�#.FP9��`v���?�4Ë/�~8��2������ѷFU�Uk���:��3��?U�
W��w�Ǐ�?(�����;�G��F� hA�](t��8���iSΞ�s>�6���?�N��_\kժ����O�in�,����/+unZJ��"���8�aΑI[�Q���A�T-��:�H��(K��,M�������=޷"E�wk���/W������Ec�\���]=��B�"�\�;;��+/
G�؈Hn* �p�O��b)�&v�Os��?�L�\[�<d�P���nE~�T;_|��B�h��_���(�
�l^�J�8{����CTh;	������;}��)��m@@MR!��+�8r6%�NIX��������a�Fu��Y���,%Y����T\͔�	[�D�I��0n��P@P�i:�y��M�x�#����LFuy��՞�=s_y�&g�.д�(w"���"�y���$՜Y���9A�2A�1�3��C�W�SC�Vc�v�	(++-{�сA#�5����E��v��p�?N��?����8��":T&ӗ�x��������t��U�-�!�[�V�B�r��^31������g2̯��&I��.�!e��O:�\x�r\/̛#���ơ�����w�-��W`����'b��jd8]�k>���YKK+:�z��3�c��M�*��i�0�?"cS]#�8c�oێ����.�P24He�O�[᤺�< d��̒bA3ho۫ĥLd��c�}�))��h�PX:[5��DE��;ԝ -�
�̹��������6�V��cm(``{g���c�b	�d�2ߦ�`�l$��噠�ν����)ZL��nQ�-o��D���Q!���$&��O*��pӍ��^C���/��*j�#�y����Hg��C��(�N����0
���?�aW{:SY>R�������"&�9��?tڔsf^���ی��y�����H]�΃���EF*��V0�C� y{2��beEI��d�T�"���2����(�Hy773�F��a��P�K�4����ť�蚊�c�c���yk��/��\gw��h��s<�:��բ�T��e�p|ʇ���{�4��!�C2Y
~�K�b�J�AX̠�j�ץ��J�\|�06l܄;�v�辧i<B�)��0�憐��,`���?�	�a?:�{]�v���\�zU�V��������ц�ݭ0�҉���i�Be�u[֬_�~��*Pe�bta�1h� r�4TV������f&ϟ!�(RT,�G!��3�
���Ѥ�Н��A*���HYIHf�m�����7�BJ���	o�ʥE�#�ѐ��P���CNP�}�b���"ҡ`F��L<)Ւ�OV)��;i�D���.^�vi��WV5��u6j���I:Վt/l�jG��9�v���$���?+�E��]��g���ٌy^*�P�)�W�dR#�J�t0�+e���L�:� Q�e8�s��/�gh����'�d�����˯�����m�*��?�я0p�x��X���F�y��Y�˖�Eo����n���I�샛��Vjm}#�t���P�	����(wb5Ri�ް՟7�ho�.�u�9�4��#�	X��UR�\��/74S�b�b"�C��hVx=H�3�N5�s�th�[�X��zn�$o��C%?䞳ÒW-mI�u�$����3�2�t�7��募��2��Fmw��y_��'֠
�!�q&��سY1��Ӑ1�bP,|u��ٍ���+0a�X,~{���2g'�]�-lʥ8�Q$ɖ,���Ka����k��Y��I�5,�'#��@]�v$Ӥ�v!�B��G0"���,���a�8r��so�>�k1J�ͷ�i���@�����:��S����іaVQĤg-�BAY��C��ۏ��	U+A���c�3��{�u�{��k�5��#�?�����1���8������y�f���q�w�	'c@E9�șא��'����!R5H���ݐr4��e\@ꞃ�w QX
�"�q�f%hP�'�}��~�]qQ^"�S*�|^���o?�gn����*G*��^��)�	�n�T�� ����R���� �)ө�r�o��� b����tfϝ+�����(C�V����$����F<��wJ�DjR� &�) �,GJ�R��0U������E�]Vh!�W2��������r��C�7�+�tCf陞n��M�J�5�)��L9�x��@4���=G��͏z�?F��h4�OV�Tջ��dYG�U�Q;9R��w9V    IDAT[�N��|����e$�V "g��ϝ`���9��?���S��e�$�)FD*��v4��nX��]���(Ԣ�gV�"*b���L�U��$v��g�.�u��������Fj���0����D���Ɓ��3ޡ�z4���e+���a�V�~�&��?^q���jw���3����F1�!>F���T<�~���q�����6ږf2b�����F�ګ��/	"�RY*���t	����z��5y3ɔ��S;a��2of�H���8�a ��8tA�:x��b++��@;w���	N��R0!?�_{���4���h##
V��WmV۔7e�,�@�!�9���݀��!��[�+i:l���ڲ	�W����?�`�x�Qi�;�LDyoED�O�S�`R�|�\�N@���S/�8#�텥K��~�N�i�Mp )\g�X�.�>�a��!��5}�y3/����������j}�_&��/��M��k��P��-+����>�O79|r{,
�5��+דN't���`b�'�Ye���vG�~�رc���w�z~Ŋ�G��7�7�=���?:�P${���avK��3���n	�n�E��F47�k~��rii�;��\F�>E��HV
u�>]�{�i��`�b$��s�"F�_\�34>�[�7�]�:)���P6�^�p�HeҢrǪ�t@�Y�!+_��U��윹h��}�ə�+�s���ƍ�e��T�ש��V>h��fG��	���I�����B��h4�񅔁�aJ�5�����xT!�}ai���V#���+Qd�׃�iv2
t#W�3�<?,3�W���` �L��#4�5;f���.y�}	,<V���8	�c��i���+_������i_:6QM��;�&Q|	�7�)�78,�U�Npw�3j����v%�=��F�"X�ʙ�/&"}�e�Uѵ�t����I'����?_�U^z�<���e}8�KS� R�O�)X�*]t�9>���H�#dٲ���yH����I�r�0fn��j�E�q��4c&�5�G�/�ݧ��)N?�d\t�y().B*���hQ�=���C>�o��e�A� �,]�~H@|��rW����������G#�����
�����e�5>����_�J����^I�܈�x��'`w뭷b��!ؽ�U,l)��s�g_`�]��eᘗdi���2R�왎JsQ�P:g�T�LpH��$���i��& �A�+~�+L�w<6����f��X����b�ҍ��ջ��pp"����}������l��J�ˠ��g�}�Ɲ�DL'^��r���Q��;�1�'P��P��eݑӧ���\���[�Y�-}���Y����*��\�2��B�Pd���uh���<V^3��e
��]���gz���ݷ���о�����UՏ�e^c[�4΁G�Ԡ,�'��n�|��8��)eI�>7<:����:i?�]$ܘ��7�ٌ])20xt��p&���Z�w՜�f
�JW^��2����A�0a�(���lL���A��)�n�B��'�!�<�Π��lJ@�4�����k���=�B��Ri�
"&�@4rh��CX�`���#ʹ��&*"��v���v0{�߳�A�
�2����j�DC�n$҆8�I�^����^X}gRqIX�R3z"����Ӥ|+Ĕޥ�mO�n��	i������L;p�(�-z�M�Jƺ<Ν�r��f��g�p*wg3t6A�؁���8��k������T�N{��P�*��}�>A�l��g���ܪ�.��-��n��� %�,2�:U�r��H�=V�r�lg�y.8�g�eNS��~/evC���у�(���jt�a�ҙ�$����09 �|������U��>cF���]+3��;q����"���r�yA�ϼ�V��v���d�x�y���W�G�x�|�B�����y��k���Ï�9������AC$i:cQ���Y�|�����uKI� mp�9i-Ϻ�nTT��G����-ҝ:��31�����c�(.��"����!�#�3?��"ttw�Ιwb��+E?�`>���JT� ����q��)�,��<�(��t�(���h���`�&����	l�v H!��I�!�L�%���ו�x��{����("ZJ��1a���d��74�f=��o &�)}k'��'�Dܿ����{��~�M��������˲�wc}���fI� 0��ԴCU��oz=�����^}y^}[�Al[��.x��p���9f��z%K'%O��]:��0�L�&����n݂����K?xҡ�&�U2`��l�4.f粑��Hg���<��D�3�O&zEq��z��1�3�/�ғ�)�C"���m)z��ED��`��~^����>yP�`D���&z���(�]]B�#���>���A��@![�����n+��~����c"aӲ�IH�)
[nēd��&І6
l�Ԃ3E~��t��0nX�H�F��J[���X�T�k*�s{
��$*�	-8���)�蓕��n��Wmj�t�{˖�Z�N�b�gx\�,����Н��zn����Þ�cg�)ɀ�v5E���I�1�)�����J��<���x_����ű�[p��u \@��u������z��[��:|�>�BA�D����m	D�D��H�-%IEI��H��
J�
}���q�f��1�1|(n��*�mܶw�G�T*!r�d����"o����i'��V4l�!6��ӟ0��Ixv�|���JT*�7���j�a ߺmn��v����8����\�˟�SN���?��s�J�ˀ
�:���ˤ$�S~���@Ss;������ �X�������ŗ^F:����)���ɧ�A�`���?~�QyNn���yK�<�lY�w0�`7��M�YdEQ2�N��8��`5*�ql"�?)vAR�C�U��R4���^��{��'-ǒw���Q�U�z��z�=��S���~��0@�*l�G����jp�SRQ)4H�-����"�p�V�]��0�%�v��	(��!5��5}�9��o7�������}{�����ym�܎�9��bW.	3�#�-�O��ɽQ
�K*t��=�t�q8���}�Y,\�y���4�����+�P���:A.�Gٲ���T����4��Y5e�qA���N��!�P��\9@(S��8��VD,���[H��Ec��Yt�3-tg��oi�'k7�WT�iz9KW��|]CI8�N�������_���1[�ܐ8D[�� Ќ*t�K�T�T���T:+�\�?^�Ξ� �8�2Y�$�<����+���X�n�݌���d�˙qIq1��(���M'���F1�K�������k�z�'}mo��<l�3�vf�N��17��q���:펷97QY���t ���{V�}���<��2�����lΤ��-�&��1����WjT֪��FOw/��2�!�,��g�!���7���x��e���v�!(.뇱�N���4Zd��c
����궣;��ۋ�ŦM��h�>���*�Y�in��.l!m.��������a�-���e.���eD��1c��w�$���;��;$`�E��#;\*��&N����0�wc�fds�6 �R=3�6N:�x���G�y�0u�����u&�D�hwۭ@SS+n���ev�O�D���S���7ޖ�~�Ǌ�ܹ�/���ǟ�5|�m����I֖ -C��� ��y�bG�5*i�����u��Z��"�?_�-�*1ϥad�(7��+?\�-7`���	`�n���?*�ɺ������w^C��=R=�κs�3��9c�����.dhl��#7r.�$tГ��Ї���?t��?����}{�����}@�7���Wm�~d�sZR��B��$�T/��ψ���톟մ[��Ϊ.�ģ���G#ʜ�^��o�!������q�89?��4�U� Nt(Q�?q�-G��1ӷLi!��(�EE2r���1q�x�5�S�YVM4u'Òv�$:�׆Tu"�A�LNZ����v����_���<���e,��t�·Lq�A������g4���Tچ_�	�-��W�����?�@�A/�o����{u�"Jf@�����/����0j��w�xq�����1w�<���꣩�A6��zz�PR\��#�]<ދ���&�^&<˗)Q�Rq�3���{���>Ip�����d,��᝹���s�e�����g���\O剠�4|7f�M�;E���N��������{��ӧհ����x�w���U����,Q��]��-<�ģ"JD�DiIN=�4�&��K��'#���Y J<�LH۟:�ւ��\�6>Z��`���K.�(����mR�{�	Z<R��:����P����$z{�;��n�GM�SϾ*:���n8��J�)�6�e�V�:�v4�j��!'��\��q�qG�G̙g��:$2'Vk��e�>ukp�/~.	�_�|֭['���t?�@|�|�$���/{�1���Kr��1k���u'֭۠F6>5a���V�G��JPO8�h�蘣�r�����s\A�Ao-~��[*�
]t��ܸ��kQSQ���/C��ZlX��E�Ǣ2`'���\�,B�h:�^C��Q؛�����p�X��"
&tbjĽ��x�b$L �ya\�Q�5Xܿ�΃����.���s��m���>���oy쳆~����-���ܤ�tR�y��C*���.kn�R`����]	�GG��<V�ܗ����âP7�2e�.U�T�jsv�@��n�j�(j�3��fB]Z`�1cp���bP�����S�R��8��Ǌ|&;�B�mIC�J���,�xu�մYN��?���q7R��3I(�!g@�1{����s�M� O�X�|�00�ꕈl���I/�}M��gh�A�M�_GCsf�yV�%����)=�/�1�����/0d@��'��H�H.07�-[����x�di�lH����^~�%twӴ�������U����:���C`��ȫV��.w�Н���;�|��۩��R�z˝AO�gqi��<�K˔k�=�a�D�����Cgg�h�s-]r�%(/)� H4���ťX�n=��aa00!8��q޹�H�����g�Ą}ơ~{�UW�왂,����uR3EH��	b0��e D�������+d�4i�$\{�5����7��glڱ9i�H�����{��3�j�Ǹ����%�H{��{�Iº���lI�؅�-������o[Gn����;d�cM=ng�|"~yṘu�C�۱cƍU3i[�W<�=.l۶�D/n��F�ji¬;�B��FaI�y�8������oH�}�QGI@e�kr����w	��������6��{}~��Fo�ޤ�:G7�&����a�+W|��vI���v'�7~"��7�^��^z	�[�؅�?��:�9.}�7���W�(�u^�O����l�Cv�A#�c����8�\����{^�pmcǆ#.��g��-Bܰ�k���=�l�{9L�U�L���]��7��-����W����o\$'�?�����i�gS�%�`d��r��� �%��l.)H��H�vN9�GH�2xf�<���"l�+[]	�+��:[�l
m�lV��Ga�@�7L�������d���X�Dv���]6�,����B���fTx��,��bW���l���+W��K��&��:zz��%x���ȡCe�PU^���{�(+�t}��:9t�M�$� � ��*`�aĜ��3:�8FF�QF�9�QI""9HΝ�9}r�o�wW�}�ݻV�{��8ki�O�ڵ����7N�ET��烬����NfR���&%%�A��t#g���	�W˭;�����a�ƍ�&�9ɓ$�\*�i'M��o�	��F�؂:���X�����M����
�}yH�sp:TB���*�WG[�l�?|�������LU���j�[����'-o�M���ժЕ
��WZ���,�Z�V@��@����R\vɥ1|8� ��	��:���v� �@�y �����'`HV��^7U�$|��1�b�O��~���Z{�w���a�a��~������Ȉ�뇝"� <��\nV��q��-�n���n�)#���G����ʪ~�ki�]��{����S�JR�C��N�������p86�馿��3Nƛo�'{\��T��g�����9sB�(�e�>�`� ���@�ǇsN���^{!�9�	�_�@�Wԡ�v�Ka8�i_Jz��/���۷��9����Qf��_}-�_r^}�u	�_|>^}�-���k�䰻5���$��z��2���NЫn{S��}sS�%��o�=7\u���>��}��4#�	n!��c���������ԌY�f���Q�p���=�|��W�i�ؾm�

��wt�.��x��FY�k]Y�Vaz�x��uX���o|߼�e��d��G�X�)j�6�G04����U����1#G��ʽ���[����p��>�$���֊�?����P�DjM�(b]�0R1qH�hv��Rb5J�j�(���	&��3ϖ��o���/F���a�����S�����i���<�4+�ʥ2҆s�2"(�j�@�������,�1��o��9��2si�ї�/I�p�&x��ie_+�h6'[�:g�-�2e�P�ަ-�~�n��y��M�x����h����&���^�H�._h9]@}��p�r�pb�������QX���}�����X��gq��&R(��#G���l�E���s�X�K�Ȉ�g"bw8%�Q&��9����j9�.K$���b%��#���4)k�B&lJ�]�ڤM�z�*t>�U}[ �Fd�J���+!��,s^wk��Z������wÆ�K/����::��� �nw"�	8#P��fv&�j��Ȫg{:M���C(�uG%�o.B"��c��믑�1��/���9t8Z�3
J@g=��c%����- �±8��B������w�n���ŕ�\����`�]x�����@���e��v����*�J����	�S�����ko}���v �RA�`���p�o.��t�C����N�[%�{}����q�9���s��w�)�:戙�h�s�Ϥ�R�5�x�	�s��y���&�{=�~�E�=x饗d]�s@p����W�]zŕ�
v��އ��V5^�#C:�dn�t#��K.ƹ���7^~_�%b�̡(D�qAM�@�~�]�'�r�77��C"��7���=���0::�dF����ڮ$�ͮ���֔�J�֠5O���ޠM1k����c�(O'%��D�Б��!�����f��ڡi�_Y�>��7�t߭�q�X����އ��C�k�=���onk�>)���̥�u!	 	�A	U�.68�$@˦I�΀~�E�!��_ķK� ��Q1� HLe��V*�t��fec�윳:��\6��g�N�U2&�-�O9C>}��叿�N�xL��Y8�&m�._��Uѩ֩s� E��H)��E�bk_Lgrtq6������%�����A(���#��h�[Q�R�|��2�8���E�*n��N+]��Lo(�I0���v��_?̘q��K����|���z5lT������8�Q�s�i�v�DDm��M)WV�|�<��H��B����~5��{�n��lomV�f��̙#��|pӲDW�� �B�������W���	Z����cal��zXr�VKު��6��'S�����	H���KQ�ϗvi{[�s���}�����$�ae{�Q�1@��[ I����m�����D3�K*�,@�m[7#����|Q�0$́ѣG�.ej�3����عGf�L�t�����;w��p!Opo��!ؽ��X�Nc�I�te��dA�yg����:S0"�se dg �H�g�L�e�/^}*��':���W���ǞDw<�h*"��9�gL;g�y^~�̛���;�%��(�b2?�����/Di�_p	�1���������^�ܗ    IDATw��E|��^v�l�ܭ;��F8\l\�[I��0z�G;�p������.���_��O>@S]=\B�����O8�\{=�����Y��9:��|3�L��7_}M�����w&���Jjb=���wﱑ����[�P+r�n�*��)l�x��Ƃݍ�]�М��B:M��U71|�5/����}܂�և3�?���$���F�����7�R��H2�x����n8�64Qk��X�:�����N�{��8�䓥��ڻ��ӯ���� !��j��Jι1�Թ��U#��V+�������XRi��؍\��S���[��[sE�홧��g�}/-��&%���!FJ��# 3V�v��gx�����8��Y�0H*٦�i�f2
�Š��$x���6%�o���9�o:�$p�W�����e�N(\ �Tl�>7��Æ�{�EEu��B���X�i3bi�R��αC*ڍ��b{�h����Kgp�kSP%�6t4.���U+EO&M��ÇJ���'IE�J~�����e=R��w�L���s�Q�5s�Z��1�l���;�^LE9K�j_Z%ׂ��V��ԥm�R���퇚�*%�cr�[�ڤz&қ�g���ɠ���|�>�ʫQ;p��`�]� _|��$mtO�r?����[��!#�K��N`�^�� |~/�x�i΃�T^A��؍}�2?�+*Aye6o��V&'cv�HC�\ęU�l��?�T��()��Iq�2�k�ZwoC=��f���8�L�py^�<7�[���[�Z�� �ҕ"K��񣼤cǎúuk�/�� &�"֓T�.��I�L�Q���C�����������Ԅe�W(9Z]�nи1cQV^"k�C�e4���6c��hm��_(�X��5�B�h&-|�Q�?\-J|�y�Z4�C~a>��A����GK2������g_���Q�Zo��fL;�|���hkj��=��������(L
���HQ笊�R��(����Q�I��N�w,V���@)e�i�	
�Y���?I����?�����������?�g`@��I�
�>���O>{�%�8.��!�B2Ў\��t
*#1���ȕR��G�q�)���9C��w��������n��g"�%*s�&��e;�;���,4��ۖÙS���?�=QW���CX�lT��6{<.矬��N���%��׉<�D*�I��%Z�7uUu�
�n��e�)*,�p,*�jͮ!���tР���H	z:%N^��$h{ҩ�XF&�QL�/�Q7%��r��6���f��_1v�u�Ė��щv�z:���P�x��U``�jI*Xe�R�y'�*�NK��ܘ���u؁��Z,Ɗ+��:t�T�˖��_60V�ܔ<�{X�_���
�<WJ�L�Yhvv`�-�j�[`H+�[�$|&(΢1��1 �w9"�	p�����wP�]�����0
�.D���?_,>�A4��K��׊��|oR���'M9���@"�����nI���Я��4�!ۅ�0+�n�S굠����EML �2��x&+�E��rB�!sI�N�i2�f"QNԾ�K����!��'�6:ߓ�������3��|�'��D*g�c!MXb�,ƍ��;w"�(�$�2�$v�� ;n���tJD�<�"-o��8EJ[�e���T�K�k�3O;�i
Iq�fI��2�b@����~�p�{�)(��"g���Z�vZ���f��x��O��܊d<&�0�w�q;�;o����E��=�ţ�]�ho�sf�G��p���N�;#����8KJġ�{�Lx�Z��ǁ��P4{�R�n?2�0;>"a��0���cƎ�Ã����>n�������p�xȫ��~O}��;�iǱč���jE���T^
w(%3�,R�\6E~���.8�t�'���'x�ӏ�Ѹ����
��o�j�~(s3�S#����$���J$2���5�$��O�K@�x�'��O?	�����="V�V"+՚�C0���d�ݸa�CQ����Z,���¤4u�<��@w h���Ê����-�A�
��`��ަ�_C�2��������G�?� ����Pڸu�����ܢz���ѯ����b�#���-�DҕA�M�����KH )?܄���6u>�S�4���ԑN%�UJIJnfl�9�@�b�2�7�5�Vx�޶iq����/���g�b�@n�ݺֽg㿮Э�n��U���xT�C�6�Pt/�8b�̕��RU34;��Mq�afɊM4��!+z����f2I[N���NtG�@�:�,�K�f����W_�CSK⩬T�eU5�8D�j�Ȥ���;���0���	F#�����<$"1�qM�<�ƍE���$��Փ$�|�����H�	[��BaA����kk%P�"W�i'M��C��4�i'Al�dR����N�J���~b�jΔy�`�G\� b�4�a�ݼ����X2��FD������Q-[:�B���K��¹3�p0f�A�!
c�}��s��E�����pҤIx�7�v�J�~�C
�y�۷��7����@Z@8����FT�ĝ�x>�5 BW6���QAm�LB�n
�
�:��9�HR�\t�@d�৺�l��F�4b��Uӎ>Z!��?��g`@��)|�-R�ܻ_�Ӕ�&��@&F��F�](ln/
��ͤ����HF���$ߏ)��N?�P�}�	>��d���ܼ��m�7XWČ�Vl7]HU`�a����f@Ϥ���q�d��׊v<iO<�$���{��JJ�1��cQU^��&~ieJ**Ek}߾:�Z�^8���Co�h�?� \u���YQ�����f�l��<�b���5H�U���|��[� ��%e���?�}��E��C&�C����_{�� a��q��w������1�_������3�����G� ��;�;���Tr����2�(CU�!͆<�8��>��C\�d��dDΒ�}_Kc�e*������y�5_ע���������=k������&�x>��U�[��`�4�)9��}(��&U��crE���(G�T\i��Š�'�.��&e~��F�{d%d�T�k���d���E�9&KT9���k0o�<��Q��|	��Sx�Ï�p���磰��ͭB�d�EcBe@����H����m!�k��`���P�G9w��.T�� ϫ#L����Ģ�PSL	�Y��gO�9�J�����U��	eO���L��J68��g������$}l�1$��!Q��KM�ޟ	&����cq�\� �?�[�`P݆(a~ފG}�w�F��A(J�x�C��;�x]���iǤ�A�~���A�啀݁�6lĻ�/](��3���kp�y��g��O?,��|��{w�@,��(-��Չ���Ny���S���Q�p�Ǌ^����W�����c���A�&dv�ਸ਼gw�Ќ8NHg�^�9&�ኲ��tO뺳d���9��]K�Ό�ш^�ٲ�l֦�l�]��z&����0���r�\ΰ�9]��9�-'?��6[JӴ���i{ƞ�:2�\�e���rV�e�%����dr��s����TLfs�����z�4l6���Q٥��� �p�\�0����%���i��%m)ݞqس��۳�lְk��g�
��k�tFG�T�t�x���\l@�c@�(*������ٓ��6mM�"]��R�Q<�Uo2!#*�_y.��ܧ�u�;�x��w��Ws�aF͠�Vh�� ���_~im��/�g�j(�{.����&���]'nL4>yꩧ��A���]x.

<�,-BYy9
Jʩ�&sm"`7�ۈ������E��?�lZI�z]��C*��rV->��MO���D�.��b��|��ױr�j�V����vN�:��>l�y��>g�L��m��+��ȑ#q�]w����a̘��/Z"�9)�hoJ$6�Y�3�L&ϏjG��S�k��쬔��7~���f��a�6)x��c�J��U�+�n�&mʹ�d��k��um���{F��{	�浴��_5=lJ��:�[Ǒ) `;���O>��y���W,�.U�˴�̤T��5�X������*�:�	\���Rb�$##�Vs��z��)H��8�_e�����6|��W�9=��WX�}4`�x�b�RZ2���!��-M�2�9))��@+�#�8��v�  ƌI_t���5� �Jl�Sj���G�5����+V��ھ�Iz�c�f�B���'OÌ��$��<�\*i7�i6��=+;]�"��T�Jƈm�����ȈϺ//Ox�-��9�,^���N*Y:*x�69�6-�������	��y�,-\��4��/œ�>-��<?�X_t���<�ԓX�r������
J��h4,]~^�<���A"��Nr�P����S�L��i����:��@���H��$p��vg�Ԅ?�~`RD�����9;�"
ih����!��1���h 2@�*�L��fP��[��в��4�z��\�٧DT״��г�8���f��0%<�
���iԏֵ�-��Nt-�BES��$σf�6C���c�t]K�9�d��C֡i����	����s�d*�kZR��v�cQIa٧�ƌ��ǰ���?����}0
�|��k{��ӭ�jn�	�o��~�]A�RY1� ��E��%�2�v*�ۂx󭷱h�2�Hcu���+@S�[=ԥ���T8��!:r�� W6	���i����h�x/<�<�Ν+weE)���2�\T[���R�&Xͦ����ѡx�۷�D$Ƨ_|�ŋ�P�X�ћ�� R�������Ya3(��;m�4\v�U��������E�ɚ�)�����������߰��?%��}7x�³-�(A]s �?0?,_	����ō���%kM�y"��B�����јTՌz���|�n��MG$���'���W0G�ԅ�L� 9�YЭ��%
c!�-nz�klm�V%ϟ�v<��F��
���.��h�)���zl�s����3]'g�l��F�gV����2 ٮX��7�֨��M����%��!�D���"�]%4��_#�Q�	� �X��Ob���d������E�]�T=5b�8����^����6��~��h�~�H�w�?p�%$ �n_��޹�8�U,9s�jy��p�,Z��6l܄���@���3(��M��c��
�r�T;h���9S��E�c�I�&�X38c7#�	^Α݆@G+J
��!�;�C �̇ł���Y�����"����p�x�vӟP��G��[�垝{D!�H�[T��� 6o�!�~v�hfs�y�J����a���"�D��t:�[E鏟Q��l
'a�I�#p��E��3���U���LDq�q���֌֦FD:;��!�dm�	�8� ��A=)�p�I�eg+c�r׽�bSdʲ����_��?����3��fo������}�馕l[	��vz����]o&@ﱛ��L`l��`�k�9c�nl��pn���7s�qǿ��5��������`�u��)��"�j��-�W7D[:�4U�Xyg��$��~�8b�(�_�d)�[[��g�J�۔�t��nv��c-h�$gJ2r6�Ѥ�p)I,�8�X�t�U�e�x$��^xI�ۣ���_s9�W���_� ��l�r����k�BWF������{X�z����R�,:���]]]_�{�����yy�w圝���?ߌ�G�Ǧ-��t�
#Q���;:QQ���U���E�y=�qr��|�)Q�br<x�����QTR���v�s�X�a�ۚ�ƤY3�{5�]<�ܬ��*I<�e�����.;�dr� �$������c�#�a�U�u��=DX�J&]��p>,�XS�j���SZ7�5���w��Y�%�������pX}������	�b��t��8�9M9(=ʀ/� 
�������H!g��0�Q�>�,��� �w7�҂b_�D�-\*�)��.��X۷nC��C����'c�����oVg��2i�s�M��r`�A��+��@X��)R��cp%4��v�5WȽD�;�阋�_.(sv`x��#8�X&�4Xa�O���dR����!x���ڵR~�U:1b3*��r;�#��z�Lj�����%��"%�M�����cp�o��tES�9{��fhOO,ߧtG�uAUeŘ���{�H,[�XDl�M9	˖.ſf=,�IIbQ�2'�����mǕ�_�I��ￋ�?��:+�E��{�v����e�Y�\���6�80@�<'LD��`��Z�V���A�L���z;�ˡdbr�����w	qlC���&4Zi)
�RdϴQ0+��̶�u� ��}�kԺ�z��,��_����ֱ==t��Za�±�:���a�;u�y����{�;�$��#�&�_�z�������#�;�U�/�zO�[�P�3���!bL��p A��=p��0�x�N��-`v�تd�0	ɠy��4����"�!�L�؟ʂ`�05��=�3;��d���^�`���*��w gM>7�p���X���=.��2\}��8x�A�ׯJ*ZjMS��-'-S���\�RZ{Ͽ�v��-3�c�9F��wl�%����DW�E%Ţ�EyɃ���\�)�N���{�n�z��uH�!�����P^�W<{r��^�=yx��װj�Z���eϞ�(���b�z׽3�f���������*��y��+7Ij�Q��M,CI�����/�ǥ�9(	(b��"6����'
7x��KT+_9�H2�k�kɒ����Zv�2��_+o�w�:ۘ|X(w�
��0XZ 3'q13g��k���1�nW����<^���َ�mBCc@g���!\��\B0����-)*��(���:
�]}� �_}��Z���b�+4�HX��]:�tu�#����~�N9��K��oA1<y(� :�f<y��⚫qԄ	X��R|�����T˝]�HX�RN�t���Z�a�W_���ު5��&��9
��0[�V�����0-uUg���1T��k�)3޳D�_�k��ߊ��5�O�E���/u��(G����Dzv�K&"8e�<���;k�J�'������$C�=��y��3O`pM?|��X�f-�rӟ��o��=�|:
]dV��@D>�~n��ZL<�h,��|�p�r_�{Q��a����6�۸�����FP��J ������{�,4���0t�5�q�t�4�"�#-|�gv���t����$i:G��ϿM=��AEI)X���-��*l���`�_�r5v��tɮQ�t�T]=&��7��b����7�)��bs���l�S��:t~T�����yg�2�L�;���5�6�s�k�����^Q]}���S�0�}�N��?�����|���6Ƶ�3��cq���hk&�vd^��)F��cT�eyR�TA�֯݁TNe���%�X	>���̗�y�tTU��3EEri:����3��υ���@��X�`Q�P]���C���R$�	�u�*X����UӰy�V�|^~�e��	n�8y��<xȁ��ƿf�JQ�z�w�9v�XέJ��'L���{�b����DB���JG6��|�D	���;S��e>��K,\���n(�f�e�hl��=3fb����<>iw��ޥgz.�Q#�������*U�wu����w�??_6���&y����f��MY�pQ�����Gv�P�֬Z�6��6I �w�����fUnbB{2�2����m�w- �U�+�B���a�E�
�|]>�.��7SY.�֯�&A-���͓J�:��o�������z ZVdn9v�̴3�-	B,ǹ瞃���[Ip�~�9�x�eQ�	PUe)��ރt"-�ᡇ���ɺ 7�t'J�nڲK~X�X�@Ye��*v��'�m���[o�Y��m;0{�ر�Ni�s��,*q��k���-���v�"˖��CP�*X�<���b5h`��K��� ��h�����Y9�L��nJ֚�k���,���t*�uQN�ipI��J7��q�E��t���f?(yF]k ��d�    IDAT3f?�%+�
 ������� O��<�\wťH'bز�g�}86l؀O?��P��J����&c&@�x�\y��,}��X�b%���++*�N���=^Q�S������%-wޟmmm1b�0
�3V�l�1�܈z��E��M{�J�N�'�Q��x?�� ��P�;0�$S��ѩ�mz.����#��A�leS��3o�!�#����]�#cph�KP7�fI���us9ͺ'���Nl�7d�p���?}e��.�<�+��r�P��	��emRV���ܙ��|^���[ϓ�i:�*�` CoMg�Kkzv���~�cX����x�^o�V=?�ۏ�����D�5�CtI�er+�df'�\���\M.e�-��T�\qĳ��"J���]��/@9ڍ���c��,�$�Kv�8�l���4��6W_x6�$�����cذa#�\���o�(�cVd|n����# (�jnݼEf�/��n8�O�,��r��G��u�q���KYaI1�x���Z���^+��\�v�K�j�+e��K2�F��r6/��_�V������!Cp�]����M���l�۶9�G�[n����M:Ə���U�)H����u�蓏)�'7R[S�TC6͆kQUU!���83$Շ���a�Ŧv�ҥ�A�͛�r�͹��b�-KHct�-��y��ښ�j����A��ằ�pֱ�F67U��lV��|mq������KY\V)�G�8�����㥥Z]U�@[#B��T���,�[���'���믿^ѹ_~��^~�~�^�U�����mR�r����!�BEE� ��.��	�Y��x=l~޲���p���w��"�{�w�}*��P@<���TWV���[v6�;�A{s�:e2i�	��T�r/�mZΤu0� R�Dm����B�	8�0�/9�}nUsL�-��� ���3�%+<I�Hus��(�nc��/���\
�:O?����κ&<��X�i����V� 3�t9Ԑ�qRx �M9'�0���(/+z�hI�h�mO#���C�;e���?봓q����>Ǫe?J�N�&�I�67���	Y�ѧ\}���&����)?/�R8G~�܋�7�k�qa���@;�ZZ囹�3�^u��R��2�*�r�R�g��rݮ-t8]]Hg�4ʵ���岆�n�@�f��a�C#Z�l��˦���5Ùc�Ěb��{Z��5Ct-�Y��tM�횦��ɽ� t� 1��=����D7��r��Գ|sPO�	�#4-��z��q���q�5�Me���ܱU�&џ�_vW0�6Z�����'���;?����x����$�����}|.d�Q�c�ht��)�����I�*�~ȩ���oW8ge�$l�����T�T�SIm�=s�^:�-]�Xq���6��~�4\?�83@W{yx�l�&<ރ����C���Nj7=mI�#��Еd�mع{7�{��5��,�.R6n��͛q�y�a���B�c����QQY����˹seFw�����K@_�n���4Xfu4Q!�U%]w#������aņ�{�4h����Jʱw_=y�	l��G�N;F>��<��cHr6�N ��'[��#�(��?iz�f,����"�L��XcX��r�X���q�H�Z����`P�i{����Z�V@��jֆ�k�Moښ��̠��3�[s���7��� 'N��*�h^��tF��Xm����i��=�yO<�Dyn��4��^���C$ǜ'��v
�$�r�86�k��z.^x�YyVQe�hmiB,��C`%`y,[����;�Ņ�d�N�nF�<������x@�D0�o�+v׷H�v���/�?��+�C!�]~|>wf�y
��m()*��Ï@S{���٪��n��SIL�x*�K��H�%��L��f���x�*���{*Q*�� ��}g�?.�I8�Iz)�="�sJ����� 6����Ç㹧�|���f�|�E�ظ��� ���#
��t(���� c?$�3ð�������;v��_
�=�"�����﮻�>��-�έ�JK$k��'�{Z��'@7SĊ])�K�בk�םA��#?��z"�"!��tBX&"��Ӎ��D���C�yx�e�I�����|j���s�
:sl��dK+N��.�3�����%��wk�:��^X��'���'�{�y��3)��d�lְ����ެ�I�r�Lư�e(�բ����1��c�=����������}��g�5>�u�u\�(�D:��)d��>�A�C��0cd2�����8�����K����x�^�F�^�d��i�Q)͍$U���`tu��j[x���qӥ,��
��
��9� 7Tr^	1bZ�&�8%�*�]́��\�i+j���r�?t�Kc��S��K΀���s�<��˗��v ��~>�WW���Bܛ�JlZ�[���ۺ���Ė����R��}��G27=��DY�k�c
A���_]n��o���<�6mªU�d�8h�'c�FF� aP҃`,�>�?���ˉ��o�*+��{�>����k@��Z��H"�����A��v���i�s�I��R�W����@gwX:���u�V����;Ď����oK�.�m�f���hU��5�����LƬ �{��,�D[�Z�yi�ӵ,U�;��
������Ce\�cw&L�����ض�ضm۾c۶�I:�m۶m��=g�g���jͫj͹�QQM+�����M���X�%9���{��?�c�v��#Da�ɻZ��v����i��y#�7=��=B����Κ�׃8X�`���}!���mʿ�GG%�F�Z{�y2�v�m�(�@2)��gq����7]'rЗSUt�_/��X��O�5�Oi��e���{uyC��Y�!>���s�'Ɵ�#E4h(������b���*�����R�2G�dӤ\���i��r!�߀��*`�J�q�t���^`����*MM929H�u�J��>����v��+؅�6)��k���s�������2���#�w���[��|�ܯ.ܛb#�xW������Mr3��ցX�T����y������U�ݤ����?���+U��`�OO��풗�c����r6:z�����#C� gH�pI��",��`�-�i١�7�-�\���bv�G�L$�<�ߋ���X�߆�_a_q��)d?�+� P�{��)��S]Ԇ�h/;T�kU�Tt�����l!k��օU5	{��Vʳ�K��)�}[m�v�
��Phr>E����1vZ6���[6hN�ǥ�Y�P�����?�=�DC%�dyt�-K봌�Z񰳲n�J�$E�ai:�6��d��¢q��B����]�.������7V��>����pL��ˍ>	[�#���(�q��e�u������ym{�8 Aa�����B�^WD^.ȍl$c��ƾ"s�C�]{�OPo��#�/pe�ik~[L��H��I�A��%�{�)A���E� "��Ll��U�����Gr:�8� +p+�w�Q��%�m5��^��.���҇yXx���6G�8}VC��*�^�0����]��L���k���,R�ب]IK��/{�jv���藄&�6nLx'�Y�<В�J��kyin�EM�bb�}wnE���z���骚R6C� h(��Ϲ�����aP���Ա�;klN����IAM��!�|�͗}�v��W���vDǍ߯�e�D��K��u��Mu;X�n�7"�usc�P��"&��jQ8KmG?��)�X]�ĵ�鐨
��6I&�LhD��JT��}�C���?H-�ވ�:�����n���%k�n�M\ॆ`5����s�B�V{��Z����K]i�d0�=CR��Ӏ��l|�:s0!:���s����N�Jȣf�d��a��v����Ք:��K�g]yj��6�@��E��0�B�럣���}�a:���?3�/�ܔZ9�䢃R��UV˅�{��c��t����-K$�?u��S�X>N���c�1\P�Vl��܃�yx�k��>@�������B���\G�x�_�巑�)��+.t�>m��稊���'�Z/��r+��q���l>M�op)(�B�>锁�̫�H�P��F����w�v�Y@)fs6��{5tқ +j=�h��|Ey��[��LDR0s�H�u+�N ��݊L� |Ʊ� ���M�긽�Ş"����v���o���]�c�a ^)��`�,�aw�+HI��>[��C�Fd���3������Q^Z[�-�kHz��m'�h���ʺ;7���*V�g�}2�2����b����%���C-�i�+B�X�J��	䛻����U�����z�4��l�x�θ�v��Q�Hԓ'Ci)a�\p�_1�Ѐ��n兹*3z�����.`�R�����o$��P���. �M�d�w�5R���I�q�~���Ǿ�>@����*!�O���]+-7���}��eGTX9�rX���Y�}�5���ʛ�csat����`p6��� Ps��/o�ؔ.��R����p��-$! ��~�-w�(f`v��s���"=fXώA�g+�[*=� ��vy���a���L*Q@������� ��wX�%�- h�v�I�w~TҘl���1��$��w�t��/�0����UR��2F�<5W8]��ct�FF|��L��o#*й�{hB����#��kvX�h�x�a�ԛ>eg���"q��mr��~��,��.��߅�Mb�Ń%�Lk�{�>���DUY��c�v##p���T��@s��M�Z��A�-�j�x�� �*}�|��s��6�;�~Eu�@��D���@���c%'��En7�y0���v�Q�N���Nq���4=U%�Z��[П�q������T�n�[�Q�g����elxyi>�ŋ[��c�F�T���Qbfh@�8Z��o^�>{a9*��>:��(cx��3�Y��+�h�I�?�U��j���dK6	K3Wv��<7К��YF�q����j�$9���i��<l�%"�B�X�����Ԕ,PC�+��Nx}ږ�Nb�פֱּu���%7�8��o��O+��j`?O��7��a���g/�`�ND�������-9����78�%-5�C��T�L���A~B��_h0��ڪ���"�����I���ҩ�a�u�(]��f+�߁��h�B��X��(_#`DJ*�����av-����	�m+���9� �]>�>|>eɷ��L��{�{UK0#��'����Nu=~���&�KT�V��X @�%��r�`O�Q1�һ����ϴ�#��%|�ʼ������	l���[����Z�7��VסOtީfm?���E~���9D�.�b��M[U�j%�ŵ�_+M�Sͽ}n���6a���0m�WпL�ͧm-�@��ޜ��8S�e�����O�i�#����[�IO�L������V��EԄ��:�b[[;Aq��Q��������_no��ûҪ$�v��Ai���q�(u�K�"!Z�ø"���[\�O,ϳX��Ⱦ����w��A�F��4�~��"���h{�p�r��s�u��)��B�F��q&5Y�T���Z�!LzI�<�DjN�x�-K�3�W�kQ� ����h���=	vXI3
J���M�fh�"V�jj�S6��$Z/�k&e���Z�Q��^;��<�X:��]L0t`<q���tm��b�m�_��OϏ -�����N	x�6<��(��EKr~/`Z؊r����5g�q�����u�����k�~ڒjE>��	Ov��4Z�$�µy��J"ɶ"R�^���ſ^��o:;NV.��4��U���l傒$�F��>͆Q�䓑�L+�i��\[;K�|n���I�zM�n)N���f�5ҫs�<5�ҮQ,0�!��S*	,)QT;�!r��3��9q���3cDw�[C�1b}]��%����R�Q�E�-g�_zel�Z0��p �=��^�Ў1
�47�m��|������?�A KX���jx�9�)#��B -(5�=P��4A]]E�i��1��80�aq���f���"�TvL����%;1�lz�֚���f�.�(ZS���ĩչ���kg]mrD+�R9����%R�� V�Y�Y� ��X�ݻ���	@�^EE���Nsgc�S��E�����]j�^�n0[?5�+	R�@(�h'�������d��E���V1�����n��&���k�ɥ/E��E��s��[6q��2ۤǭ�j�m���s�7�I�SbzJ������b�����~��4�W��0}�5�G_�	3��iSָE]ٙ:���=<���C&l�"�m�	�JZ��t�]�L���z�vp��mi�7��P�>��3:y���j�;����w'�^�В�#���Í���91��n���sMOP1U�Z�(**��,��������@%��J=lb�_�*G󸳗�^2"�$^���;�r�F��6;	ڥPv�o:����:�5,哼c�G�6���D����tS�p��|�l �3�S)����59D';�D��Px�8yK�U������������g&����� ���w�N��[��;�+=]�-x.��@;�%������/lY�`����������?*Y�����͘��fga�ϯ,�@�r|{'��S�l��	UgV>(Z���H�/�j�R�{0ɩl��µ̟�t<�A��(�d;sT���ŕ��}��c�KW�S�c�C���F��
J�5�'q��=���-f3F!V4��$��C�.Bێ�ϤR�p��Ǘ���Q� �_�>�w#����}ӷ�UR�i�c&C�َ7|�xO�Q-���
H�ʨ䘜�F�bP(��k��L�����T�/AK?�d��))]d���1B����U�$u�Hm�P��`��t��u�f�//n�|���z:����V���!��Z��W�
h�	��?��\y�HNĜ��-�P�T��g�8�&�������(TnC�>��$P���R��81ʏ���m��n7�C�L�j��΄�I�O�_lZP�8���M������a؀�B��>�N`�v��	އ��"Y�4����u"L{M0�uF�; �c�\��n�2	2�AP���M7��lOrO��o��J�V	�P6���@V-�2�p��@J*���4��g�)���Z�y'
Q�ھ���h�yN�ϗ�[|
ˈ4�`B���b�Ki#՚�pD��j�5:�vDS�;��C>7���"���D�U�d�������&�}�.�K���40�	�_ʌ� 3,T]-Q~�j$y��v@FL�;U,���Rti�@ F�/���x�}J����CM�
KE�ld��qߡ	)��)˜����ge!�xm^	�5�̳60/��UY'2�]e0�-���vH���`P4�'�~���@�@:wA|�xY��c��`n���o�h�|t�H�#WB�K�mx�*j(5����v�:����nЀk��n���G�p6V{�@GR��	��Ԯ*���[����w�1[?���%g�4]��
�8!�i����z�I��F�|�nn��
�·����zu�K6�P��_��uk��7@W�TË�_dپ��8�`�X�'s�ijO ��2`8O��$�/'m�hݷ��wtC	���E�����_/���S�/{u�#�tHӂ6X�t3���pM�O:R� ���SXq!���>c�Ԧ�P���*i1G�%=,0��r�q��DĆRuh5F4ms۝N�҃^�X�fnф|���7�����j�����b�ҡ�[�,>�Ӣ�y����)5�p	�Qq2�rC9���L��~���p��ys��4?�E��K�`�xQ`7*A	"9u�V��d��#�D献��s{mi	j�_�/������'c[:��/w�4����5�ۃ�#����c�]*�K�R���˾���#�����zw��`�@ɇ���%���4t�����I�LZ�P�r��8Q<���Kg��L�'c��ET!�1��U�s���N|/��mul�Ȕ�&OEN��ة�޲�}�ad]�;���-�Ϝ��o;�t����x���S�o��`�rQZ�8�Ab�� ���Lv"Mأ(m�B�Q"�t�n�?�N&�e�{�z�	�o��=�����n�nLm
���g�K�%+�%N=��ߙ"]�F�l��:+�aV\�v�T��
:�F�|Ԫ툯oK�� ���K(Nc���5�k�<����!h��
{ڃ�D<���9L10����,���Gu?.�͜��ȍ�B�W���E��_$=�`Ρ��_V���:.TP��P�8�&vk�}����W���RMQT���G�RI�1݈�X�(�0���S���ݯ��X�m������L��q�H�3�N�7*0��%��n��Qr3k�����qÑ8nw�����D۝bwJ�x�h�#j� �5�D���O�����	��@������р�s�h0)��R[T��?ߺ�>�\1z?�� C��ٍ��"y���+�s��XR�(�ҲmK.��)dֲ9�x�r1#z����<�u0G�m��|�`�?-��r���?�ֺ��;�J���2���2��Ño���9&�!�2�?ݞ�t��Ziܦ~�,�Ԃ��rjT��Y4W���)E��d�Ur�.��������j�2�.��I���*��{�ހ�W���Ŏ�NC��j�</� !̬_�iuDD�f�;����Ϧ������w⑀I.1���j'0��uR�sb�^(��?\�|�)�}،�}�A�~A���jbʯ�<�U�����)�k�dF��{��+n%��z��h�4�N�P���B�?h�@�'{NߐH)46��0���9"����ĭ]QS3���[�
���D�UWL��V��fp�ꥐ�OM�y˙�2]��=ӭ���Ft2��O4��u6����b�2U��p�Dy2ieA��Vz!O��	}J>1�D�A^�ٖ*#$)K���.Y�X��(S���4��%����1���dm����zT���ـ[(Y�֡�'ʫ��;�f�ㄝQ�N�6�EL��?���e�՘�8 t\�i��w�
�����k����"������'���Us[����{!!���W��z����D/��r�u3�ܳ�fd���/2�U�⭷Ս���P��_� �?�E���h�
(���t� �X�T�:���A�[<�i������9���e�f�"vTհE-�G�
&V�g���J�*��TnPv&hrN{]�����T5˷G�������4�r��*Iq]����h�
�������ȫ%D��@��|��nz� 'w�p��S�S��y�b2�s�b+���x�7���Bm� 6ɅC��!BM�y�v`@H� 0��4g*�N߲�

���T��s�q���R��O_%���X�u��w f�YoE�����RY�~d�cn")�I5��.բ��iU>�T=�d:�N�k��%��aW"ܔԽ8+����v����QÀ�M��U_HR��0����5*1�3�c.]��.����Ȩ����  q+T�Z\Y�A��	��.�Jc���9١׍]��*,�E�wA�o}@8c�K���	q�v���c�k���儾���t���:��D���>k=m,���W�$E��_�@���S&vS���o��V,�`,�h$���"CJ2D� /FS��= ���9IE������h&�ע�	�H%c0�}�+QR�0���g$r�9H��=o�Eu'����P��ۦ��iTۼ���9���F�K��(�B�ѻ$��hRC'l+_yˌ�)�d���roY�mH0��A)���3<3Vا����� �1\N�>�4��G��/Z'[�-I�s#��B�k�:P_nj�kll���eW���v{4L�q߸I���>�^A�{�e��?~�9��c	��89�a.;N�8��2o����h���k�����
"�K0���3# �����D����@w`� �@�[��O�R�R�Ik�l�z�n�SYd��w�ٴ��8�Q%�"��r�E"���ev��@'�ɕ��@���N��3�I��`�Fh�]���;��ޤc"D���" �]\<�=k�G$�Ť����x�n�-���k���nle�y�ٯ�)�@��q���] D(�
���v���u��+��N�B.7v�pr�E��r��^;z"̔�v�
�*P*�I;���->EB�3H9q�(}�*���ۨ�/=B����gc�V����[�k��Σ�dwS�6x�8�(��<5�֣��ge>9E?����e�p+/&R<��Š��(*���=- �OyW�T)�Z|�=F�������qg�^����\�����S���\���'rQ|�ta!#��J5����Fsx�K���h�K������Lp���x$v8�g���g+��sDwU@��}���}˕�k0"�j�_tV<��8� V�ǈ_�<`F�$n*�"����$r�-9�OY�����^WP�by1?���^�c/��>_���o�$*�ƈ;X�D5Z}�o�+C�֌���$��U��jP ޝPo���a��"��&�\���ｭuV�8�%�tN�WMLV�Vu)�wC�P�ӕtպ�O-'���Ds�'�A�ElLA��m�r<{�|��-��a�o��VFs�J`�?!��/1�c��R�Ѕ����f���d��$H���:���lf����+���!��?��6��~�Ol�a[��ݕ�+Ͷ��՚2U7���ઞ��/�57�=q��;SC�Sg��a;2JE�&@���V���{ц��|Amdr�N�uO���� J�
��f�i�u�Ʃ��&3��{��o@��IӤg�/��tP.� � (4jgJN��^	\<f�|O[�\�|n�ݖX��G l�0i��LZ�m��pL��ξ��ԟ��ǤR��>w2ڿPٺ�[��$��$ԸN�L�'�)�JA�A����vq5�m��_�]	M�%C�J���&��&Čo�Π��#�@�&�����C�����6����*��;���h���я{ZL.͏�`���5t؋�[��>]��0hi��+�������pV�L�a�ݬ�������" ���e��O@J�d�Ü[ߗi��;�g���z��w��I�Py���)�� ��٧N�ۜz���m����4������f�c:��M�����e�.���H�OD�>
�Ǹ5$Q�Z�l��A���B{�����.��gB%�a6g��'fޔ6���A����f�%j�X��H��C����fۏ��9���қ�1ww����0uʸ��Jb|0iM���+k������/�G�4I�ן�eS��x��� �a)j�r���
����+��i���ד����[wS���y���������FQ%��ػ�=�ޭ��k���9]��M*��*�f�^t�by��ll{@�h�<���\]�)A��0���jB58�vr7@��`:X�����ц���!.[���v�TѸM���aa46��2�r�&��mR?�3�~���^�i��Y�_��>��PEA�,�SN� Erf�[A��J�s�Sވ@���*��.i>�V84�����,�^�?�єG���k�Y��P�����9���Ck4���FuF�Q��E���vX#b?��T��ӱ�#h}�����y��	|����/�B�y8=��<�{;z��vU��o�B-���PO}=��KT����*���#Sx&	���"w���Ե�,�%N��7�\���北��5���D��zqq��G�ZE4Xo��9�|��	)y���d��F�/��6��\�����`�ե�-L��8���>�*���w��΍��;jfv�>�?]u�%g�0q�H6��-�y��cnW[H�������0և,���z·0������:�t4Z�Yt1~��?�P�Wp;b����v?z�Z�� &�4��r;hd����D�eO*f!�V���&�R�Ip=@u*I;5���?+}��+���l�ƥUz�:_A]I���]�6\�A�w������"c�{*8���)��T��ǳ��ަ�Jä���A�(�6Eu�N��6�u��"�m0L�N���*�yLD!���¼_��|l�\�O��V��h>xp�r�",��W�%���+�e5������?���ݛy�����m�l�Ag��Sⷹ�1�V�/;����+�Le�䲊��(��;W@�z�[TG7Q�%Pm��3�d���;�1�ۅ+�s϶e"G��&g0�/�M�����w��.|n�ǭ�a�8A�5�{�s.�cऌ��y�Ĳ��v��e��g��]��|��?�yW����F��E=h<���[����y�r�o���m΀EA�3J�B����$4�l�H6Y����ب!�ߚ-�p�%W��}N�����}�M��̧�����q���Kٰ��4a�����rc�o�N�,ʭs�������)Kqz\���tyi.
�R�)�ɮ0�Gp��?m�B���Q�&9�&�Cz�����r=kΐ::A��;�O@�Qd�Y��H-�a�(Qye;�T٪�j���v��g,��xۇH3�7���zJ����Ź�m�x��)h}�/veq�?�d;#M�\�M�5��sC+♗��R]�r�"�z�n�nI�@����RrN5M�Hvyg|��EV������X���z'���	�}�ޚ�l��е����X�2��ۙc���2z96�eA�p1|��Ǜ$�pI`��v�Vgg)Vle
+3����WԪ��sٸB$sd�NY7'&�Xe�XE&����h�4vZ�g�˯(�i-g���p4��q�ư�ܞ4�+޹��7D5,,h�΂#t�3�S>a+>Ն)��+����n߮%��Mv�~�rZ�_WS���w�Y�Dd�<�~�7���lq,��j�'�������=4�0����}_���"�a8��=*K��Z�$�p@=�p3q���"��sŸ�/D�R���ğ8�f`p�a^�B0�]�4z�N�%��㍊A����U˯��.oɜG$9�Z�>��а�z��,���9�qz��j�(�a �3�{����>�71����#H��p�~o:{��3����އ6�6��E H�KH�!�Z���(�*�$.�Y����ޚu��~������tC�x�Gst@��߸g��%�]��V����4՛���0���9OZR��:@���zb|��Nd����6���t�x�m��7�RKS��̯�Z^�]��{~�Q���6ן]������E�b?��:�eu�z\�{JrD��㮟�}��B�៖���b�:v��WFw�����R��*����_A�K�'�u�o�Sy��?�d��p�� ��;��K��1&�1D����#S<����;�N?)ݥȞ����cx�f�6)��x~����q��y�F��}lf����P]���QYx�ޝ����p>��}�)�a�AA���Awq�h���R���"�mb��񄚀?�x�m�-���O��UE��r=��u_>�i2{v�j5�s�_���W��i��m^�e�@��c"�������J|�����J\.O�x���m��f�㡤3AҦ�Բ3�F�eOL^��ٌ�$��\iVe�l\I��X{�-�+�}��������b� e�sR���&yt�5x�JQ��F��	J�-�� "+,��-e]�{T<������BX��u�/��j� ��Ya�&IT��`~�MH<h=/9b0��޼���{v�����i�&:VF��D��X���ee�w�4��V'��I6��~��x��	�s�~A�Ci�s̩��eT�M��$�22�[�צ�۞o�䨛����q�¸�!�P	q|�z�f- ��WZĢ���t�l�U�:��ӛ+��Q�E@z��n�0��Zl�C�5~]藮�t�g�d%.��s*��ݎ������u_/�O���4dB�M�R4�3T�	K�:�:}�^.P�S����&ޯ�(/�b|<~���H���y�q�V�i��n;Jb��'��!x��_��*���$�;��-����^5�$���1����;�
1��3m���d;�H��m�����"�eΓ�T����j�A�&Sl:U[[��b� ���U�flx,[v�Y�,�Ma�
 ��n_к	��c��u �T�/!�& �d׷&&������iO\\�;�#Q��	�g#��c���"/��F���}y������c��`�7D�ۧ�8O�b���{����s�NQO��7}�r�,������g��~����rU*�$��{�4�(�Y�$�ow�%��l�y�k �W�����=��יi�C;_c?Y:�6���~����H����ƚӁ��#��D��Ql���Mj��6�΢���G�\?��G���[�>8�ƥd��Mrm6[4R{N7��):��Q�{k�e	���l��3{��`�<Pi�<(㭗�o�`�-�`�Q��F�i����;Y���9�&Q�UO�C����d�akg� ���?u�#�pF����N�i�2���]h0�~�db�ja�a����3�:�I�Fx�H.��~�/�{��Nv>:S�?7�@��b�Z����o�9��&O50����ʮ�10N\ﺿZ�����Г���F;�u���ѣ��H
m��j�������m�3;�&Y#�D�?���8t��77|��wc��|�S��G%N���;��ٓS�pǓ����MZ�_oYU��W�>�+�v�oXW1�@:����{����"��D�U2��i�E�k�w���0�Č�X6�%m�� ֤��:�dB�*:;ei![��q�Ҋ���I�Y7V���i�m�;G˘FS��CО������%�3�,��R��<���	��3㰣���9z+��s��� a-��dfei˒����Do����iA�~+I�����t�����F6"r;��jq1�^y�mgX����;ѷ^w3��4-W��g���ff�U�N��f��z�Nŏ�Y��6���2f�Wn��!���{�1���WII�6���F8�3h�'Vp�X�)�˂b>���L��^J���c�|�}i�ͺ^��M���RD�0��oixԁ��T�:��d�r�{tc��B���PY��fz:�����T�<^����=��
u�����߼��F�����XWx���Yr�k��Us��t:�%�BaQu3����I��/�$MG4�G��J�8��[]���y�����E,��(Et���jE_��؎�����|�sif��¶j����IXd�����#��
D=����I�j��cg!X��]L��Ůx�8�-�"z���)?51]t��g�����ކ�񮻝?����WH��'Mh'�C����Хh�Ʊ.���쿘,�"�YF�%Ѥ80��GC�&ʵ�-eԳ�n�ڭ�.�-'�<�Q�����[GG���{�\OaH,��b`eȺs�J��E��#D�Ǥ��բ��4������iX�RB�����N�h9�)�)�ny�=�����wk�|����
�`@����(>�</�v���!��O7x�k-Y�y7�0�0�S�����2V�u�8���Mb�|�:�U]�렉9����fa;�x4S�I�,�@���n
�cxM� 2a���ef�/�U	����?�����_�?w�7�?��
nKp$ۖ�����O<մ�e�}ؑ�x��~˫W�M���@Ʀ�������.u�ƹ*�uv�;���r�8ظ����_ޭ�t{4]�Cs"�"��Z��"� �S��6���[E�<�����m�.$iZ�K}��a��39M7z������]�"r&��R'e=��ǟ��
����>�)�-d��d�ʮ��f��m��~lZlӼk:P��StT�^��ı�P*��zC�*�n��x��9���!Zx�D6e��.�^C��7t�P&Ӫ�����a=B�>�r�w�χ�`u��33�����,�D7{���?�	2x��9!����X�K��	�O�w��,��|�y@��ǦS�:rt�p>9�I.v��eJQev:��P��a?�E�V��9
��x�ݻ��=��iZW��1�)���}�W"1����'B�rp�E �������D��-�� ���З)
F!9�+�ɀ2)g���j�'2�3���Q��Ң��~ljk ��AS���v�y�89#�g�&=��U�y(l�c����W�>��i4����W%���RMN��S+?R�_
�E�
?ݗQ��j�V��D��/�	��]KW�����8pW ���3�f���~.��q�(Ļ�瑭��UU�6ȅ͸x��������������r��#�u�d!̃D�j7��+�G�`&����|i��x�ad{�~�y��D����}�v�nV��(�6��'��eb݌��3Sp�_h��؈��ny���u�Ʉ�x���<���t��5D���b�d��A9���:���qvz��6�1���i� BCދ����g�y�&�(�)"�A�4������2����>&�n޴��8��O�i���X����V�&�U�ؤ"�ګ����Ω�,!'.��N�'/$�Dn;h�2�D�q:��j$��j���u��;I�3[�����&�d����й!ҩ�V| fN�}°ݯX�J�%�L���3Ϳ�����
r���˛�D*������w�&-�H��L���kG;�
�]��v����H��� �] �56a1�.M��p�y��[?\}	.+�:X�*	�?93:L�0�^�bݜMn,�ӡ$:�Xn)V�-�=�bVA&XA�UƐ����
�x��qZ��i�j��M�=4���g{!1&��u��:&�J�KGv�`G
:�V�Π5՜��&�2��;Qx_�6��{;�j]�i]�-<�V$�5�u,#=��L;��}3��A���<���$�������-�YXb��ᮅ��+\sv���]z��G�)�$�?���Q�)P���9�
�\4^nlq7}t�㫧�����������:��c�Í�v�����FmY�a�+}�0��@C>�Y��y�!�]��>_οx&~�#����W<�`d���;=� �+QFLZY�����Y��R��X�pmvmc�D��tO][�Hx�W�d�����������h��(���3�
�w�ç���Ⱛ���q ��c5U���#�d�j�EC�@���3��as��}!�� R���x�i�Nq���V����$�!�'�mLZ�| u^3>���dIB�wo�&���Kd�ܐ��?��I���jD�*�j��#a4�M���T콟�G*���UϞ���܍z�ʯ�>%mL��m��.�{��F�͡��T������Q> ��L�:r�Eȃ�6C�t��e�^�g�}'����'^���t�K���M�m��v�X��tR9�4o����U�{��rT����Q����a�������1�+CWi*�
	��N�]"U�,�"#	�{UŸ�t��5��i�b��KQM�xzL��~�1�����Ԯ.�K��R�5���r˥��έtCu�e>��/)(
h�@s9����f�(E?�ޒE=�?����S�<�5�m�{9}�Z��X�g9h�e��9[���#G��|m�.H+�O3�F�u���y;�8��1��si(���=f���	}��Ӈt��Y��`��ȴ��0���˦3�L���A�Y)�� ���S�������6�iW����2�^�*3꫊O��ɞ�#��ӡJ��P1���/�.W���j�Z���6��X9[ ��v�bj.\/� J{�$�B�������1�=�����o�a���~��e�f�
��ɰ�4N!�g1j������̬ص����B��w��V��#Z��*s�1]Z#�ȱ�L�WϤ�8��A]�s��v��O<We���Y�W~gO׍�E?5ֈ	�3�5�m��?�������-�_��Pw2ao��t�@�'d��2����'3�=��d&�T���`o/��߼���\�'�,���?YBA��\�����+�Sr�$r?z ?Zj�&��0H)�(�rJ�?
Pף����5����es��|��w�)�)�x���7��V�^��o|�pf�N���|�~q��ҽ>�\��Sf�CH�S^6�SP]���I��:�hhE��2���ys̒����$����zЅ�{��U�d����h�=2��b�'b�vg���}н[ʏZ�������5\��w��O銆�1�>Tf��q�=�	TM{>/b�%F'���,�4��>�l3���4ߢ派jmd�lj!��Y���v�������0���8~�|1s�P�u�.c뚀��Ϫ����zd�3om���w	�a�v�&����\t�;2%������tz�b!�A���c5H>ffy/s�= ��Y�2�ir;��SI�=P���Ha��ve�\��S�n�7g��Ke�<FQδx)��s4�.?#(���9|�wH��=WnJ��[gp9�
�v5�9K<�`RSKQj�Aq�^�:�<��`�� �� �S�v"��[2#Ri"�Vl���J6;g��e��S+���K�ۿ?��)Lㆣ�\�㽋$���B�g��p��u:7':���&~�;Y/H�)�C�9�5)��3� �库v��D��� f����?+kb��G�,�d��L%gaP$��Od���:q�z�
���;C�r���y��C���.��S�J���m��F�9�Yr��2�����}�.�f8�TR�g���C�]+J�lxxf8)�iA�{��թR׈����k:���OFǷu���̡0�n�m�9D.H�*2�pȵ�ɗqP <Yf]��;;	�OA^�!�'���N�ch1�Xy�q�����:���62r'����u��G�m|�oc�����-T��C�i�r�@����哔�	�)���3v����x�؀/S����t���k��l�_���(�����j�ES�5.Ī+h�֦B/[�تV� �(���=����6E�_��������y�y�_�'�s^�u�ۨ����;5���պ�췜1�'��	P�/N�,ng&S���B�}�	���.8K�=/��|�6J�#z�=uJ�������T��#nϗi���n�v`�����4��SD�[Ya>p���c�/�U(b+q�W�p��!ɏM��{/���:��T�* tu�L��Į8ziF��
{�/Ӂ��~y�fv�"gO�>�En�At�/�ki���;� ������	��>�������!�ɢ�xƘ���p?[�qq|�ʷ�C&��-K쾀�J�m26�1^� �8zhxh#�]ؾ�	0)VR���o���x�� �B����~�X����r�F�,���E<�����\\��٥[`=�ך2北�oZF`��zy�c��$Л6��Ƴ��1�̋o6k.��"��6�;�a��O��ߧXn�$EV���r��^�ƙ������
a}SԬ=�Ɵ\1�Y�?e?ӳ�:��]��Vײ4�Vf'"��渽��ᖲi�v������w�p��ϭ��~���io��z���Fe���=%�LAJ���Q!<5�ۃ&�Ra[ïZ��_��
�Q��7�?�������[*�v�ç	E+po��}G�wN���h����~T��<���PtbEk�]~;-T�a�YkM�ũ�D;��,);�L��Ƨ�Ie�[Ͱa��� *��i�9þu���TNc;�����{�W�?��sU)��	�V���W�$Gy6ԋx��*�=L8�=�V��RJ�"�}� [ðt�&h"�
@�+������P��@z-��5W���{'�|<_�+.��=>N��]��X{G�}on�F�x	��a�p����ڠ �%�u_��}-���ه���9��b��^گ��Yb�)W~΂8|]����͡�>u�e��� �u��`�  �C�p8Sen�b7'q2%^Y`^�u�ܰ�;����]놹Vj���2,m�Pk�nc��Q}�Yi�{�'v؆��..^d���t����@�4�t'�������ŋ9���᭐�M��FL��R��/���BO�SL�Js!-�We�*�ݥ�YΥ����Nԃ8#g�P�����\��r�S3ѭ/������)a������=�i������+0NEP�}�����zχ'�vC�[p���\1�}�̄&ɼ�4;�-G�� 6i��o*�t��U����y��ԛ�qtl�!L����[.v����J�`���Ô���l���z/�P~^�\S � ��H7�2�����}G8��>����F[�9!�7�{��$?��ڥr���W�ހ�56����?{�����q�TZz&���R�|�� ��
O�F����Nl)Y��<��	=y���� :B8���m��n��8�����R�|6������C�g�e���y��lcq�x���v?���;<;��e������tE3M�!TtlR�t*��l��]9��r���U�MXu(�IzzcZ����NɍF7ww�Z ��«l�A1��r��dt�l+��@��R���l?1sH���?,~��qP|��A�k�B��j���{���@�Ht��K6�D㕟�
�3���K[N���T�?y�P�7�o g|���);W��L��=f⓵�Wc��z����j,���Y����y�� ��[�D�~����9�]£K��^�����K���U!�J9�C���C��s �E���P��J[yޟܔ��ւ�K����ƒ��Y���֏��+aYV��˗;3�ᩛB{P"�yӶՑC�Get�6݃ i�4E�o]���������u��]ݟ��s�ԗZrV�[����>�r�
��G�����MH��@���~��)���T*����s���u�m�g�sx-9Ki�ōL;s%L�3��r{Y�f}�������:����=��d�?��Jߕc�1�h- ����ݺ����	/�lGc�߀����,N�(�F������d��|�'�1���~�=�fc��>^4tf�V�����YT�;R�h�N~Ê2����;��?*o��
�;��^��\{k�u�����'�.�KK_;��m|�O��0�5�^�v,e�!HM�n�#�ng��Բ+,dQ.��a�]��qz,�%��`z���a	./C�dH�ţ
�H�B��z%hn����,f3==�rO<h�� )}pno샶�.�0ӕ�Spp?\��������S5ШC�g�f���I�;//��R�Buh�K$EC� �#;f��+�ާ����9[K��Y���;��l�1`Z(>��Lj=�n��X�;UV��/�M�Cٹ���W.^��د ��ُ�0;16v���	��¡Bj0��`[f4�5l��3������T؋ N�h�����a�N:]YM�����5J��@5c�n+r��Wr]K��E�_��#�
�n�=\�����+��mʇ��16�2�
��ә��� �	X�-Ɗ�PVȡ�<K�\���#4}�A�^-�%c������IԂ7�w�21c�*Y�}:T����)��wv�!��ph��m%^1ҏK.���(��w�`�}������U��zjH�?�����y�6F�)LfSט���[�����#Ż8^~%��f�nrȪĦ5��)�O����#�f�n]�uN�TT�٬�=/���M�{z�gmX�I��d�/��	�v����8���W{�7�����<&Aݥ�����i�k<�eK���ns���(u�-z$�l��R�9����O�����\�0Nv)���4��2)�C>��[@Ox�P%1�1��ܒ7��r�d�K}�﷖���%�H`��P}G�k�"�� �0�8�z�п��_�<��՜؞	��+m�S8X��P�S���导(�$�u>�J��W)t���U]�4oǚ밯���iC�(9ܒ�ll���}���9n��!c~Z��]��P�j���c�ڔ_��2���N@�Bd��^��ء93��=M�� �B�#��n�up�7����B��^�|�<W��6~{�E�p���UJ0���*�9$z-�d��&��9;X�aj�CN�9�+W��p�6���i#o���^��A�L�����x�F�9�Uz�+��r�oxL�A��I������^�(�{o���_S�⁏:gu����U3n]��M���|U�󹼚|�Is���mp<u@p+l6jo�ƠU��H�Ձ;j�o'�V_
y��ޛYW��3�P:�Ez�ڕ����T-�=Zm�LJ�7_����j�3�F9w��
J3i�� 8U�W@�81����gkX0�iF0؜�>?Bo�C�;��{�Qӗ����GF[K��	^V�'���jv���<�Jr����8$Q��Vf�8n�0��Nr�fr���*hUn��I�����1ԭl��G�2�n�q�kR��A��y�z&��=���6��LF!��H�?� �S�]�b���M��'Z7A]?���~�d{O�q�D��IQ�O��I�䌟�b�/jB���\bRN������tS�R�fI�PG��$��m�%M�<MqJ�@�ȭ/�ĵ�k�	*v��C]�-�]f��gۙo�Z��t��8c��SGX���}~*$e��W3:�iWqm��Z��p��+�����&��ɹ��g�)�O��Of�d�dm�XA��G7��n�կ	������6���_�F�o0Y����2��C���T�����i؂a����H�׺�Vg%��ڴ���;�	�wR�W�NMz�5�?�������`[%/���У~���z������gOV��8O�A-ͯ����T߲��PK   �<�X~��k�6 4 /   images/663b53f5-e86a-4272-a51e-f5b809259b46.png�yTS��6D��U0�*�n�4JTP��� ݠТ�
A	CP�y��j��mQ�L�4�@ ����@E� 4$"B� ���пw}�ߟ�ֻ����^<U�k�g?��u��/������[��O$'nE%���W��o��� ~,=󟟏|F�W>𿿦�t����G�ɩ#��/ׇڸ����;�7:D;s���(��_��b�	�3��G"2G))�)	�-�H��[_Ɨ�e|_Ɨ�e|_Ɨ�e|_Ɨ��H�<�/p�������/���2��/���2��/���2��/����bl�9�Ϸ �?��7��S�9gζ���Mт��řv�����'�6~�t�y뽇N�ugKZ����������E?�G�'���O�0^}b�r/��̪�=9�����g4K�?E�d06:�b՚*������2��/���2��/����6�!7������CSoo�Q�ا>�:��3�"�ܾ�yT�_Ƴ��1\�yk8�v~�V�����g���d)N�.�х�I�3L&�}z��U�B����I����Os���:�O�@�bt����j�A��,��YZ�Qr�p��`���5��^Jt�l��3g��g0�������ҀŌ��~~�hcG����a{	|�K� ZZ��,��%�o17�����2`�`�~r�p�*3�������(�w�2"Ɂ���@�hy��ON�����x�*���/lU��b���].�?W�-�H$+
?����%{�1��x�EF��*�2��K����AZ�� ߸�����4@��_0+��r�� ���g��O���D����N�ʲ��\�C����6t2*�vnȺ_`�",������Y�;����Ui-j����L72{=��H�5����CB�:�F;���k*�3{vaa�q5���[X@���n�2T7Nah���-$NTײ�ڐ�����	]�8�scO�*�XwF��)(7�x��xλ��r�	�F��(��s�����1�QP�Ƞ~���4*��M<7p�'��Q�A�����"�t�A���t���#ڇ����l4}����c�v����b�|bTx��DǑ=���M&BI�$������.�k��>Ը|�B���C��VQ	Z���L:gO�]9����C'�K�Q�x��ߵ?^˫�S��ai6Ǘj��:ٗ�`4|x��Ǐ�_�~��*Z�&c'ո����L.����\쓷RE���a���<�g�$ݽ��̈�r�3'�0J�����:=�3#��a+�^�V��65�Lm4�����Ne��w�7S3�9�70^0�͈����Y��K(��34=A�)WB�ێ����%`	c�y��j^�1��!���Rc�	1�'��p�<�M[`L ~��*3���gϞ�~zi�����'��&�\f�1#��4�j����]IG���C�������<^ֹn̎�1;�CvOm4��bD������:����xY9_"�ğ{t{[!��9�	�9�^��I�s7��'�b<IT��V��1 �y��lb�H
�O��ƞٍ�݄(�S@���<H����$��Q���������*�� jA2�Zf9X_c��i/Gӵ�����={6(���������	�#���Tr{��@y�?~�O>����~c/o����J\��ê�Ȼ��sQ�T�&��`j�11�<�C��,��
NW�M��}�*��<�~UhNHLө�����N/M|z�u�~zԳ@��}�<9����>b�F4����eЈ��Ӎ��֧6��0��D�z���j�4 'O��
TL&^rd��z�s��?�iV�c���4˼��i�����^�� w,>�qt=��c�H�����¦�F�������To�z�b�!~ԅN�m��m���NAn�>13��wSEB���H�zE�^`M��F����W +6fo��I(ƽñ�5�!L�~q�"�qP�ܞ̜��g�A��m��+*��-��f����-t�3�B�u�9��`����5����h������;�s�F�,���Ը���3��G_LY�f6 |G�����#��n#�[K�Dp6�x��}�o�=�{��x=��b��r8�r'6�̉������.�\��]��wz�;Ñ��fG��l������mG��C6�$�'��]���drd��ߘ�F�/�M&&�3�/|N�^���7xօP=\�ۭ�
2�hƩ�VS%�w��>t7�ޓ�lu�;���+Qm�YP�����D7y�s^N+/����{G_�\��F����x�|vv6���	e������?lf�J�����ߧ3���_��- �:�~>�fE�Bp�:�|G7ӬEIĕ�@s�&9��ͼ
Q33҃t�b�\v��=��7f��Q�n�C~��^��ӯ`K����4d|c�3�p���2�����|+3���MhN�+v�՝==D恾_��.6��3p	��w�t��(�EE �B V`��Z������-_8��w4ՓL�VJ��gLSɱ�eq�.E/�v.Ϊӛ`j��������]���	A�u�ݾW�jS}RwCu]7/���E##v##��-���x�'w��}M�������r�E|+��Ң�����A�@Ɋ\�Ew�{��]G�p���̙d�a�t��,m�_Ѵ�����������_w�F/�PW0���Idjw/�/��0_:���}��9)�s�
?t���qt:�SS`U�jh�����]��?�ÀBj:�'��/0�����q�<쌮7'Zs��u/�jF�>�U�,�T�;�O��E�t"�qF���o0s(G�FzQ���jpئ�sY�c��'�A��)fNkK*�}���ݶ���ej�W���p:0�
n�I��,��،`T�QR��W^^�>5�9���=��*��U�쩔��mD� �y��z�E)�lA��i��v07��r�m+������X4�;� ��?�ɖZ��הhiSS��%�%X�C,���:\QΏ�$,���.������?�.*�*~XW'�KVw�1���s��C�J���|ud3���F9��{��̈�EZ��B9�If����O���0�O��K�B�W��6Y/�>��X�[���]X�|a�{����x{ژ��~-��b����@W-��z6��
a׾b7A��=m ��g�26����6�K	�bq�H�	D�	��6�dE��=���f��0��܍�!뺺�ɽ�F�������_��Ved�%��<��陙>��"
0v�:b�(Z� �F�����cG 2T�ysA��0-�Z֙�O�U�Db��L]��,�Ί�֫�����J���+B��&��>�e�Y�X����<��s��y�,����r3T����H��ŵ-�ڋ����y���ڨ�eO�Cql��G�a�/cz�f�l������~�����ݻwS�b��,d��n���0Am�:�R 1���L�".?Ƣ����w�j��橐�]������+d��b/�S��E�JlA&R=F]8M*�.�Y?=�}~W��ѣ3��l�t��[ I:_��,���S�NBG��S���Y���"��o�E/ߙ�eJ&��#�1�% �0�t%C��y�n� �G�Z�="��K���LФ����?���;�`:H���pc(J��)�`��bL��ئ�ZW�c(G��`%驲v��j.ڵ��������B��@>���k���\�7�,�h��յA��{\56P�O@Z�'��!�Ȭ�@r{��H
ڷ�K)�!�L�� �;d�f�i#u�M��y?���A-���,���W!��x ��Y��ߤ"Ux[�'(̌�y��Wi�L�DD�u"##�o�R����N���"��&�����?�ݎF�"��p�U�6�E���"%���u�s{}�C��oѳ�A�����踙�7�C8�VO&B=Ȗk�Ҭ��o2�3Jk)�m�k!(�̒Tn��h=K��L�6a�X��Dn��)参��9}���Hr�2�b#"h#���
���Y�bՁ�G�g�uT"���+��Z��U� ?7rX4y������<�vP����u��$�F�ҙ�.�71��
JH����}9 #6�'�@'�tHc�B��Ħ�>:@��xB@��fjY�?A؁��M�ΉN�aY"6W����1N�����=t�����{�Cn4d'Q^���Rۋ�b����Ug�ꔵ����������[�V~���s�1���Z���⩑�S~���'ZZ��+�TFo��O;�pZK�J�$q��Q����U�j�0Ys�I���D�\*sfpp|Z�p�Q��%5Һ�3n���?�Ŝ��{�����n�1;�T���0,Tl�Į���.��oMd��%Q`���ۉ
��빯Gd�FL���=�O��+D������C�y�`��>���D���M65�&ƠV�3��_&g�2����E����A~q�_��j}ʹ�vR(�ܿFP~f�U7w��G��%ݩ�w���J�2]�z��`���-TN�-^=�葆�R��Ϯ�K�7:5Ǧ�58v2/f������\w[f���vl ժ�?+ ��M��U_a��@�y��TF]P�J}��</�o�d�(b�'��Ю�yi��k����t�RI���<x@�bo�w4R�i�z@���t/L,�l��Ż�E��9��#�P$̔�r�����n��D;}6z�:�aC]��r����^�� �ÿ3��:GA���������0p4�A����/>�=OKcv��'Y��>=G��:'XO�}܅y���k02^�-�>�T:�z����~4RN��蚾=�=�x���\��s�����4����ⲟ�u�\kc��e�X��&L�a�_ �[�sl<M�u�yٓ�,�S\��Y�41ܪpk�	ޖ(j�������"ń��>��xG(S<��]$��s���T�؄���o��?���~sÃ�#��= ��E�@�����Қ��b��Ӝtz!b����t!�N����ǟE�ȟNv��������� ��.���ZW]z" 5Z�~i��co��5�b���ͫ�q�y�[	����R���%F�b.�|	9��k/�&.����������Q
�ѧ?1��g}䝍�&̘(R�-i�s����5��W���'���X<��1x��_��'DNM@��tu�u��#�W��a	��������P�34އ�`�'��R��I��!�ꆔ��쓁��t�jl$���"6_k��xqRV`6���l�p��Ю+ Qe� tW˿yr���!�/���'5��c�ׂ�4J� �S��G��#��7�D͑�>���`]o=�,�t�9��=R&�MC/ӭ÷k�rѓglb�jV�Ps7��t��1��rF����A�%\��9:�}����g.>ygo��E���|����n��ٟ�~�QP�4,`	y��7)b�[Jpq���1>��V��,+��w�^�l[�e��,�U!�4�p��l�쪍y�-^y{�9oP�E�f�o���*����͆���|���^���X$�^�e������`M�K�x|,���s�}�Y�T�Z|�~��_.�)�j�̴bī1�E�
zvG������`�\�t���Fz��s6��0b��5��9���~�_o���	���?�h�K��T���k����կ��śĀ`BZ���Ț"��wQl[x���	gM~�T��&�͗�6��[+�	}��&�Հa����0�K��=PP*��0^z�n?����S(���1So5S�Y��E���˜I	��avS蒶��ܓ�/<D�����#�eޙ��
M6$�m'�c��݋9�gw�e^ڧ�:5ma��o������b~v�C�{�W}}����JK�UY�
�Jc�yccc����<U���E���9YL��Ւ���wA�e����Ë=�E�����*	��XY2P) ��-��t)8aKj����ж�*�vk�dS��XZ�@�x�SSr����D��Z���,�x�M�}*;�0p��iqjʥ��o�y1� ��G$#��N�d�zK�2�}(��?�|�u�V9�'A��1B�nG6���kD��c[ݎ��Ps#i�b� W ��->M�,?�'�!�� j�a�[�`�8� B�8��W�/j6��%�C���b���mܟ�:�B{�����������MaA��Cq	�k�
���&h(%p��a��AXR��~dM&�h��uR�������,sٻE�H:
��GDߛ*g:�	�_��[7�&1l��u]�W�2&�MXo�u [ �p����d�Y�C�d>��w2����@+(��T�2�#�@ �)cF�#,0 �^�K���5�j�D"����;U��� Egȏh��}��B�t%}����G��27"�0�(���I%�:�8wGd�fUUպ?���6�8�Js�
��)���-�@�ʟ�G�ز&�~T�C3��^��suc�4�]�ɖ�Ѥ{�"@|3��Q�&�~^o�l����x��%D#Gag��n'�@P
#���u
����b� ?���(���13�~K������6LH^�o���"�Vh��c��?����#5�QNiڧ�NM��JwJ��Z�#�񿃏�7��𨋙����.� �l�=�")ox­�$s�����4�Q�t�0����c(��dJuT/�tCI�Z�kP����my���E7����zz�kC��߀~3��>t�ҩI�� ĸ����T{�z$~�*�z���4ˡ��?�٩�,�w���h�m��B
�����g��]Cc�YT#,�f�L����"�<\b�h�͟�+�5MihWTG�am���E�i���a�B�O:	�˹��y?�dc�a�"�Ƙ�,�����&���d
�Ks�i�@��v!��6�Pq!9T��3�U�U�Y��j���L��2�o�1�ڊ�[z@��������S������lz怒���y�!����������#�v��)�A7��ߓl��[�;=��Dy�d�`����@�W�|�!��a%�H��+ȉ�m�'t��1��0�	4��E�^���l���#̾�ݖ#���yaA+]�ۿ���O����a˶�㫀�ܹ�Ҕ�P���7�U��U�����P6�#w��'J�kC7�a|�Z��XS��A�	:�'�9�*'^<31,��;�NV��2#� t��;O���QpA��%q�'2��<g@�b��G/˴uu�� �]Z<�������
�=|��`]W���l]|{�E�	�V�d+��Uw�r��x6�-��h�����*uтj�j\O4�ßMrjrFHJXr�xX�F<�A`K�P�x����ȯ����T,_��Xm�N
Z�Dr�o릱����cݘk�%��E ��:�fek���N\$ ��ҋ{+2^(kݘڨ����	j&�\_t�vJ�Q�@ģ�v�z	Q�$�
�}�Oj*C@�pC�`Ț�'�{��k:<��q��&�$����;�����޽�c��S�T.dB�2�`�����o(ZR5�Ӈ��ݮ:�H$���X�y����j�T��wj
����.徙}���kTAY��TU8����WKKK�� ֗�|9.��t�ZR�e���D j䥁�2ѩ���8�{��p��I��kv� g{�`�l�%H� ���NfjѠq�:�s��]�{m����p�3�����N;��*�%�����1��;[4zT\fJ&��re<����^܍�CB�5t?����.]r���BI8H�i�4�P�W�(�|�3�`���N]��� !�v����q��<
�?����QX��k�G)�M����ԖO���c�K�k������I.FU��=�YG_��kD���k��n�����
�ljh��&dHۛ�#
��֎m�rA�Am�`~�a`&/�$����bs�����0��˥��6��l�!�1V�� Oͱ̥��#e�����\w��A�1��҈�ҋ�|�����K���_'�E��sCﷀBQ}�\�����I�?k�&/�v��Bv�M��2[R���~mo����z���sf˨L+4ӎ�
�k1�J�hٺ�=]�!�
�Y�����N�ꦢ���0���6�BG�)ׄ6��Kq�& :s��U�#zĝ�țnD��k���{$���}���y:�>,&fn���$b�3�F�T�f6?�������N8^ָ�$B�5(�d��c��g�C�����߂�V��
3'���g�U���O^gm5���@��x��#����_��Pƿ�u`���_	���������Qua�G�0��x�������	� ��)0������{ī�o)9��n]@ݮ�������ӸX21Pm��
H8V:���a��|�ۀSl�)�a��`�
3%�S���'^+�4nq��
W�T%@�m�;7�$#͗`��N`fa1w�C��3�/���%�����P)�झ���	[�]^ܾ���ۋF����ə���t������@����)߿Mw�(g�f{���z��1�~|�H��?�鬈���@���V�܎p�}�?4�3je���^�^��y��pKl%���HΝD��ô�(������myl��2�Uf�sޠSS�Tn#ޜ���>��w%��T���aq�0�P�kk���s�څ[	�91?k�]��Y^��nV��s���Vtm���js{����8�yF����ů�˃������X�����X��E�#f4�Yp���r���\�|��&��/ �S��Ry�~`�R�q���tJVVV&��O��0Ǭ״HGGk����0%�#��VRr�=����$8�mĉ,aW����)�y������W./�/ȁo�`Q�f��,��`&32�	go"�?p�y��V�L`ַ� _8L�rCP��C����U���V�N0����C��D����w��(o�.�l�"rL{[���B��NI�J���"�q�S]�s��G��=�(�yi��7a���B�N�6d�ks�����a����;��C��oa�\<���O��s�7n9!��qV�����P]X:R�)v�����
jY��?˱�@�Mxq]��mp�J� ��L���f�2p7�1\�ূY����tY�OX�@/{
uKEJ��^itgo�v��X����3� ��""t�N9���.���A�~O�p:ل8���(�e| ��h<9�"8��B��M`������CuP~�_���/�����N�֟�V~�}(�KuS����)M�Ť���Ϡo��@�Qx��7�"Vux
j�Cq��uW��x^'�k��l��u���k�l�?��������S L[z�@��;!�]J��)��"E'w�����0x�]��kCE��r�vAX盛�o�?��O P��5���D�p��	a�O�0�9B�� �T��iM�|���[��Wl��5�ƌӉo�D�@���)�խ�	Mt����9�u�E���yi��Ņ��V'>=0���#��!�T�5sZr���������mE���C\���w^�K��x'l%w�t�SS�u�Xf`�~��1E\f���si6�N�G�>jTNT�6��ۧ�po��jGGGb����Adsj"�$z:��{�B��r��>���a<�e�$����p���x��s5����!�9���0m�5�.2�%�z�� Z���Pu��})J��̙x����˰:���W��᥽~ry�_�aY��zJ�"�;dj�i�g��Lk����Tï��A��&۟V�k��=��mi�	�N���;�w�Z��J�sv��ّj�>~�����Y#���{���|j�>�������a�UNv�������q���+�ԸO^���>{�uC�#	�@����N�n���<L��V������e�,����ss�P(�va��֜��'�H�/ Y,����E�/��+�^�v�C�<�mꉹ@2���+]�"��~�KP�5hs�,�/ZlUev�=�����i+�^%�G��}���pa/���Ga�	H��d7S���^�0���d�졉U�v^Vq�`m叫A骏�Щ����(��9g��ʾLf*���R��TH��I$�(��2[��G��:E;�+E��X�O����ɰg,,�����#D��{K��;��B��,�Y4� ����ҴO���R�Tr��a`A��Z	�Kg'\z�^�4�;�,ςb�n��VB5�Q��f�'�0��������^�ϊ��	½��˲r��i*�Z*�s�;
�������U�X��:N�����J.�	�Jm�ވ��E���cK�78�Uw���s*T�*/4B� �_����?`%�׮,���P��o�\���}���G�`~��2} V.�;֠7��~t/��p��f�"�����;v�\~�ͯ���#ĉ�\��;�\~㑮,V�p<b�6ݏU�
v�:��\̮��Y��u�#���Lv�	t�?�</�8lM��aZ,�9��1j,�l�MƁ��cՒS��U`9�H6���|(IP���;*�5��%$��䍃���.���Jl���0`���E����e���!$&8�z^���	O!Z��C:t�=z�(����Ϙ�8�"�`p�����ea+K#�������כ���T&�T�[���L&�771uRyn����+���	����l�p�n�j@#:7�w.�ڝ�K��-����S��4!J�aKH��������?f�1����cR�J�tz�,|�+��lq �l(�W��[�W*NwLaThkiYTayv��d�e_l|���,�ͯ^��ޢ�@�ZW�H7r'K��t7&�/��.}�؍#T��@P�,�С'�Ń6������R�g�d�����u�}������5���.���m�Ɲ�qb^Z
�{0���B��}E!��]�����'��)#�ʷ�^��a�6d��ϗtvuE����<�q�����U�1#��
[���R�u�]��
A:����sNPpp�]Ҍ�0�w�lMq7h%�)J|������w�ޥco*7@7��ߛbq�f�kXCԱ^J��֨Z�o3!�d�)P},,�ſ����x�yԯ�3ն�]˹����]Hk>1��y���9V�8h������a��L�̨�Y����8l�	��Y��oD�K*��P���}���)֟ڮ9�ȘNB���(�N�^i�����7CL����J��$��맢^�4ɟ�Aʤ�*�?���@o�E��/�͊˞<yR��+�ӿ��~G\���������_cƿ�����j��CR��_�`'�k��G�w�<�W*�Y�
���﫽�]��@��?�n��n�0�4�C����Za�e̪��8{�W`� ���/���(ͩ/n��P�b�[�}��k�|-��C��e�c��6H�!�,��Ĳ�^墢H��X(M�%�����MΈGFFV奕�;���=���X�IX��a���6d���;��w#��1[�V��<k+��M�',��{	�v����?�p��U )�@Juφ�:6�
z���huê��| �*(0pޝ�[��{/�ĿW�p3a�N����0�fjj��p�5J���vg�z����k US�Τ�rI�:���ψ*���D���j���+�1�d@\��=��Z�=v]�b+�}�?�k�H+3[_��`(t��ѹC(�ϼ�X������ٻ�{��L�r>�ty5�c�:��������Pيtc��TT�"(
̖�|�;5�֍��"ƹ�艫�*�ހ�u~|�}zL���7q�g\mgF��ޱ�@�3,R'j��Y`� ��,Gk�-o:oi��m�re������-?�����o�D6�]��tn��/����t��i�b�#,��`��B~�X����4�)J���[�e]��|�f[�4������F�@~�B�ʍB�cV���~�Nw�+B�zwd�!R��0����_�f����/������k#Bd�6�i��#��v��x[Ľ��}����M&��ߢ/&\�!0\�u��
o0s�Ql�� SѴ�26CJ��J-�(�p��wnH�^��[	gg~)ĀN���Q��?o��b�|�v�e��n0����k|E�����o8��י��h�; W-?�kY�]�3���v��|�����N���p/A�%O�0���^�Yi���5T�_�4�W� sY![U�xO����9Ō/�>Ü9@��7Њ9���2`��v� �����E��y�o�7H����?�d���[��`�G��������: ��1xZ�;)I������b8W5�dW����L�#���TE������<iψIg��w�Z�R� ��>?2���!O�o���3��d����+�
�T��� �YX� �k5��Y����eh�%8��e�L��^�8U�[����RΗ඗;�F�,�DK=�K�����SӇu{�(�W=;���;7p�f(��ynk�_��<�����9�+���flHI5��.4�)J�6�4da����u�rww�K��,//�
���]q��U�dQ���Nv�q4c뀱�Э��"��7���w7�S���C��A�f������8���#9̒@�`�mh 魗��-t���E�=�ܜb�7����)���=�'�'��&�_~%t(�����l|4�5�;mm����K��p�E��_eÝs0�:�Ւ��Y�r�䮝�j��������Ty��͗��K�ށ���Sg\i�O��G�s"�E��Xa��Z�e8�u3�n��@G�^�I N����*>��蚷�1Q�FLݝ��%CVs���'&e6����oT���cSb勳� Mg��6y8/�Uf�,���J,K��ݨ�jY�z�%E�Ӟ��;�%A7dv3MfUG�ni*#�
CԚϏڀ�x���b�����	���p��]����m��_�pt�&�j�L'c:9RND�I�L`l;��Ҷ�e���Z%9S8/�?��j��}�Z�H@Yg�*�G�<��?ȗ���b7����-�O.3��JB"b�U�~Sj�����<s�ڸҍ�6]�Rŵ�ɾ{�l�>w_¥��x����P}a�4��WZ�3��TB5$AF��W>�3��l�ݱwi�&~<Z ���EW.'�o;����4��g��d��j�p�����HV"[fff���/�aG�-��ɩ�ʉ�#�Sf�5���O��r-�{���t:T�.]X��R�b���?��΋�nooW���5�̜ P�τ�lT=������~E���*��1�`�ҟP�^7������g�����\�!-�{�o�ӷ�5O��8JZ��e>Zo�Ӫ�ԃ6����te9��B��tj*�B`zr��c�0>��}�ǻ��sL:?8�����u/������d	Ď�z�X�;�������^g>����춾Ɯx�����\5\�)c��7� ��������G�U`�
-��zVR�Oh+).��M�@.L�#�MLLT���*���"@o?@�ܻ�����V�����ϧ2�E��H�I��;��G}D����C�Њ����o�g�y�&�*I�*,rZ�	sI�ύt`�>��Ϟm��[o8YE! �SR	�*�׃��/y� v�2�`[�ƚ��$��(p�7?\�ɾ`���3-֝6y]��Zځ\c�8/������F�zJ��c0�N�,�{�z��2�Q�0�q���Tؓ�G:����Oܜ��k�8�@K����h/��bL�ē�[�me�0��}RJ`���-���sQѹ�Oݺ{*T�t^t5�T|zJRj��ʉ,sb?��T׽_綍(ܛ�j���L�kH���T*;�6S�l���#��[b$ ��I)0��ውR�?9(Kw�
B��T>�L���?�S v���k��I�TlbjF8P�4��v��14�����[v���+��k���8��R����P��_���h4�#i�9���IW�&�N�Ɗ"▛�"�<��HO.M�k�ԉG��I���=,�TD���n�Y�G&~��;񂗳��j�-~s��?���7�'���7��8�Y7P��h�,�K6�%�%��D�C��O`��L!��6��d���V��8����B��8��򪢰�b�i�i�L&N�u�$�a62#�`��N�i���7�G���]� ���؇\&0����_�ϱ�^������������}5kzΙ_g��� ���Wق�}U��f�.܋�p"�w��y��P�~ۦ�g}_g��n�����&�m���~��>L DK3�� m>0!��Gw�%�_sV3��u�P�l�ٟ��ͷ�x�,v�GV:�{"'櫞�T7Z���D���^T�'�Ɨ�V>�,�/��2AD���¬2�{�rPf��e���bn�j���F9Gic!�ɓ��o�ic��,g/KD��E��@�q��� �8ƾ�g�\-�Me��TV(���v�Ut�Cj�c�Q�H��O���'�V�*3#���+��W�:��Y������jX:�[��p}��e����\+L��vL�ǡ���-[c����@A��2؍0@$R{�">AҲ�Z��r�e���"��/b@���`���q3��骹@�e��w��2�����l���.�y2��S������A�,�m��ڗ�S���'e��Axl��C{��kim���~�ʪ帞���3C,v��S ���0��!I����:�����P� ���%1�n�͕D<�-�SZ�"߫f�����GQ[l+p�)|��~O�.���O:��i?�H��fP+���O~���2น�����+��[[#��2��F���'vgpJ�N��"���<|D��Y��(��5W|�6AC���!tSu�5|�+'<�����6H���tϨ������Y��?��:8�d���={e���� ����]H�W曈�! c�J~�mՌ�ԕ]l>�߸�#�	.��]!$��wǂ�"������@�iY��j��c]e�!�<<�u8~��~x�"Z
d�C�,�l��J�6T w��WrҜ �U.W�E�����:�x%E-���z��{��S��G�3�hN|:�g��Tk�:�)�♿w���Z��f	�$�S�N�qhW�v�Ŧ�͡��o��mx�.!Q���������8�
������{���w�Oj��'���T�9�B�����E�:��/�{g�i}�g�/��?m|�	�əŶ�����Gc5��˟7��k��=s��6�.���w�lK���V���C�(H���K~i2�������V�ϯ��zy�'o�jw���<�P�TP"[���u �;8�Z;�::T�G�[~Wyv����9�ف_�p	т�;����W�H��p%�G����Q���EPAZ��o�j�*�B�x��Iw*�z;%X���a���M�b^j ���S�E8��L�d��%ĊD�����sX���k𻀄��1<d�'��=3�A�#�z����j>k��{$)Fh+X3�_Ce��]��AM@z���<B�xKI�Xx�#"Kc��pޠ="���CWr7^f�r�&�\ ��;�z�IX�D�ajn�t��(��E��#z=�����w��Q���KX
���o)n���4˦����ꭻ��y��JV<E4ō���9l�-����TVN����>j�hH���{���A���Q�Ұ�Z�!��Ȑbj\v�ۚD�r�=���.3ŕ>~��Ȇ����+�}���bhc��(�7��Nu����F��yP����%��,��ІDE������D���L���P�U`�6Mc�UW�oZ��̢B/��i3�qX./Mx�Υ�ƶḌ���ڦɝ_T����i���g���$\�_��h|aڧ)�?�g��95��M�8�T����>B�Cj a�;~�)���}�Z��d���Q#�i�FmX�jZ�#@�����츖��R_Pz/�P�T@~�H�Ix�a�?��X$�Kj�Mg���ڵk�:15<a a9a t���w�QՉ�Sjg̏Tn =��֞vmM#�_�����_��`/aLL�\8���Ӄ`��@���9�Ņ����Ye�mO�l*�]x�'oQ��<��-4�ľ��ե���)7@#��/v��⒒z���h<����������k^Y��bM�5=VcE�&�֒o��"��N�`��?���H������m��2C|�n���Ë�\���̳iP��~-/�w9纕��<�f�.��OdP e�=�7���~��KSD[���1×�\c�r��f�;5�Q�V E���w�b�j%/�Q��/?}�O6p��_Ɇ4�gʑM����ƛ��,�ih�^�u���/�T�qP�=�fց�丸����:G~�Ƥ)/�%��e�4TϏKu^!�ѼKW-���<���2m��ψwL�)�������,�����=�V�$�E��΃�m;��Dw53���ܝa�CA��������wj����ȇ���	]QZO �������3#_�N��w��7�a�z]����	�ࠠ��ϟ?����	��)��j���$��U-��AmJ|���m�G��,�p�#kr�����ˁ%ʝ���lA�+$;ʡJ�*�����ǟQ1O�Y��L�؍�5�9^>"�H����0�\t讃miǿ}V��g	!l%-���5-��[@v�������*���g)���,1�(��i�d =�(�{v���DJ,��A��׹���Px�gڨԏ���{�[����h�]�俈��~c�ɩ����="ԟrb�%���QH�����V�z ��c&g���FFF}!@Ӵ�],�w�"�]R�y�L�a�;�p�'�Hq�����Ι��k�����&挱z�S��� n3 0�G�	�0Y��6�DćPb�O˼��N��ߖ��u��	"|����s��O?�	r���<=>~	S
�C� �� �XA��"q�B-�HR��΀��چ���
���}%wOE�ӟ�L�j?�1��[4;��2P�kl�ŀ�HP��G�̙`�DSvPÂ�h�Tא�=�I	Xnj��{y|D�'yflW�8Zs��R�.HA�|�yN+(e6��h*���(��d]c��]j������� �'���S}e5CB��S�� g��eM�w��A�i	cM�_���3wB�5����:D����Y뫕[�KJl/qo_f�[lK��̜�An�|�in�(�Q~�c��f9m������O�+�G�Z	o"c��"�[�tPkY�L�U}f�4	,���:˒�Yb�OXp�<$k���2�;}Q�>@�PjR���}[��~^r��Y~�΃�Nv)��'���~��{���u�3���8�0�h�2�oÚ<2_zؤ�Oi�����SuV޺;��5�;����3��e�+�>�5��3�.:Z�t��%���Dqgg���Ҏ��j9���,~�^ ZDI%�37�|�_��|L ]s��Q}$�}I��U�O�7)�݈��p3�����A�wD$T����`���T*綽gFvF��|�DFKK�Bb툟 �KmA���`�,>+̓�/ׁc-���C��^��w����?M�^���0�Ը!��[P��[����ڹ;�S�yi�I�8��;��� [��CPF�u[��������aP.-S}���4fnz�5��K��]��s�������f���ڐX��u�/Fk�@qBz
�]�`lV�n�m�:�[f(��ù�����\���]0��~^�37"
�@���ן�΀U2�⮫u%@�^ P���'1hEl��o�%�$�6T��YBQ{*�Ea�Y�������{ a���npj�	��넷�/5��)�[�z�$J�}�lQ��L!�}���ߨu��J63ǢZ��g6{�^�i���~'��N�:�]����'���o�U`�{���l�����qcO�>�݀.�e/N}�+�¹B@���6�?J�T7��y�* ��\hY
�Ö~�E�#��1L,������2*� 2�d������@�07Hf-KҜ��Bم��f�T��^�� ��|���i�����l\dkɭ��p�'�Z%@�m"��|�`�?������h@\PAr�@kX'�򧥋��*LrZ��If���8���J��L.���I�S��Y7����#:?�:�ɬ[�4�&/	^9j��S�8�L�`�A<���eI�� T��C��ޔ�����<�}]ϼ�ނ��m+ùw�7��S�X���a�(���b�[a�N���h������i��H��"�� �ςh��
�a��������5�@,Ő��ݥ����Rw#ŏ�1cu�|%��ږ��'|��H>���л`�X������MP��5~ĝ�q���[A�*��	8�6xA:5���������u�����o�:{�K�ڊ�m7�\j�]��!�]%���P2��Kr�M��"�M�vkQ4(M���&]�&+CaL��eH	�眷�����k��s��<���������Ґ��K��M�$��Aw���i{b����`��@-���q$�kq�e!�b���6��4���t�������_�ΗFVg"6S�װ~Ov�hY��?�a/@�|���LFM!$³�#��˿#����332���o� $ j�L�{�!�z��"S3H�T�K_.L�
�vg��;V�Ul�{�\Cgv��!�z$��Xŷ���⮐�v�+V�&�v���u��V�V�N�{r~� �x
hPKR4cC���Ɉz
������Q'�G��J_+4A�\V�e�ҹ��D;w������OY����@jF�~aKw���
�X�R?/T�XH3�5���L$�#�(R�=�.q�?
P�_�&�2�a]Q��(RH�03�~V�{��6����� 矠����I��|�X��Xо��d&/��lc���ެ'LG�%��z�y�����W[�S�rj�{F|�o�W7|��jii�-�;��G�9�@Y^R��yx���Cg�f�#��:O3��kb��H�m�`Ψ����u�1��9���(��npKV�+c`��I�*�\.ٓ'���[����S��D���H��#`:=6?ڕ��d���.6����H�$�4<�m���7�t�,��W-7�����TA�7��i%e���[�6Az�J�V�t|F�	-:��R0�$�(�&S�*�B5p�5��[x� %��|�C�K���z%s�
��0{RZW���Y���k�S��@�y�͠��!�'�%�b���}�m׸���߂k��sZ	�
�~�ȓR���G�TQ�x�/n��,YJ����;�DZ�h}}����:�t�U��ji��_��%xÆ�����hZ�B�mj�]�h�U��r�^䠘��2z��|����Ѫ�����j�d_�n����WK�}�����'a*��E	��9���VVU���}�#(nK��"5�`Ah�U��o���1/�������"�I��}�T��8A�%�ۨ���|e���%��oq6��|l%��+ӆ��ž|�޺�њ'L�F��7���S��[X)GӤ��ܲ;��:���m�L�t?b"l����7MWԉu�0��}���gtRx��ѵ=+Ge���po
Z�D }w5���q����� [:����?��#t�755��:U��->���t���1���dYXm�D����|�� ֢��nk4�@�8��Ldk���N���V��N�����:��H��=NdU
{�A� �Lu�|ŋ��������>�>��Q��.1����;�z�Dښځ��+����+#��y�5��<0߰�H�ڹ�xT���ka�ͧ=�rU-C�1��.���]Ƙ����#��sd� ����<JC)���v��5��c,�f������S�tDai���?dS+��-�'����ԉ�R��r�e�"4*�����G7�� st�o�#4�揦��U�]�wS���(�ܻ� VTGQ�ea��OeБ��?���`�Q��8Zc3�{\��1p�_�U�)�	Y�*���:F��}��)���IB��Y�����ƶ�����@*�Q��W���Z�T�_�xa:���g�)���mu+�%��@�;A�c�͆�;xo���b���c|��96
�(m
la��2ާ���)�@�S�������Ĝ�5-�ãr;�ܟ?8��2����^a@�ru~s��0;���ի��H��L�	�'@����&�FcZ*�詶	].���,Sr�:k�>���s�S�`z';�Wbb":�YA� 2�����ʗ(qgqF�́E�h�N69�ri��P93���[�/��BW�@L:�Zj_�^E��o�X�ʅ���V#�Ɠ�y�+E�A�Z��c��^o�=߰��XA`vbD=��%0�:%�S_���gl�]� \W�ŕ��J]�ڶlҦv���u��C���ZrBT��=w�0����۫]�\H����#,���GO.(1�����C�	iM1�jM���9��9�w_\���a0��Ӗ��Hti�.v4�b������#b�I����>wa�貈��w����[Fi��OO:�wQ(-�����.�*�p[�fϘ�?B�4-�]�-#��a��s^��dGVEch�>�
(���W@�q�L���]!a;x�P捊3Q���x��&sK-�Xl>g>5���p[�ߪ�Ӡ���ʋN���TQַ�0�3\�o^6�Y��YI�#DQQ�#A�ԁ�(3�zmkFq1`,i	 ���%9�F~q[��Őa�����Y �� �y��ǧ�b@Υ�;ܣ������Z�����7�0H��iK�OP�Z�	2Qr�in��~(�w��k���K�09re��f���.9�$d���H��ɱ�'Ն~w�y�V��.H'�Y	�G!�wzݗ?��5���������T��/%W�S��TPi6��'�T'���F��݅���#�	�_Q�ָ�xi��Ps�W��h@�)�{h�whm���zuJ���ܬ�0�]^c��9�o��]?��i�~� %3 ����v�2��I>Ƹgl鷪��g��(VL�Ku�_��Ϯ�M��T�zFa�
Q��hP ����ɗ��g3���mlfڰ��W3�!����c�gT��H���Ooo�x��AȾc���b-��7.H+O.v,���N��㪻h0�ka�Ç�>�����y�FUP���u���В;�!�N�.�
�T:���	����8�u@E��db�¸XWGgj@��N�U����;)e:�u�8��oe�wW,;u���Ө1���
�)��0���7���%�";J��,�,�6���
�x�A&C1�n�I/�0?�mGt�:d�a���V酉���]�[M��Y���y�>�)c����s?��F�+��V49��a���w$V�j�Z���5\�jv�Ü��
i���hٟ��i����<��^�����s���J��]�l����tE���{��)�eG��i����1��`��I��(��Wv���>��Z�v
�HA�Œ�hS��Aȧ���4`e���;_��_Z3S�C�d�Ξ��m������0�.�����#�f(|{M ��T�Z�Q��{�/uȌ��I�!uy)쀬�B�|G^�9�E�r��!�!����N�� =�v��=� k=��f1 ~�*��5ioksKv��GH������|N^ԙ�Ǌ�`X�� Ai�O]d2~t���4$8�%ga��v��i�R	J-�+���q�s���"���u�u2��C��Q~�GC��5J ^�tF�3�W�VF{P
�3.:%�=_p�g�bj�6r�ܬ$�pN��F��B}r�>)��?L�n�Q� ��p|"=�2���E� ��Q6�	ɳ��M��|��o!�*���Ѥk��9���qJ�iK�!����ʼJ�	e�癛��u�$�P<��������
jg�Ƀm�q�hcƨ-�tHS�l�?��5$��\ȱZ����gؼp�"�oԓ�_����(���j-[��°'Q�[h⭡�u���@�҅(�/�̤��$�ѐ�8��j�������Hh�Ը��%��:c�Y��|p]ѳ"4��t�/9�Ȳ�L~U�`l?�§M=ى���=.�nɊ�x�~~S�A�)��	)�L��3���^�i_�ZO��wl����!%�n��=��x��fy쾵K=6�C�J�C���_2�h��p�Tx@.(���G�V�{���9}�m=�!���7vAN��	�"]�4���C/�-��VF-v�]���o���YD����|ބ_P��]��/}�=#���9�:�� Z�h	*�ĕ\�$�Y�zH ��։/8=�H�a#2쾆HV'����u�胶g]���̍�xI�!z��Kڻ�uB�q���h|>��"���<2T����a>-��.�?��=��S��T^�ۇ����]j�w���ť�(�Ԯ�3sD��S�>�x�F�.��h{g��f^r@!\^vgp�'�0U^��și1���j���nI�*�߮�1�к:G�'�3��cB��N\i�`
ŭ=����P��!���pg[ ���N�@�\.��h9DGSn�M,%����D\;�
'&r�/�x���L���^ȕ#��^ˈ�O�kz���\�d�P�_�pT)^[�
Uz��'�D!����Ј����9ROV��ݢ���~��{ٟ��آ*p�xϩ ��c
3�/�4�A*��wAk4�W,=�����<�!��`2J*��!�@�b�
�Ə?/e3�! ��Ͷn3���[WS�<!>�0E�2#�!-XH��~tD�
���mޢ��f��O�v�l��<�d�i#�jM�	e�X�rL�#�X ih-q�;C��6��m9
�S���״T�y�:���βu��%��W�c�����`F"˸���c4z&:vƧ��m/�\������i�Q��o?s�_Q�P���V�9g����eG��/���r���{/揭��w�Y�l�9NM2g��ymǘ�[c#�ё7�oDG�X]�H�"��s�Y�	���T���Dev�q��Ϛ�Ɣ�
2���I H�����X]�`��rp9��?�)[���"u�R������v��R�_�"M K6&|�{]�Q�Ԁ�iP���d3�����
Ъ���G�:ѲL��i���v΀���c\�8@�@�������S흒�-���M��}�h�@�P��Lsǉ��@�Ƨ/�l�M���	�hj�ܹ���:vfW��{A���c���'��T�Q6��*��@x��������=��>Q)jDc9Ʒ�[-���x�c�S\�k]T��>���$.��(Z�q���s4-Ɔ���Y�r���x B�%r��!�S:�?k�
��-0�c�O�&����� ���O����&Hy%.��,:m��J�xCW���x�០}in8ȃ��	��@�$@�՛���[�����:&���;D�?�n��P�� �k{0 �|;Ϭ�q٧�0.0���='��?�w\O~��;�@d��6�Rd���!���lH!�m��9n�Ĕ�%_�qH$2�ᇆ�<�L����m����G�\�(�9m.�Ml<rRMt�˽��{����8�Kjg�4�vB�µ��9��Z��g��w�ƕ-G��)�v�A]WQ<�6R#8B��]=u̓�G@����e=C7�/3� �ė�s����
��9!;�K73sQ�h���f��s���8K�Z��ݻw�8T 7_�6	�ѐAâ���w�!{5��z�	�n��2Ch��.`�0DY�ה����HS�j�-`���8�ܲI ����������xT�J��54,���[���HcI�Sr�A�+_���-�	iXK�ڠ�a?�گͩx�8����m�u�k�g֎���c�w�d�-g�e�w+�	ly������
׼ ��A���A�"IJ��;��>QU��2q��qS���J�u�@�|��D^�F0��f��HuJ����>s���9'Ba~zq�������"�3�b�e;x&!%lk���\��ۏ���YZ'�����7 `��(����w�wG���6�]�#4y����-���_УV�U���p+L��@D�1��d��tWs"���JU�.�l�����h���ϟ:}����-8ܒ:g'�����$ݜ8�興w8S	CW�f�FL�r7z�&����晗OX�sb�o_�ۮRy���� �	�pEEeeT/iMtS�+�q�����c|}�sU��m�����(H�\�[��M�]d�5����b�5�]����+Z.w<�S�M�2�(�*N�1�����h��P'��������M��ȑD��E{
m(�#�o���i^'狎��ks|��h��|hrmC{���o�������I����nx	���ݹ�v%��ճj��{��o���&����3K��x�R��0/��qe:��v�PD��A�|8��{�ft3���lr�щ��!n��J�w)}}}J�nJ��}�R�9��#�@�{p�]n��T��5ϛMB*~�M�|��ZY���u/��߲�_�Z�^sIh��JeC���o� v �pM���5�
�c����z'��~ym�׋�+�@@��/CG�b³U�%b7w0���C���\�)Е�|��&��k�e�*�m-xx�]ځ����3�n����t� �u��K�*����� �}��o� �¾��\Y�yK|	�z+��z����r���=8��j��N m]c����R��V���d���'p�s	2���6��H��9_����Ge%�&1��k����P*T´G ����vn��n�9��;���?@�Z��ܪ���T�Ӯɣ�d�(`9O�J�X��W��9�rǪN=r���Y70�5�+Zx�O/mN[���#��.����8�v��}ϵ)ٷVf�Ǡ�s}�H��f��F��a�@�Id��Ӡ�����G����C���D�U���Є�B�D@!��QX.}�Б�¶Z�m~PK�W���B����d����'�0`��T��w��\"�������&�y#�i2�������c�*�Y8*s�V��㕿�jRl̳$�����D��S�SU�Gk��)�.�ۄJ���`�9����zA��G8��� �G&�$b��9�w#�r�׏ʚI���9zB���:Z��2��~L`�(�D�>�Ԫ��_/K#@^i�"�#��
�&��6��{�	*���H=��I��R�kbЍ�y�)�84򏟻m�⅄�ap꪿�,"�/��M�-��
��O��� �*H���0 J��:�7@�"rr����7�/pOv:�
m`&�&�c�pa�I��mG��x���ԉ�p���
���5_֮��t��9�� I��6��7o>�@p�NM���`�zd<�߶@�T{\Z���XHP�%��u�7�]�9ҟWƝ��Z_�,y�ie�\]�}���m!zPe=�/������m�W�����t�-:a�G^���0{;�5��W��1˂^tޟq_���wlA��{#�F[V�ҹ-N)dGF*Ȩ(L���}^�	�����3���W`bj@+6�^��,�xx�S�x�;��l�:�v�L��@�Z�dǧg�>�T��_�í�tw��?3�GD�*�,p^|\U~^ }��h5���	z�PR����ɳ��d�+�.	3��{��A$�-t)�_;H ��h)����*������ԍ�?G���;hai�0��*O�L��\n�0v��۷�x� ��˹rg�s��/�ޭ��+��A���)����`�t%H�怪�o�oF���G�Ңg�$%%UӨ������U��x�%;�P�}ݱ��'��9�y7�6D�n@U�A��>(��uߤ�/
S�WF2|��?}���l�����Հ�7K72��(��w��Bt�/���8�a�ϴ�W<��Q����n��� ٢�S� z�%�ː*
�������?����6���\r�V5u��A!��� :��PR����G��X)k���tM=�I�$'�c�yИ��]�KB��|�]��5B��m�m��*���5�b�m�|��Æ��+ڍG,h��M���r�O��RY�Zh�M�@��,��G����~'��a�F��Ի������
GB�jEq�#��*-�T��Wo�l�2c)��ro��g��|ǚ����W$�����J��9Bc�E��ָ �X�X�x�Ω����TV�~hM��MN����'�B<�Ğ���I�%��"�d���|A�C{kO@,�T�3PYJ�ڷ'/`0�	�w��M��-�׿#��Pt9i"w|g�����}��H/b�g�i��]E��!��z�W��Ya9�5�{�e�.vqaT��`ٳީ�b��y	�y3���;8�C[�}̩���@�[�vP�]*�)Rf�a���RnM7c�����k`�Gt����e��h�L4�["�z��'��n�; [UlE��q:{AL����>�B彶���Lmk|��ym�ď迊�7���������e�!��=`?1֠�� m��$;��BZ�h�g7�����ĭ�EAe�n���+���
&�y��իj|��(	��b�5��B{�g^�i�n�(���smD�qvno|����KC*�M�gcc�6~�4��I}ڌ���KlP&d�1C��
��;�/����4�-�U�t�t�Kp��:�%��zs�b"�w�`6����_P'}v�w��ڠ=#j(�)N�&�S8�����*�C;���r�پI℣i��'��h��:��.��i��˞�Z�3+����>��==
�R�F��O}���E��ND�*Zڠ}5��-�ͧ@s<�%�U�E&{ OBHѽc|MJ�I�i��m|:=C�<8v^��P2���m�o��n�mv��&�<����,Օ��סʃH�!R���~+F��{�^�Յ�i��
�D2S��N�A�7���xx��;�m^��'��d't�BєqPS��:�3 �s$���1^�j<�Q�	3����E��+�D�bҩ��Ԧ��\;}����M ��'��?���v5U{^�W�`pd��/�ŏ��n4YgŢX�xV��%��h��채2sy��g�>���7�N�S��=�ro_��k��4�v9yO�uvr
������9o�:#3�*IM����9�]�C���C~rwt9�d�'�钠��Y�K7�_f)L~����ۤ���w�Bͮ9Ƕ��Q��	z��c�OU\�yU}{,K��5C�v�������i��ڑW�%;gƮ�H_�q�Gqh5��ؓ��p1'u�C�~�^MLT��!�+?T,o��?v�����5���C�e4�e��=3#?��=��6Xix6/[;g�WH�$R&ZSߏN�D��+^��;�3���u���e�'���`&�m���oB5Qh�D�jr[�����'��W\���&��h��m�5�wzx�c�^��F~MӘqzk�z�9�,~ґg���G�9|_c�[Ԡ��+D+O�D~��[6+�qS��M��FJ��X�؍�C�YrK�#T�UL�
�M�u��΁��hC�Nۈ�����3�@H�������wɜ�,�[���a��M�b<�܀�H��p��o������({�+��B������mbpk}���!��$�GE�2Ԉ�,~��k�E�Sd��W###6x{UQbf~~>��u~1/U#��0 ������r��o2!X
!R�z���	���j��?��C8���*��0s�M]4�;�/�BU�2��ߠ���)e���S�y<���Dj��L�g�Q9�ӟQ��vi�q�*O{W�>�`*r���q�I���u6�Zę*��u��z�ם9/9�4�l�E+�)/<i�{&6����������(g�����-�6� T�5=8j��D ]����{i���f��Gb[�����c��I��	��SOC46�D�i,4*j�Z���^�������Hk��L(��"��ڔ^�	�ƺ;���m�M��������R�q8ףm��N0Ζ����@�L���\�xAV�j��*>�r���/SX	Uo�8�$\��@f�q�oB�t1�K�s":z�J��}�R/K�{�RU6쐈/.iS!�?U��pD�T��XV׻����F�(�R��O�|{�r�����n,i__��jT
_�}�hZ�A�&�Pg3��V�
!x���ՉCFRw����<}��̖\�1�����8�/f���<���)�D.�X�R!2�aɭ-@ޫ�nd�����JT$1t�^�l]�]$�C�
Z�LN`wB;��2;Y�޺� }�P���d��j}$ґs@�{fW��T�N{��S	��� �S_��+i�js�!�M����*��m���޳��dj6$�np�;=,�<���}7�@W9�vĩJ�罄�1�{���7���&x�yԘ�7*꽺�?�4~��W���B��$���7o�,����@��|��[��c�g��~�~CK�v��l�w�j(G�$LWzvr#���)���E��x�MH��n��zC�4���G�iي^ǂd��O��d7�j��"�e���h�f��j�B�m��!�K�U��;#�#a'�j�*�0��ȯ��׳��(I�p��mM����lՂ������0_0�t��PZN�8�a%�_�
r���j�8�7�?緜WKpy���S�"�If���i���S�S�ހx6R*�;<��5U�z��tq������h]�)I��9�Ӱ]8�e�e�M��M��eO�^A��>�:�[=+�d<Zop�p�P������SN��.>�M�������*qA]t{�ɹ�$���:�N@د�`���{K��#ϲ�t�s^�F���%}Gu'{�X@'��c�{dV��'h�cd�&Fٳ�%�I������L��gBKZ�����ai؟�}�+;�?��dz_�Y+�j�[H��M`��\�S�U���vѩ�H�c�)��k�A{��h��S�C��z�Z���hf�T	␭�`u�$�D��ˡ�m�hL����-�����W���[kP^��(�����=�����v{�/Q�����yhM[ܭ2�S�zw�y^x{��vT���ÞR^�TG�3�'}w�a1��>: �N�f��s8S3���NɵlAG�(�f�C���HxZ�2R��ц�����;:H߭�E_9�{X��H���Po�GE.�����#(�"�^���ŶO�z��/��9���u�.�Y��yV0��bj5m�4y�n��&9�����;WT囷�D�7��B1�����s���k�Ӕ�"Ϥ��uʋNU��k� ��1����;3���D<�`:�[�7K������C�E������	��6���W���;j"�1��Jp��
�UT��!4)|��?����_��D��D��ֲ�7�fe>oL�Voϓ����GiJ�=nCv��y��ф���Ԩ��W,=;�������EM
�{s����S� RG�{U�{RU����U�V����I؛��w����N�� '��;�x��3�v-�C6�ɕd>#�s�lL�''`.�]����t���w�q��E���Y���b�m#<��֭R��Y�o�l�q<.�]4�o��w��Cќ�������I Kk�ǃ����qܣDZp����n�ᚭ[�ą��m����n�C_塟�ۑdі.��*��dv�6�r��c�j�rt_�z���W�}�2dꡫ�=Ws�Jp�BWd�Ѥ.��3�ɔ[^ ����h��mnX�K� ����D�
W6��es�:�yz��k]n!�� �q�N�<�0�i��8T�ǘ�'r��@1	q�a������3RhFVS���s��׸��n��=�����2�C�(]����mZ��~�c�A#z�vptt�#*���߇��m4�_�QS&誦� ��-�p*�#�˟��K�kh^i9d���r?B8=*6����$9�յ�z ��&�I����Օ��˱#�<�I��O�k
���rձ��;��Ӟ�)�NY����C����K(����ڠ�Gb�ϑq�U��8|0à=�R�,���=�!�Y�M�XtJ(�h�X���h�^�$ONJϥ�c?�����<��O,�є���`[��?�<��� F�vl�&4E��p�y���Э�-2����%��k�L��"�ſ?�-ɜ�&r�?���M8��M�A�n$���7ԧ�:��z[vS;�\Y����׬^
=P@���,�>��L�X&�_�Z��Tu���W�3��}2Õ="7��]jzX�v�	M�(|o�O,
x>��L���aƔ�H���
�ė�\�;��W9���O�]��Cl�=�5�� ����}l:�+]]]	~� WW�%�3\�AS�"B����݆x4��=�#��0������%}�G4�����C��
���&'������o�OԱ���h���r#�U�@>��h�����(�y��� k�^a� ]�ӟ�~��˰����Q�^!�����0@ލ<��o0v��$���4
f�0���d����fM}��8��n,�)�ŧU���� lt��y�3~�頀7��9i�c?�2����Bȴ�7�H�#eO!��"��"IZѠ�2�_�&W���7o���3��x&4���Hcdu���� ��G�߿OV:u��!R�!�bChd�Oi��|��	lL�#?�XuMP�O؂��|>o���=�s~�%x�+'u)�:�$l�o4{xxT�`����{����24�w8���|�K�2�G?;��	8���nN�������^�|AHӿ|���l"jz�K��"��W��@����O�ɜ"����Y{m9�3J��&9~x�"SD�h���1~1��2��4�����U_H=�$��/���/��3j*�3��*7��4�J�.�|/��K��.��7<���z���~RuU����K�v0ޢbִ'i9�rf��g�.����A������m�8�=�(�!y�!���hᎼ��=fs@�*;��.�U��fS��~y(&�<N�I�ܴՓ8�>�f�Rb�%hn!n�A4�wE�&z lEcĸ��w���@��H��`a��W�n��0�C�$	��5�~��C�'�ji�}�v�xIa
)�'ZvgDՁ�&w��B����æv�x ʝ�٢�c��6�O8vN�b�0��A>���|��3�",��mE+�UO}{�J��Ҥ(���{<��@9rR��L)Z��q�L�H\�����*l�_`�V̵K�+m�f�e���h����ÌM��J�GR�w}��\ׁ4��1��W��C1D�pV>���p��=��:���T��(N�5"�D�}��Xxl3�4��ox��j'{��?��ag�����sT�����n7{����k�M0-J9*���l^Z��_��}�˗�'o�%J�Ю(��cSI���
��6�h� ]��{ܗ�&�~|���:��;ft�9Ry���/�5J�E������VM|�$v���S��@1f'BW���T�k�G��͞���K�P�� �Z$B����ۣ^	��uD�sKT��}����t��DS\��t��8�2�W�&�2&|����9�|�:{�Z\O�LLJ�1G�Q�s�\���G��'�j!n�(Q�,�$�<#�y��E�B�RW�DH���>.;L� �p0+x���\-D¹Â���9��b���6u-�#l�Q;q�����G㶚�Ł`�'2jԶ��
��,H�T�9��/\r�dEL~U,�R��Aѡ�7��%r8��u��D�&�-���ы��#� ��t�3�d�%��{��a�Uh�(��8A.7i��v�)xޫ�7@бԈP�lo����8h)E�%�mW�g�+;��th�x�]-J���Uj9{T����P�q����/t����t3����&vj]7y+_�=0�R�s~	h ?�؛܀KQ���G�Ll��|������/�.�{I�@�ܳy��uاȀ؀�6��}�ҵ�����
H�(n���{�����ע&��j\�j����$�~��|}�=�rp!��@OS�p�@���2̅:�e%���%��B�������nD�k�,=]@���}�i=L��-���� �;�����wH�����Fo�t�736�ʱ/��MLG�.�=��r���s�(�߼qꔑWK�l_�f4cn�#�e���k�����h�ɗ�t�w�5%xFxM����j�����&Z!��AX�tA�`˛�1q���^�X9�/��i��U���Ǎi���3�/$�6Z&�<#+k�Ͳ�ծ���=:�6���+h����;>�v�L�!�S����Κ�(wlr�z����E�G���{�ծ�y+;0A���g��><��&	�(���H/��J�F�$#Q�&cպ�Ca���1�:�2}���>��V��o�n�=u��O�6} ���>>>3�����f�,�`���"�B;�;~^�J��M$-~�~w���=�����9��\����Y�}!����8s�%�h����q}����(�6XM�mMie%�n{����r�M�щX^a�(�6L�n0�/}D�!�)���8e�Gn��#	�l�{\%Ϗ�� s}�j?�m$U�t��c�ܩ_ �^�L��y(�p}l���nz�R�iU����HK��ڋ�C9Ż�0��E�q���Τ�%�h}~���Y�:0֊���X5l.F�G� �s���=1	����91�L������44��D{��'T����Z��^���`<JQ�+a�!��Ρ#�L�`���d�]$��&G�<%	��FMM���Ĩ���l D�75���nBkt�:B��'����0�>�;ohhz�'x��d鯩=F�����]g�K5�x�^�ul�ϣi�9�*Љ���W�Z�ć7���nu(fب����W��X�l�����P���}g��.y�\�Җ�C��zn�T��ccc����2�|T;4���C_��'CB�νV��3T*������|�����=f������jK��B��hZ�n�ki�.�ѡ�mgFބ��T���LӦ��)��_��s��r�n�ЀΡ��C멝zy�=��Ao�����lg��N]F�g������R[�[�:�?-/<��{`��i9�R1��A�<������0I���V\�:i�R��T�"F����g�'x��6�g��o������ڗs3#^{  p��+/�h�8>�h��a֞Pb�.Ȫ3Ҟ�X�q��-~�"{;x�L����[F��kuN�^��Z�M8�fה�OB&�������t��z�:_r���_�����3���S����
Y��;M:EK)����S�Mm�^;�~[���.�nE�0T��0��mO���ݘ�b��.��/�%䦣2���w0b��������?�o��H�K�jy%K�Τ�k�'ԳF��`D`��g"��B)3��ee�34����jMiv��W7����h�(�PZN,�ptd2)�(�+�nv���X����=Z�߱v�
pf&8�qP��o#F��$6�Y]�Z��}��}��I[��+��xn)��hC��9e��kߧ��U�0�t_;��f���h9x\�k\��|Q�>}�Pp�f<rF���.BQP�J�\��d���Ka�]-J% ��T��2يk@�\�,2��Q�_������A1��g��D)�*�yC��/�	i�wV�$��4g��p���ݟր뉶 �𧦕ձ�U;!HR�]L	Y���}m������3-�����wO<��n�i��jW՚����}�
���$kDQ��^�J�<J����K[ƣ��z�u2!�w�q*f��߇��KZ��Q�P�	�ড়P1� OF�L�u�NL�}�����Ʋ�5��Q*�~�dz^�f�q�{F�<�3�[����B ��r�C#r5�o�^	�g����!�dx��-��PL݅�>}4�x z|��M~�X�$Z��� D���b3xHZ<^���ŜߝX�LvP0�ۢ�у����|��v�s] >-�P�Nk�5g�­kK�����~�#}X��q�ͮ��>��[�%g3�4=������{���5Ԙ.���
��������Z�:�,�O@��q�'��ح�y��I�:Ѓ�z�.2�l6�����I��[d�-��&� ��j��Z]1��Sy�p�ƕ�;a�[�q�ѤL������<�5��~ק�GM�8mn���_�l&��-����_H /�����L�����k�)ʘ�߫���z�SyWHT���q�C��X&q�}��uk��J��ϕ�~K�A�PL-��lWd^ý]on��8�T.��~d���1�(�(d�S�&Ɋz��c/��W�<틈aQס7� �-F��m	$�͗R��$>���Ӓz�^��K�xe��W�W9��_S��Y�`��3��|���㹖ȖD�� Gt���QV�: ���R�P���=��:��)
}�<����ѡ�o�_k'&&lJ����i<k=�n%�D�6��l�Y5����+���s�BA2:��z��W���Y���*.�utC_f�?��
�~�)��P%�K���pV����=��"'�EVw�x�v��}j� �Gvy�t�o[c���,���Tn�⢀&U��Z]Q�rސBV��W�,���)ˀ!�c��2���01��'�($�I^�����R)A��@*\َ{CE����7 �+�{�7ܕ�(+~>�jG�υ�'<Xum�f+PE�-���^�΄쟸A�p��3Q/��}�������S^��Ρ���ה��k�Z��0�Ïo�Ү��s
_�����*B��Z�4���3�,.Љ�,��%��o���������sI�̔Bg�*̤��yڷ��U��� >�*Z\a\3k�?����V硿�oE�������M8���K�^��#�¥�]��v�`�:���m��Ya��휣�b�R^�i]wD���Y(-1��h"d�{m����5k�U�������Hw"'��7�`<��z������D�O������~>.����#�ﴞ�_�'�����!���F`۬�]1*�)(WIY-+B��2�rL/� ��c>�N�`��&��e\b!	�����ߥ�6�(�l\�v�tq��/���5���xe�*j��)�����p�^���Hs@L-ߐd��C�����
k�'m��]�[Y�^0VO�e@ *]~ ��5���"�	���)��j���Z-Pve$r��"c��Q��v����ޑg���)c~���p��|z�H��Y>|V�K>>nG�v�t�P��Q�T^�2�۶����
�1�/T C���f,��b�� Ib�Cq�Q�7��^�,�K��Z����if� 竳�FqX��S�*Z�,����c����҆<xSO�p>,grz���w?(܀H�
e�����[��|�["${����!r�Άƀv�be�W �-���������3gu$��/�j1`u��q��?����bE2�P� �f���Id��B):��N ����+�}�
k�6��f����v5>�靁H��@˫�9�P	���(�XB�Z!���[�jXJ<�]��`�Ѡ)�v���l,F��I�)��| ��@W�1j>c~���ys'��i��'�M6�9����?!0�C$�8E���D�(��a]X ;p���"�3�__m��`��3.]zO��£iJ#�^�C����΋��=�[���AyX��?+Zě��74��*���4�:�[G%�s�y���M��|��(�m�j�� aԞ=�4�0���r;�3��<��X�`TZ������L��m��@�{5Z^���Rؗ)�ԏ�l�ދgO�O�t��lE�y=��U2;y)�4���^5.^�%��,�G'&� �ٯ�Y8�s���/{�E(lp, �������F�뽇{
ʱ�s�㹅{�+�S�ˆ$��B(0����]�����|wr��,��~�v�=�'A���y�,���}����0�n�|�u��+�D�u���çQ*g!�Af?"}���)E8!$�W#����e;�T<ic���>�O+�N�uEX��F@��\�Z�E�4�ߌp���!��ЏӦ����9AO����(����8����/ �&������Kjg~�(�Mgo��R&�WҰ^��^m���S`�:�f�{|:ς@�-�{�.�D`�?�� �mF�������aB	z����Y1[��lG%�r�D��Z��0�@��:�[���[���M���:B��\n�7�l�N�i�}4���3�H��!��������߀�tm/�k|��Њv3䡜>/x���|U��A!f#��ku]��jas�F���������0Y�9�xZӁ���-�q_Ѫݑ��適>�ղ���l�#����O᎟d=��O=����i����y��B�>�ĪO��?�������<Uσ;�T	ݻ�+fg����mL4�@4��I���L� �3�d���
���2�#g���?a�Ⱦ_e�9���V�54��Q;yG��/j"�H�ajg+�՗�@�C�k�V�nuZ�f���_0����f7��4S�E��$�1q��e,��#�1�r�n�S]VV������I��`��O�Eu�:j�%�F.<�C}x�Զ���	s�r�5�oA����Q\�%��6Bh���wA-��l��� �8!�g$	�&��d�����X+�+����>S�xd@���\E~�Q������̡�#9R��}��������}�F?�NϞ	_�6�|EtȻG����[*fȸ�Z��J�l�+1�:-	��u��0�gB�hFT�@���kh��1{��Ay�7�(�'��Jz�������ձvLL�`�xTr�#}��|oMħ�zy�3Hu�O[�@SH=n��rq�E��m���Z^�2L�O��i8���zm��~M��Ѧk�D�/\��"���ˊ�A\��'��:��P�l
s�� '�^�n@�\9�>y�=p�+c�����r�cͼ���>b�Cp�mA�?���W��B"�J���>�5�p	����ȿR||��_��5�]�Fs��hÉ���A�!�RY�l����N���7	Mm2.������|��0K^��Ð`>�1.� �.�~�a�Zi�-��2���x{mJn�*�束�O��H_l� ���'A���E�v0���3W@�נ�׃!<t.�垺{b��ub.�W����ne��&�A��K	�9ϐi�$_U�C��c�� |2�\���Q�H�0�g�ΚC�J i5�DW���#�q�xᳲ�� ���zv=>Nh��c��ߕ�����j�4?�������-i-�I����d.�����Tc�dVa�w1~�=�9�:8��1=vM�l���(��x��1kroHA��p�#��mt��F�g���U�w	Ew�Yn�U�!����>j'h��r='롸N��mvlI�����k���:���Qu�å����d���{޶I����s��'�����S{����F?瞅���S�(=�bTV��.]A=I��n����YzV����|���2n�:�ѼQ�Y�&�#{UR*H�S�q������U<���-��@��-{ݬ"���v>y��fX(np��<���W�N�ko�CWK+-�E7F�H�ӂP�����+�[X1Ÿ��kd%�����SΨ��d�#WO~(��EΝ�?Z�oٌp�t�T#8�`3{�0�J�����d`Hq![=�<��r�!�+��W]�)eS-��;z�<��,TҼ,~���Ktg ��ڳ�o�+��J�Y]]��`�v?��*@��pU����ޟ�S�����4h$�Q�J%
E�ШdHi3��%)�$TN���쎐�:Bbۆb2O��Y�Y�:�߿���^�w��~����p߯�u��{����%��K�o��}ς���PͅKKP߇�b�XC�Jh,�J��a'M�S)��k7���J:�|�f&�O[��h����
�Do`E�%�Ⱥr"���y�u�ڮ�i�L���řV\K��H�E�dIC��4�1ִrW�Ps����9aM����{%�Y�]D��ޕMu�jY�[q�Խ ��]�;�m)�F��!�/�
��j#q#ٺ���Q��y�vXta��)���f]&#���É`�8�M__!�.ӌlxB�'o���\�ՖEtdІ5��N��ʝ�'���=�],v�tw���Hl�K*��t�ZD9���t�0�#(ԓ���ͦ�1��H�:� T��t���:���,OgJ�h�#�1��V%ئ�
�]+H!3/�������Gtb�:$t����ŘH�6���gf�4A��٦s�m`���R��:Y�]�ҧ_9gpVk���\-q�?�81����������#���w�%�C8�FS�PA�2Q�ѓ����R�k����&Ժ�LS�B����v��#؃͋�A$���1Ã�:��9_��^�g��k��<?_��I�Θ9x i�.�Y���+�9@g��Ϡ�x�(��3��$�&�v$>y@�I�!�e�fG�ڮV�%��IlN����W��O�C�Ğ'���?`h�Ǔ��z}+v�=�]��i��Zsf����[E�_�����b����3��
�Z�x�X�y��a�-Oi��jc�f�}m�tU�0�2���)��T�X�`1�v�s@Q�(:���XD|��@g/��y�j��"ZF0����/��C����G%��_�?dr~�$v�r1ֺ�a����&@�����`YR��ŏ��%��ʣ�=�6 2 zBm-NΆa#���H�e��,B]���W�g���I
'���.��'�b�Dg�k��e�/(*���ق�����8�Qq�V��ںM��)�,η����\v�����ӳS�.�������'d�X��+DP?ڸ<�jw^�,��S�>�A��c���i4�%�y�F��#��3a��	8�)lSU`m�3.(�,S1X�4���U[}���.�7y�>�̾�_���5��:��j���4dp ���Do5�[d�2F�c�"1�Vq�j�cdb�ٸ��
J�E¿�z���3�׍�3�z�1i0��]p�U2��q��H~S�B�B�w�G�"�
��*�{�?f��h#�������	���m8t
������M��0,xj^�<�e�#Rǯ��R*�qV��4B���]�[��l�:x�ʻ�Y�Q��y{�L�2�}��X�u�v�	���}'P�������@I=ϿɈL���O���Y
�(�<����M��C[�T�z�Lߊ���`��H�����DL�#�FFze�H�
�2���@Q�7���B�Io��!J�X��b��Iڴ��ӹ�Q/iS>Q�_�0��=Bh��i(�Pi��T+��#�i��~~~��*_����cۨ�w� �)9?�G��e(O���Rw�&:���=!���=qd<,�zx�2e�xł�2'O(�^�!׊��Ǔ楞��:� V������j���E��O�Ǒ��H��]�&�T���V������)���X�Q9J��-���ߝ���h'E��Wgo�J%� Ü�����y����%����8#�$��viT����y+!����rG��VA��I�E$��n��n�.�S;�&����Y*�x������ۙ��'���kb']��-t�J�
��~�%���7�˝�;��o4���Ź2՟�W��ؗ�L�����XG�|Mw�^w6oq(wP�K����(h�/_vOs������f����ʇOt<�y��l��t���ӵ�S�/+2ӧp��7+�/w1�z�/lMc�����}Ip���'� Ǫ�wH�5���>J|�蓶���5�Yo��㐡��t3�\��ʽRMK.�ǂ	e�m^�_}�7!�Us!Π�o�ܹ�f�f�P�:�f!����cT=P>��u([C:e����o:�2��;`U,�υ�+�^�ki�2��2���A���]�m�Apr;��>gǊ��+���ΰa؆��7������m�uO��������_HP��c��>�v��R`�o��l�C�����cLdz3Ф6r�8՝��-|.)����KX!ո0]����E�7N��-��=ޝ���P-�Kq�<����;+,�$b����ҁ�錓HE+ksH�������w��fd��$��˕'�?�ܫC�|S,���CNx�y���N�Ng)9��K�Kc���o�瀧���.�?�3լ��'��u����+����JNE�#A�x?##C����=�(�ؗ���w�~S��E�t�K}}=i.�?����c��1�� �GCV�e���_�������@��=E�(�m��/��h
�.�R�JZ6�	9̆�iCgg�OۂC+�B|}ۖ3����V�����X���1t�be�h���R���	%�ju��� ^t����`���ӵ^������9�.�Q����Yfn�&j�݇T��j�H{V���TL,�Q-M=�!s5�C-�����ɔ��<B�c�I�)�g'g$��1���o���k��	J]��<�l(9���C����6\���	�-l�z���>^��9�ӊM�/��%�=��lxD:����ṛ���կ,W�k�P�]�~���ٽ�=n�ߪ8��j���˛�w���\!U���Ef���2̚v�yυV1�[f�drQ����yv��u���̯��?w%�)��+�;����]���]���j�ΣL��Xyl���������i��xC0�\�]�]��&(��F>���x;0����qΏ��狘Umtx��`|�����Vg�@�B��y�)��ܼ�,�L���W�hP�Ӓ�?����s�Sا�� Ã���\�˝oFz�)(W�ǐ�-%�ۮ.'�}ؒ��_lE�$��=��|Y��*��oM�o/�`��+M��\'�'�w�W�@>�qt����ѽ�Qظ]N��a�=[�6���xԼ���>����P�X�0�5曆����v�w%1ӵ�{|�m�h+��o5!�_K��P)Ͱ�9��9�n� ���WY���pִ������YC���R���%ў����o6gM�L!����T�Pp[�����o������k�G#� l��:�j����n'�C����2���� �ڌ������8'f�L�Ȝ�f�r������{<F�r}�L��7�4���x�����9!��� #���BE(�ր�����辅��~ju@�%`�j�풙d|m���d�lS>���#s�m�fΥo���M93\�'ݍ���n�Si�֮/�%�&џ����Hִ����!oB�y���Q�zJxq5DvcP۴C��9ūq��7�t�>J�_����(����8H�ڸ�S�>y��H���������t�b��bF5Ѷf�R{�4v�_�K+��P|$Z�m�;ў>�f�]_8����X�f�1�IK�y2��}�>��*]�«��-�	W��:-`�M�Hv��F!��HS�&b�8%&Q�̪��[�pS�v�o6�l�\��ʜ�v����N�������C���BA��Y��#v��SY��⼇>�}pZqY�Q8�8��j��BKc)S�A��@��^�����]0�O��s��;���]�QNv�ei��)ĈY��ZϚan�꧓|�.՗�J�:wLĲ��	ɢ�?�q
z�"�[0��]��1g¢r�k�/0P ���4�fF��M���I:��WGQ�Yf�{ �mC�𯴡&A�CXE����GCv�.,&R4�<�1e�tљ��e�2������u>FN�	��WG/�a��򇶢����>^�>��y����`M�TmqP̊�n�W�q������?�1��;��v�	,L�~d�.sJ��(E ����5u�EQ�fY���i��:�`}\��T4C�c#���v��w����Œ�J�p�!(�q�c���Y!����Lm��e� "��$I$UXm�d���&$�@	�K�����c�<j��W�>��̌%�5�J��	 ���ӟ"e7��ƒ�;qХ4YԱ�㥯�P�@ˊ��)&�ksϱA�A�r�K��"�������@b��>F �O�����~3�)��9�`���ǗL�9��y�{�A2ω����~> ���k��m�
ʘ �m���BL��;�.šXsoddĂ@w �b����?�:=�ZeV|{�)���]K[.!��_���"܉}S	�B��`��*�G�X6�h%�����G(dv�y��N����9���u2�ξ)���=�6'�_P�	B39�׆��1����<�R����g���'�pS�
�;S^���[�+w���K'm}7��"&l�Ӽ��A�R�N� �v�X;u�l��֧(�#{�^,��5;�Q4��l�-$��x�sw��������]�>^�y����,��$�(O��9�ƿ��=F�K��Y%Sf�C3������$��e�{�W{8��im�}�p	���V/|�KK�ɓi��]qj�L�5���.#�5���|$%&s�=��C�1� ����Z~%�2O��+��$c�Z��i����s;�*�,�	B��rR[������KBii6۸4��8��)It[�(�4�F�;��&�5b�kh#M�3��(���wn�>lZW��?:D,X`�"�H#z:�|\���{S5�Ub����b;�����\]I5͝�װqF;e
�8Zg���X_�@��6;��HEWC�<2�(:������~�ߙ�KO�����yyy��"47�$���������0��[��[��Ry�h���F��
E��;�f�>����@�x�2���S�^�XJ '��`!�d�Sʚ�� ��ϋ6<��uo��)��J����u����6�K�o��-��%�����K>�$��}.�����o��-��%�߿d]Χ��d��8�k�,شtQ�k	�w��'?�9���NP����l��b��/�G���8�E�b��դO]���YS����I3�a������N��l��_��=w�=����_�����Ԅ��<�x�΢G�9�X�x���xYeŻ�p���lʷ��Lr�W���'��+�cC3Uߥu3� ��X��%⋞k�r0m���F����+�
�/o�Qx���H����=�0����Ig��I��Օ(D���u�'����3̓��ȋ�&o��}7uss�����L�n�1���ϒxmК�N�:l��������L�M��͇$Ѓm��.%��1~�;��Ï�S�u/�X9�<��kj'���5�r-�G�q�o�+**X��sx'N\O�u���fr�����|�����!�x���߾~}��X;���e����	�h�Փ��O<w�ɝ���>������!��XK���&�`����yy'���S�=_
�ք�������'��3�6�T�VR���/�?WH}nP���G�w�
�M�7|`ZC���hu����)\+#q��;�sVV[�f�]mt�'�����c��]�����KľL�q����޾w���n5��8�u���())��}l���>�����<��%�t&O���Ŗ��$��Dٽ+��s�c
��z۸F�]+�g	�0�����ݓ5�L�z2w��Sh�ME�*�՗s'����Z���m>��K�~���4U%��d�](E'�<����Ν����Y@��e�zI�K&����`�/x��X%��ܖxhZ�&/#����G���@�}_G�����/gg�E��1�8�v聘�ĜOn�x5U��[kIݲسg���7K���{�ʪ�P�j �h���ۄx��U�yRNJ��|֫�3rK˼���HI��K��+6OP
*��W���}IYY�>�٢;M�:�}�$��1�U��F@�͍����1#���l{�
�]���RZ �=�j�٪��u��a�����x����.��'$$�$���i3�6��"�����ay�w�=�<�#��t��|����P��P��5�p���YƑ/⍿��P�T��L"W��^�H�h��}�����¢d�]�=��t�Ѹr��"u-��K�
���N�
�	�]�FX����z�t:f�0�3yx�Ҽ��ɵ�����������W
��S2k\�򭶬�Mc�QV��t�o�uN�Hԇ�"��5	��ș qCR�����Ż�Yj�l�c֬Ys+�Ħ��� �`9�$�G^�g�2�Y�y}ʑ�	,� Iu8��j�+ٙ�����;�(��}��á�D���,z�֚彽�1�!����ew�0?|�p���=d��5�j�[Z���;1P�rQQ����_��"�R��h>�'�ؓ����g��QZVV������� Y�,�Nۯ��C�����E��x4�^�xx�9Ȅ�܉����x����v)H�7 O���d_y A�	5gq]��V�%T�-n�U v8�i��ݻw
�`�����H?	���e�4������ڊ�F�U�gj;;;���y������,�r�'D�ꙃ	N*�$I�l�䜳�@���TwVXX��E�~g �/�P�=f���C�s��ȓ�ʩ������ɰ��k��ҹ�o5����K��8�@���Y��\>����v�)l.�6ـ� ��l$"a�H�����>8!^�q�"�2���ֹ����꠨�"��و0���6�����[�D��kп�������UZ0e�jEp��Pҫ�4�*�77���;�(�����_o������&3D ���_�x�K��no�N����>H�J���)������V[FH:u�C����g�G^nt�����_�ǲ@Ą(��9�HBy���c�Zw�\i���颦I�y�!)���l�o�o)�eOw O��׸�e�p]�V�U'F�}����`u�h��j#h�8aE��\��I��
9A����~�@4�u��ȠT�AX<�a�?}}}e���5i(�ӭD
�Ҋ�XND��F��g�\q�;��?u�#Ȟ_ӧT�^��F�D�/O,vPШIZ�0$��XG:B��s���ψ���G�������\�Ȭ���Z�S8Jڎ�6
OĔ��p�3���3簦�8�����`_�l�$�����K=��K��Y����zezhl��� ^DP糳�S��?��z|>��
�����+㇓kX��<�Y@���T��c�����	3�F�ӹ�\�����dw?͇��SrEݜ�?)������X��X�|#��8 .H��.z���ϟ>�vR�%t�p�51�c�%�������s0���'���NЯ���Ќ	�Z����_�F[
O�6�a����0o����(i@n��H��Z�o	z9-6+s�/4S�U���l&(9���!�-_JN<���%H�6��
��Z��Ʒ�ՈWx08��Z�=�����	�����ju0����~��[|IFٖ��������|�>b����?%�>e	.�qV���>��V��Rɾ��Pv��̿�P�$� ��{&P<�d2&R��ƙ�!�(h�M7>"�=l��F�;�NG�1�"#�4+O������=_A��Z��KI��F��0z�\r)��V�t�^<ovtt|x�j��ϗ�9c/�:�Iݸ0�&-H\��SI<����j��ӳ�=]]\��IjD߲�]_�(��-�l�PeY�_����3�a-Mf��|(`��� ��<�{b��5
�q�[�)�9���<��]X$��HpǕ��ֺy�~!sI@A���_�&h_bz>D"C\C�za�����P�BfZF��cFF�6�#��8~i%?��}~����BHpH\k���˗焊'B "<�㡥�l2����u=z.��W����B0"W^k�����߲�ju=BGuʈ�|�߬A< �?P<�3���2]P�z+[�����U�m;���o�&:V�	e]�_[	�J���u�\,�E[ֳ2��4S�ѭ�����͑���D�e�SI^y�
Ƒ�e>h%��ڬ�0J�c�Z�٫x���0�[Éߕ�:q8�7��
�: ����ε3@?6-�hu��"�����X��y�p|����=�`��f�sX _�G���sQܐ�3ӎ\��O���5�m�v�@1�����7h��a'lE��`����Y4=h�C���	�$��P���Ȁ�%LTM"{��v�#��R��i�lBO���S���nd����c��pҘ�U��ЎL�M%g�h���� Z��v s~�\ �K�Q�O@ �m����J��@�/�<�qߴ�w�\n�Q�AS���|�o� �@����3}�RG@蜟�t �PCÉR%�A���N��p��Zm����D~P��x��6�0�X����$L����P߉��kyAb��SS����$$?w���E��-m�D ����ƴ8�Լ6�p/mQ9�b;��S� ­�ʪ�<��%��,eS�<���+��\4�301�<���f�!F�Ӏ��|��K;ہ��������G�Y�ś+a̡���'��$�SVvp8�l�� ��fNc?+##Î�7tP�1�pI�M����8��|X�q7��p�f8s��������1ϒ��o ��^^^Q � (ـ�,(���\%��m8z{��K�){{{;gg����b�yN�x��#vt,��U�|�! �K'�}�&�P'Z�PE1p�t*����u-GLjz����ȴz�'���T~��~���Qd ���|T��\N�-�̾Π%>�.k�d���5B�p%�A�b���<Fm�LiZ���\���5'�[�Ò�eAAA{F}x�S��C2�(-�$K�s����x��1	�7������gTy��
�4��F|��Y#��8`�����	�Y �g���sEX�j ����X��USR�K��Z�3��@q�z}P?ꛠ
e����e��_5�����j���L>�&�/P���[s�.�1捞6�w����ETDd"b��H�p[#
��䱱����p[,�@heq��+9g�8�UI�;Q��`pĆ�y���hsf����nNN���C�M��p�7>^�� �Ċ[Ʈ +;���L`Ts��MM�
�\�)��>yG�T�t�)�g�p��_��^K�t޸��y�>�tC�'x���֞#)%�IƝ����?Y9d����@��m��x�u8��V���Y��f6���ڞ�\"XsJ����%XM�f�!BΌ����?`l�Wu���(k5Z���'p�ף�f�&��!dw��[WX�BLG>�_r3���-?:D��!=�PE�e��w��������=���}۷����"�1�_~ �DSq&Y���:VHܴ�8��&t�F�y��g�-~d�%>��ضe��%��P�YXX����1=��?z
�)` ����BjY�tYY���hޣ�,�f�'�I,C� EFH�tΨ]FR�,/�b�D����͓��������3O�bWW/�
N}I�Kh�@q^b�&b)S������\mVP���Q��C���R��,/����]ڰ�����d��k��Czu��@PN2��8<KQ{�k:�O���0gB����|*\�/9��28��1n��MT�G�L�^� QU:�WUH�d@M>m���"͎���/��ֲ�xВ�ɏ8�GQd��gl�l�M���6O�t$7(B$)�?�VX<��_�I*q�'O�o.	+��&�Eo���q���#VA]Э{� 1=*��7���tz[��W-/y�% 吺H��#\�'Z=�<}]�f/R�)ݍᤴ]�.�1MnO%�8�+���9V�a}Z.6�k�__�H8��gh��Юh�#�:(�Qp�[�,��V�At[ �������}�
Tx%���豦��ka ���"V�5�^�SO0�J���9IV(��r���Ff;�<��K6:�&ЋU_�F���t>J
 wW��w�R��y3Pdځ�h5R�ǝqrrzO�l�4b�jM��.��[g�*"�"E�T�֊@��X�j9�N�q��2��Zq�j�	!wb
�c� m������<��K���p[&��j�� �yJ�r_���	����a�c\�P���#w�(#��8!iZ-��8���G���5>�Yپ_t��ĸ��xv�����Pe���Z��ə2�Q&�����[�?����{x�}�4�b��A+��C=h�C��`w(½���c�PW�����eQ���i��k�3�S�1���SS?Q�v�0!��oUD�2��yyy�'��o aXS��܃�e���4���Y�A�o�6���6���Ci'���;�##�j&�BB�c�;::��������^�)�-�ide�_ī�q�����6@��$K (�Q9߿U%eDEE����S'���M����42[���@���W.�����>2`ooo8�D��Z�/Xs�eJu~G�q]'䖖��s���x^~~~&��<����VWWǐ���(��	�[W�e���ͳ��/����8J=ej�/�A Pt%U����a��x�����J��$:��vǓ4�+��(a���S�œy�'z�	&9��� `�#ěڈg�!�Y���8	�!!!7�S@3��pg��	��ё`"@�&�~y��w��PHyrJ6���r��ǜ��B�ĨD�)){(<�6L��R����M-�Pϲ:�:,���b��U/�rw����ꉊ��Kӣ��'�j�~%"<(Z@:#�<L�.��#e�l�"n���h�9��[`,�Yl�ᘱ+C�w�v��c�qU�ZS/�a�I�s�.��?�k�iϞ��h��p�S��p�r�3��3��3><��F7Q���y�����.���!ƭ��_� �>�$w(C�B:�viA��Lv��rd)��������B��&����Ԡ�FQ���Tdd$���@�����X,���*a(�R$_���ܰ*y��4t��	����H>�r�Jf���mkKX^LLL���F��Jj��� ����	a�e8q�L�np�]g�?��`��.�o�}||0�1S�Sj=�t��8*! 	͉ll8�p]��L���|�O�ƃ�\��"������)D�IS�V��Q�>�ycw*΢���l+
��޽k���1#��J&Ҥd�1�'Nl��	B=����b�<�?�`u26>�Y�m�܅�x�:���<�	>�|�\龸p�_.��}vt��_�����/�Y�����}i���+^|8�W���T��{�$2<<gC��8�t�НOt�@�V8d�>�����[�Ŕ��^���?��p�9U
�[ww�a<���ד�Iii��N�H�w�*+QJQ��fy�'T&����f�l��f�A�6KrÆ���ʄh�Ș]L���29���"��f[AE��왭H�����$�u�)�2 6�>��{	6���%ǌ���-��(,$)�P3���144D�*�P��l�'�рqU���fnnNOy�2]K�!(����^�����e�C���'FRa%͖�2��Z��g��@{a`��šq��]���ߠ.Ȓ�T�݋'��ت�����o��}J�N�X�c`$�ܥ���
tk�H@������X�q��o$ZgS7���[F}P�Ћ�n�@�l����
�4�y:�]I	�ܓ���ʪ�	dޥ=�!�yU��u6��POS�hUU��E�%��~w�����v��b��u��l�0)��������Ap�^j[�/x^��<�Adt�X����y�v�eFHH�+����i�e�}� �Y�ٍ���;���*����("� � �
<���@!�.E8ST
g(����h����^YY��`0DvGiwrJ��|<*�s�ܘ���`��*咖���Rge�m���xg-�e=?�^*VR�p-c��ى�X��,���A	��0���̰���qn7J�S(�~Qeq�H ��@L�0����[�B��kEd��������* �����MފA���a8���;
�vy�`�VBBB�Zu�����zks�y
b��
��;)�q]�T���ɭ��t4�P���0�ɭK�:
[��$G���rѓ�[����B
=���(_���s�b��R���&3�(r_��h�A��o�⢿����Le
P&���5VVVw�\�}�H�c~/��u(�|VXX�	�&���@ſr�d��&M�UW#�@���"(	}���5���Ζ�~�/���dan���[�&��$�Y�%���=��f�T{��u}�� �Q�SX�S3NWRp����2Ț��3���G�[�D=i��z����75���T��F ��:��w���85㢂n��g�_h�ۏ��m�4��#��F�u�>J�&�x6d� �-���QY��Y����?��/?�`��|�-�"�iuP\�elMA@#��y�������&���/�ߓ��E�=��<��]���j&�ZB�GB���p^OO�~DO �/%%%ɓs�0;/���M e{SX�cF/b����ւ��B�Y*"**�Is�ޔй)����ၫ�s���6T�3~b�� n��_�G��N],Ėc�9��!іd�V@���>}�l�2u-��S�+���져�|�L!�����)�r�{zJe�x�;�7�<�Ig.�^Sb��␄8���F��q���h�ԭ������k�95� �S�11��Ȃ�@�k����LϿ��z�-]��MK���/�!$��������FAK�A-9eC���N��s�\��x�[j�s��A��{�6�� KB(N�SI̤�^p�'�?DS{{;V/�H*"�@�JC6u�?�6*I�9.��]Z��<kj�2j���͛'�a���F����,��o:f�p���\�
J���&M�uc}�<���R�-)i�8H��AW�A:�:�����Ɍt�*(ෞ����~|�J >:��6��ņ�ed���܉Ȋ�+yu��*C-�/C��?L�j͔��{	����r�^ ��k(7�4��$V=�	�U��ng��x�@qܤc�;���_�*�jkU��*jĐ������&L!�� )]��$+�E�?������p>�_]�p�����d���hˏ�]��㸮`��"u�����It��
���i��y8���f{�={���7$)���� 1Rx;B�6T[E�?Խ����STYY��8��i���kvv��^8��n��0X1��[�註�ɓ��H�ߒ6i.jř|6��5G�ʳ7/�OB��)�vv��ĩ���Y6�Kq������kɝ���p{944�:>>��q
�,Ζ4}�=cF��l���c��2Nx�������)������c%h���J�tj:Xt���^�s���� �3���>cFRYC��EM�hsNk~o=�M��RK�����"꨻:q�Zhd�_D�$vU�vu��
�-����dƜ�9��ܩ`c|g�P����:ܱ�����v݌2��@�(�;�R�[���}E;e���BB�ׯ�lE�!P���H2t���+�f�+��4*��胢�r�AH��������
s\��#,2kٲe-Ǖ����d�C��-	�v��t�רm���(	Md:T���čj����:w��T"��>n�JK-na�T��fM<�X��%,�V� ����iOi!�ˍ
�0����-B	d\�3��LF����1��G�\��eu`%����B�����.�P�M��8KV	]L�t�vnAa~����F��� �(��ʧn#䍠�,�~(R�=���fc��������"&�e��*��䯽T:�|l�+�*}98�h,z��Fc�*��E�;J~$N���[ϑ�-���f$u+,2�c�Us�m������P�Z~&y;�H������>��d	��ɘ��I�,C�QUPQ1DwlS�.S�����W[m��t�����I�f���Ѝ�j4fs�����86�v��딅E���F��`Km>|�ø�ĸ�A��u����d��Ý��;���b H���%]I�~`�)��,newi�Һ�e���~.Vl�NQG��� �R���n�����a'���DP���PE���� �&漁�???�-^T(>�#�uQ����;af�9�F����J��0&�:�!`~](�Ѹ;�Z,�e�>��m4�Z�`@:,3ĉ�j����P���� ���
��0Fe�??�I��j�o�����.��r��-,?����i���Q�n���|��.
rT���u�0�y����$h��ʔ�]��X����`��S�U��pm�S�P�� �hHS� �(�ni>���ゃa!���mSb���8�oKS���V��h�|��g�I-��dS�YJ-�������|F�����W����}q�f��uA`�S �A�������=�+9�2��`���F�F�����}H���H�ڈ���[Z>N���\��X!tQ3����ͱ��/씱
g\�-?�]RR�0�9�f�P���n� /��o�@9�~jRC-���0��F�E��F��<�e)Yp}��3NǺ�x�������f�jx��m��F���N��l֨����@{
JJn�p2�>�AB���#���b\�a���Z�b�Y���N�]�J��j�Lvs�]���W8��')��;-�s�]�~������ҌWb3��7t��y�A���r).��Z�mgt���$@�CЏ��{�pRL���!(555�������
�E��'�_��t���(�ۻwo����_H`��dd���h�q�f4���`��2gv��r`n?�Nof�s�љ�ϫ@G �W��N}�1ണ�cjr2�G\�ǣ��3���J����c�ݨ����JR�JY�7"ԸC?�ΏE)�9.�����\�����G�������e,5G���~*�M��CU� �
_gq^��E:)���w�Jbu�bG������ Nd�}�*��P.��>�4x�d"/��.�A1��F�V����W2~*#�E�E'G}H��<h�f�����d�k���erB��w�z�3e����e�{����}������p3�L���XRJ�WWYT�4w��|/�.����c�GL8t��h';� f//���˾rT���<qpwA�7r�����g��,��۱�����H�rRr��\=��0�1?�@L�����o�g5G����o�z��n͓��P ��W�but�Y9KT"K[<������S��#��������v�������>P,�� �78������s4�eTʍ�_m���,�_9G6t_΃���#��s �wU'z;2Rt��Hڛ��%$��֔3q�3���k��mB�}�l$B����K$���&��� �nnn�x��n�OhM���p�g��+W��%W�b�{r*G�#��S1{���[��w�U�┉���Q�эS�d���	0����?����P���H���G���P�&'�����Y46�?���,���.f��S1�@�����IM�y2T��b���@Y06�}R��ɓm1B��q9F���#�;�er�9�a����w˪݇CӘ
��C��1�l�N<;-�i��U��%���`����^^#sdM� �B Ta�s�����IU߂���<5o55I	�s���/��֠�F|�\��G��w�Śs(u���1%�I�'�F����	�(ऱ���`�J��P�Yvu�;|���	C+u͕5%߾Y��~i�@�!��# �L'�i��=������G��3Ô�jao�U>���S{���s.u��Mʺ�~�3Ф#��
���ohhPp�)-8�8���b���MT���ԥ����@������(��kMv��;枃��� ����a�Z��5�2�Y�zU��޼�Vi��P�37�[#e����9���L[�#�d�ɐ��S�ټ;���Y�c�����n2�"�� |�N����":RJ��p�Z�����_<{�i6k��ʷMv�R��8�8i b瞢Yk�x��
�b������Lf�=����,�_�?� d��k30�t����DmIKo��ĕ@#)����minc�㋠��N��P[H"�')Jk���L�	�bpP嫑p��1�oі�ѭ��wO��ߌ	C����������u�WJ؎���+u偑��Ē,vN�6\o��N5">����T������w6g�D~��Uw�טn�-���l��$Q�BX����.��(��luhv͊�oy
���Lg[a"�@�
�F�eg]�=�������1SH�Dtrtt�̃!�٪�*����-��E�����g6�N����\Y�#�g�:�!�RF����!�lLLLSY����m�;��"/o�u����������6������!PM�����H��<wvvVXF�kn�N�e��#����iH#���
Q���Q�ub2�:�
���3gC��a琒���ɭ��c���n���Q��bo`��m6��7�5Y�2,�N�
*H<��ġ[[��	O5l%6F+��}��U�N\�5�9K
����,��A�Ȯo
5D��x��0����k[�3�5@�q��\A�T���c�;P\}oP8 şξ�2#4%���(b�&�d�^'�P��i�L��
m?ť����-a%�iFH�?�� ��[�1�K��y����<�*,4t�G��N3��X]]]�@�Z�qR\������O�*_��n�ƞ���]��3��
]���ݨ�1�RI]��d��?}�*-)y�␻!0��3�N�U2�c#����Z�s	&9!׮]���	�C����s��ul�*���ɬ*�-��8����u˚��ZXvǾ:(�s����<1q��O��.gZZ�e���7�(~T~�qwԇ�sO�n���p<�>���(���q:�^c���ju�|n�FP�J��/���f<o*J�˶J����8:9�*|��BI�k�-1�p��0�Z�U��"Q#U�wGݠ�Z�ӈ~�m|x��*mL~�LG\��d���01.H��O�F�s[���~��VosW����i��|(���)�^�`��]�I�|x�]���szhx8����vŤ,�|w	mN�P����#p1�ݎ⪟v;�9νh�>|(���S�f�.q���zFF�>��F��H�&�r��O0S�� ���?}Z����۶m�ɰ����Ay�����f+�b��I��t�d)5:�� j���HQ��7� P0r�j��ǳ1Ϗb�׽*?�l��+d=ř2QlNA�:C����IV���qɞ?����)�?G_*�2]��<)�>�T��"�����U8[Ҽr��&�~S�a�w���u*pa�sNYD)���@�N�8�`啼�]��;g�-���^o�o��J rA|��K=P(0�U[���K�ۊ8�(S���'~�8%7\n�}��Y���R�0cU�ћ ǀq���ޭ�o�b=P[Gg�)��z���iiU	(W-���
i*�)��*����肂���U4�riiitC�xdVF�9ɽ��2+>7(�ڟu�c���]:uo6��x�ړ}c��o
6ų�[l�ɼ�|�w#�O7�/N\���xl8�|��ݛ��8������2�w���B�+V�)�M_�h���d/t_�(~������/_�|���;��x�L�;IjLl#���,}���;���MsR�tx:T��cN㥆�4��!>��}9d�c��)4?CΫtp_�n�JK�v��ƪ۶�k�%�U�.l��cF�3���vySs�/������nm�B�ۍ�eѝ�sr�V�}D������P�S�c�;G�ٜ���.o��~}�a$5fJnl:��ľ�z���W��]��۷:����Aj��j�W�����"y�ګg�B��i�9(�G���;����
a|{��!����o�������w�÷���u&����Zf9l��K��:7Z����[k��>�\ڄ1݅��ͷ��ހ�_�y'�}r�s����d��&2��@e�M��99���~5��ֽ}>6��oP��.5�	#��
���>�,�qv��<� ��3�U4��_fd��{[K�q]%�l`|��q��xX2��PoKR��,d�s&FF�I�S��m�@����aٹ��*����v��7�p�4'�=�|*b��cVR���Z���c�߾=	�9�A�@Z�,
�55߽{���uF	��ú_�\{������\{h����Ȉ���䋠ht�)�u�_3z=sTSr�����8���KS�g�svK����t��܀������!f��Qf ���y{_���ŋ��7\R���:�h8�|�ңŤ��<6�)<V�A�j�:e�r�	��~��e�aO�}$q�n��K��e]���#�ء�)�d�>D��D�G����IS �i��v'����a�z�PZ��QIA?�T��Ҡ%��w77�F�� 7�<������J�𲉿�a����`��d.��I&��K-�CG��d�M���N�={6fS����.�?���-If,��b������3��[-Q�$�Ӯ"l�KY�Cv�YY�J �_��j�"/��"��2�c��q	��wa���V��\��2	2L��6^���,&Iu��/������R�,N�O6b�ݦ�(���B�w���@��\l�J��f���Gƞ�.�����F1r���w�ܴx~�ڭޜc��taQQ'
��>��]㿀���@�-��O�Υ�����mD��V��o���S��c�B�̊�CSU�%%�$ �3rK��\�e����ߤ�Q3.�3jk>�60���%����}�;�ī�.DBo;�R�� �]RUq�rµ�ĩ��9��j����A�O]��'��J����0^�����2�2�+MvK@@8)�_�o�+!C�ގ�ᶸ�ޖR�HGo�-}�Tx��27���b/SRT'�rr�a�sw�Y⿛�8�4~Ǣ�oUI���ሓ����9��§�5�2�X �q�@���|FqW���(�yvuu�"{u��؛U��So��!��FJu� ��c�`��ħ�x���%/��0�܍��<x�`5�KC��杕[�Ғ�	{���������u��x�!_~�Ҏ+�4��U�sqI�k�P�$�3�CK ����}A�:��ó\?����գ*�+ �Nɬ�5�4coj{����|����8��CME����y0��A�JI���s�'�d��HI^^��#2wx�&;#A��zkC����2:R��]�I�|�ͨ��
��9}h�=aTϽ�7ⴃ��S�晑T��·1GpHt���1�m�>��[���G9��n�[e�<�� �q[�$�b%�d�޽���G���6�<H⤤8-:Y�m�Ɵ���&����q=�3J�SY�\���^���,�W
������I���
�	��\r�D���j�Ԍ��m�y��%$$�as��3:im�*�� <B2555姰=דz�������}�d�A|$0�c����~���e�ov�b��A�P8��4У~�(��2V-}���U��4�����'��*D�wp	�	 #Z�`�A��J����:�Pj����8ݠ���R�ۥ-d?�n�����nn#�E���a������p�ӄ?��}��m9UI�JJJeX(��X��ء&�ii[�Y��/8WX�ϝn9�W�\\}3��:{(zjrm�/S��ñedd��1�H���H�����TfM'Y�&f2}uu%C�[Fa$ �����N[��K�9�� '�(`6֟#�`�el���k�C$��5����dK��7��<�4@*�nR�v�^�����,�:����sa��j�-	�.��7ߎ���Ɣ�C�ݴ�K�X�!����	{��/�(�2�F�M�';7�S�&���26�7X�'��Jnnn��Ҵ̨�SD�	��訨���(�"i�Y���QE�k�=��ɺ��bbأ����(qY[[�'���d�j�vO&3�4��������b�!�8�b82DI�I�����S�֑���m�NF8�sv:+?m�u�L7z{�����0���D�$��pz�%Tj8!�)��ۓjg�υ���k�Ki))nz�D?����zl]<���M�	�XNS�R���d(�B�_��^wش��L�M�;$�����'r�{�p�ǀ���?cR�'�*��<�K%ۺ��[�(y�@���t��0��<גl����5'�����w�H�_cc#]?$-/{/[Q[[;L�)PwW 7�viW��Y��[i⵭��gT��:�A��/o�O�H�UA����	I?E������P���GZT´Q��V���(��W�Ț]F�'KSI�[�ƒ�����aJ��
�G��ނ~���9�����/�}����<���,�s�����̍���L��p��4�z����v��_�	Q��۫����_���� ;�{�s]J"��[+pwj�@\Q����x��ͷ��x��D���+o�ǿ���[.x��(�yak�1{O����(5־{`��1^���*�w`�ث��B*n��S+�w����$�OَʀΊ�I�-��������OlVB͉'w���ɚ���G/�2�����7G�#b�� ��g7�|N	(o�f#|B�x�dS5�lq�"��l���^"�ߒ}���G׭[���߭�b=y�u?� �4W(�O�nĳ�_ޯE�ree�E3�#k�M��d[��x�/�0��<`�4�^pkkkJZZ�	�BEQ��PR:�M�v�?z�A_W26𗯸�k�XK��O�>���=Y�q���(7�X���9�.�Q�NB�9E轛{"��Ӱ���\Ł>Cu;�㨑d�/��8�n)�0�U�W&Q(�F<�d�nR�$�
nfs��4����M���]]��� 4<��7��0PR+A�D�Q`�P.���Z2n�a�6^^^9����a�#����^�"����ߛs��3l����ب5ۼ�_�!���y�ga� � �~�b��4^��]%f��Ñv�n^�PD��.Ĝ���/J�����rq��c��Q�jR>I��A�+�mn	{z<�b��~d�b���X��]������ؽXzV������z�� d/�]��&�!����5�p�s�zn��U����'6�B�@�|�)h����p���+Zt���aX�nb�lsWD���-"��R���v�qb�V� ��v�?%;(���e�l��rA��Zy^ ���Cw��bܨ2	�f��f�"�~��Ͷ��)��+�I���{�����aL�Pn�O�6�s<(�Kł��kp�f�����v�oOyd[IP;��l�=۵1�M�¶u3��(	3.o=)t�#>��< �S�T�y��k���d�u&S�%�qHd/�n}������0�\�������瑧��*�e�B�.!�b��ح��?{^�5�T�����ͻb�y� }��É�Y؆��7���ěA�O�1��lq#B=��u�u����؅�3�=�Z���PUK4�]{�ڶm�7E�Q�r�XX��]x7`	e��G�5���5~+�e�
)l��^g�g"zI�Ph*�� ȟo�Z&(��p,�y���-h�孕3�psN����W4h������Ӎ.�Q�|�q#�3�>�X����"4=���<#(`D�������I��\��f<Oj�	E}�M��2	�5QUchV�-�VB�2G��ٚ5��~붉���~iI*�������`m�al�bD�-B���)w@f5Z�<�s)re�Xd�����V^�t/Gbב2�CO��7�F��6w���z^��
X8�*CU��CQ�z�A�]��>5!����铃W��F��"�~pJF�r$���ʾ�r�-Z��[v#�	��5=����
�=C��ODZᰤ��T�ķO�V��l��"�d+A_NBOV|��9�1c��{��En�=l�`j�g�A�/�rs���+�x	�^�GL��=x4Y ���/~RD[�эj�;�Q�ȝx&a�s?� ��D^�{%������� j���{L�<<bjU:��N��"{��M��������In`�cUUUx����^[[���H��ߔ�F�}$x%�{d؅˴���pD_��(�y�˯_�ЍS+� -���qy/
C�H�[��63�mnn��k�F��y�D�P_n;jR-�'��
� �ݸ;�yH�c�E#S�L�/<4��o1'��<y�2Q��C@
���M��0A��M6����F*"z|(��0X�p�r;b��8�yب�]�ty���M��
ٌz�G]H:��<>�H�&l�sIlZ�,��J��sm�q�,��7�ܪ�Y~�cj���`�{?�$���iy�,7�+~A!�0*%�e.6O��z��tLsGu��ː���Ti|���>�9}����rS�O.�l6)/����[�+ ��}�8m�]��xIA�K}��]�F�D�������(��h�'ZͫFPs|�"H>�Z�X���q�8Y>uC������C���(h�K�i�㘺��+���l?r;�>�P��$���+����;���]��������E%���]1|�}�T%�)ytd�l���/��C&t�&\.%�WM%�9׽@�ElS`���䖍>l�`��8l.$���ͩg���bc���Ԓ=Ӫ���G��`��-1(��T;:kh�M�� mT�i$�ȶ"�uu���&괪��l�x(co�d`��bȍ�Z�����|��`�?''��S�.c�4�\��1V��o�C��|�;s	e��IQY�x�����{� ��;���*��m�հ�sswI����f�C�[�9���+$�ʮ�V�ݺAA�0�q˘����,ǚt뢓߷"z}��ωcM{2z<*�ܭy����ȃ.��crjMTi���	O�v.�Gl�z��.���Z �w�WB�0�Kt���mgV�A�VF5ц���2	t<l�oA��Fnk:Wz��4[�o��F=D�͋�j.��a�=�ͥ��^W �s=��)z����!Yf�x>K:X>���D܎���P-}V��M�nz�J��eۅ����-AGQ'��Q��;g��o�v�Z ����ڸ�ǈk`�m�eQ��9�8e
w�)���^�F|�
��7s j__.�,�p�w'�����/i1D�I���̴���A(k�:��$�މ�D�Jx�sNl:���l���q�<tw��fQQ��Ρ�HT���=�sY���U�=f1���-���i�^��f���K�zNd�ǎ����62J����w���λ?$��Z[[�U��$#?����bS+H��?��3y� �d��d�qww���5�ޡ�-��2��@���#�5*Y�-~+�&ê(����phc�Ygo�>���B�Y�����5�(6١�
!@���x�Q���6��ˇ��ՉoI�u�w�ō��d�=�*v{$��B��h`� �1G���~Xo�_�˹�J��)���$�з^m6���`�]�ws�U��`�Q��\׍C���+sh��t��W���4Aa	����}�3@Y�~���zJ��4m���z<���)S��^ے}j>�Sa��YA>�s�ώ���R*��`���_�~����#��ΐcT0�"_籐����Hn�*���늖hH_Q��T��>z"�s��-S!!��QZ��4����������]B��Ԥ������3���=�-�������	b���á�
D�	�������@�Y� �5طg�Ac��f�U��x8�n�y��j%hFY�+ƞ�y8>0}kLOa3�P-��LP#S�3�8�;�*UR������)�rP���;� F�w�3���y2"�3��WG\�y3�����@y�P;ޕ��Xt�7&m�������N��"�a�}�C!��s��Bz�V��ړkQ?����1Q���OsA!�d3
_��*�&�ay+�V�@j�q�w9��E�.\�
X��/i�g�\ga~��c!�_�_�[�Ե%��������|�/E��)�[\u�1O�!k|�=�gI�����w�G�V6��555E�YQ�ZW:���qcwH���[_Ծt�v�"D���|�u6���?���N��!�"
����EW���A�}�{э	{���<R��th�� C�g`q0�6�I���&��h$~X(��7xi��}j����uttl���{f�ֲ�j�������$ԧ&��B	�I	�/�֓�>T;�a����ﴥ��jk�98?9Mi���	���{����5�}ſ<���8�m>���gyܲ(X��B�i	{Y/�!f��ϲ5G��wT�j�cE��=�n7Bf���[�94�����%,zt� �u�c����ϟ��v�X�����l�t0���誮��O�IAq��s����DeQҘ/}���h�(1�h��g���\�աR
@�:�DMd�o�@|���ؚ���3s
��\#��j`u�͏�6O~~���dSK�/w�\Ɉ^K����Yk���_�G���n�r��Pֽ��}f:#�<-�kW�(g�呁v�vH� �D���J�H��UE��u�5�M�����$ ��d4���$�c���$T�µ��k��7�t{�',��X>��Bs�A<�nY�������IJO'52C?+�C�i������v�/���t4���n%C��q�	֟K�c�褭<v��$�� ���(�݃���/.��)���zg^18ZQ��=�S#'����Z�4�s���k��$I��{Lq��8�C��z*�h_ߖ<��5�{<��]�*�؅/�sL3��,z��WJ��gc%OZ]א��&��"���\"��w�d1�PF��4�ou��	�������P �ʇx3��i�V�w-B�����.!�U#b��(������6QN�~�¹���Ѡ�V�� [�Ѿ�zw��k!�X�$��b��N�PaL��쉢��;�{Pz�r ��>��;lb�e�v	IC��~sL������OtjN���<�T�7:����浕�NCA~c�~Mь�?{�o�l�ӘAEC
�;��J�<��y�0����V��X;��_��}�2$8�`{��8q2����w���L��7��
Qhc%�]GB�is$��W>\��� ���R����ѫH��-:"<�`��%���+�m��r���C�M6��^�0ٚW��ϔI�F��Y�g%쏨�L���d��وi��5&��v_h����O�]��d|Muu:f�GҪ�א������Ʒo�y�N�"9���|�� �lR��ss`�����K=-Q���Y�:g�_woٽ�Tp�����+
�!����3b	m��:)��~fc`�`��'K���Bm{woQ��W\i�Ȋ���[��ͽ&ʥ:�����6��W�����4��;��e�ꛑ�}>%
A"/��uaL]�\Nm�*߼5����7o,���J�G�S"Y�����Ʌ1��2���z�C�E��\�iڸ�AUB�R�WP��=vS(�O�ݢ�5��� `����R��xr�����+�-g��<�&����c�h�[��Ѿ����g�
��X��p�:�+��v`D����
�S�ACeeecG�\<f�lQ��'�\���	R�{��+��oT��ن+�6�S�_W��w�/	?xv���􈶪�Y*<6�.O}�0��cA�f�R�_�M�J� ��9}�xw�������F���)��M��-@��4ukM�yd�H�w}o��p��[�����r�����w��6���,}=U��j�s;m���00������o1��
��M��aN�(�ns������Evo��^�*`����~++�����G"#�	c^$g�4|�P�^�W����V���!��n{_�c�]|8h8K&A"�T�	�1T&n����Qϊ��ʗI0%���k�RL��G��R������� �Z����nm�,w�a�3Ӌ��*�/���r�9���&�gL����&�tx�ܸ<��e�����<��2i(A�q�Q�D�衙�YײXm�sk>Vǩ�&W����q��Jl]E�o:���;~R�H�IE�Z�B`�6��J,�+���P}:όG�BcZ:�<r-̇(sY{P<DMvN�"E�R5�+��XE�����E����=ܻB?�t�U��0�p�`�h�h+w��.S�OG��ey9�뾚���<߁���~�
�!s,����(D�l"�=��Zg��=���
���G�3p��?@Ku����Rj���=_����^����L�8��k��^��i��/�Hw��(98я�G�t��
�|@�w��X@����s\�s�2/8R!QΨz��r��*	$ް�lM��ޚX����mn�c�Ѥ�O[��n��|ི���L=)p�����Z�-ᝣ7�~�:p��]��:��B����&�W}�;;]��R�Ie�xc�&�"��f*���lח�K"��[�U�C�t��{\��g�MGF�t��I��Z&�¥�|
[K�Ъ��x���K	9><���괟���P�d��y�����7*`
o��!ڷ�z̠P\�'�*�n�(�q���U*d��2���V�$��`c��3;�Wƞ���>f��z�p��n�b�E�j�O~��!��d��y�GW����}�St?-�j���u��_��̑���1�2I>����^ϓ>��*�J���]��d"���[��W�V?Z�Q>v~�Ґ��澚z��aa���>�
�:;��������Z[�k3����T;C'g��GcY�\E���1tsd�{	Ꝕe<�a��4+��e�|��-l�~�c�E����9(/�ۦYSZ��D��TE����X,�&�k,]�%>h��G��e���S�*1U5z���HcX�6P�u�v���T��]aU�q�4�,�-l���|�0��^־�7��~zW��{��ٍ.m��<�>�X>ͣ�j'k�*D���aG+�-u���&>��8�Gs���=�bt{k�4-��խ}����������B�x�c\
��9�iU�4��H�n���@]�=�N�h�5ED�����T��.�B��Nf[B�_^�kFPy��V�G������G�m������X'�Fcxa�}́�"�9�̺�Ci���(������s�Ѿ_���e,K�;�t�	�|% ��c�ij�*�cYn�n��*��\6��Y�k�UOKɤe58Ǘ����pVVV��W-"��#:21�{�v�dk�j���HgK"f�_��	��̶�����Vd��Zt���C�PA��1�|n���cc�49�\�kc!n� �i��K��b_�zf:��%D����iT���,�χ,���LB)��|J��<�pH�r\�	����8,�����x��H��Y�#!����A���g�L0ݩ;�.w�ws%b��6�����Bz<@O�H$	�c��yHp�]���hk��ЧbW�qow!��:�'r#�S�����p7�Myw4�1]ey1����j�鉪�K�i�FM#����i���=��8,i5�%�����kac�ϊ�h� ����ސ*1��_� �s�b���4M�Y��s���9�����ZK-o���P y�C��B	e{$�r����Q�'�E��l%n���8"��X�bUaв��[)�1��#亃��J8��d�P�J�S62w+������6V#��v\3r���ۅA�+R�.Yn/U���飏Wz�¸�o�%� ƹŬ�e^�]&���=��EV�
��i�j�c�$ �t�n�>�+X��ȿ� ׇ��,ӌ�	.Ó�G�0��J��!6t@�o@���A_��P�QOXE$kk�%ƒ��I�>���J.�MoszW�I!����:
d��m�v�r��$�a#6U�^L��y~q��xGEE���;��H�K{�1?{71�Cl���t�3p���T�.0_o��8&/�K?9������Ǉ��Ch�m�R�T���	���f_���lꝖ"���Ȏ�J��l�=�P$��-�����]�^��)��K5Q��8��w|x܄�R(�߸�@NJ�*���.I5��C�����o 5����k�Bs��H�=:2���	�:?���$���l���*F�D�&ʴ`���ÎR�c��<D� �-��[n��o��0��"p�_��1aaa֩�[�G�e��"S���u�
����+v?���}cIv]�V��["��U����ׁ%�d	
��A0m��Ph˾����i	�=m�����'�s�p�~@/b��)}U�� ����K��&K���*'i�q�.ʠ	 %n����������gʺ1B���{��U��L���^ z�ZeWd	�b{��`8�³W�l�Nt���?()C.��c����Jqs��+�}Q(��bbs8`jB��|g��P(��3n�r�A]T�)���$�I��".��"�|ZJ�s��]���E:�O�і�tT�Q�t�gx��.�Î�6��1�i���m�;����q�X�$��sQ�p�`���OGF��s�([�	�:7�ֈ�~] ��ĥ���v�����⟜�[C�Z4���X�/�T�J�+|0�޸[���Įԅ1!���Uօ�A)ѭB��EjXt֩�����-�W�g?�У�Ix��=EW�^u+����c?�%X��xB���IbQ����{�*�fi�fK#���GGG����X��WB�~WA��W�:��&ƜU��
@4����?Do�%���i������ɡ����.ז=�s�NT�
$?�L���n������w>��pOF��J1Ns��nb���9q�PfK�r*�aǋ*ҩV�#ցPt!UX\�SRbt��3���3�M$�L�n��
X10�����Ę���#� ڣ7��q�O��z#��߼R�[���<�T����5~�뚙6ڊ^�	����.h��z�VT�4�6<�e����g��nӿ���/\�rh�C���W��^r�����6��@e� ���B�D6c�z�0��(
Y�
���� pݬf/����Ry�a9�tr5c��>CJ���`o�6�ȐU?v�IL�Y��D�-A�&=WD� M��Q�pU)r�{�{

!��#�;���[7dN���mX��S�A�H��r���}Aľh!����
�;K�4���~2��	9��N7Q�vD>t����g�ea>�!�Έ��E'~"�x�>h��,u�h(1*ڂ3#�x^�r6�u�0�'�U��{�4�)"�Qߝ�tk��H��W_����� ֓�5�U��g��K�+�_4c���_�Ah�(1�V'��]UG��}����&!�gS��N<���@/��І���R���b��S��aJ��"�h�M�[`�6�s�*�{V$Je����tH�Җ	dC2dT��cnj�2���8�H��os���x�$�9GN��Kl��𢡊B���C��R �x��0׃�4F��u�)���mH�~��e��m��|�y��	�*��>YFF+�6>H��-��N�/����~+$ǵ��x��f��Py�ڏi�5ȄBTr�t�.�p@1� l�NY����\�9�'�h��m�22^�u�y�U�^��*D<.�6�\�Q���c�i�<��&x�Ω��gMT��\�p�V# ��;L_AQ��؎�4�C�5j�K}���U����=;�A��H��+���T����v���>�gBm+J����^�d�ᎇ�������.·���`�}��#��m�M(��92�"\,;K逎�!��̙�'�k�I�׻5Fn��bTݲ��D��"�iz���z�L�-�9�rfF����~�
�S�<b����=��Z��<�4�T����[�-���DT�3B(����K��.m����|�\
j����0�\`��t�������C�Aa��>�+�6/��,4^�����*��� ���}��}d;&�����xJ�ء.-�sx�.B��N(�~#U�>���}�a}���x�7g"Bh���+S&��P�Χa�{�\�w#۬A����Xc[����X445'O���>:��j�4h�A�D]J�E�	=%ƅ��t�{D��]m`W<_��K|��-�<�I�u*��.1�C��)x�Ia���Ȝ��Bn^�6`�je�x�N��r;���\����"�	�1��_�⓵�kZ4?!".S��
L��h3D�⓬TcbD)��N�YY�"Q<�D��AwM��A2j���J7eKbX$"ǋ��Ί�>�D��V�v���(=���d�P���o�նP^��ߘ��zd\�⏅���n���^�6����緺if�Y��,�/5M$̭|S�.�V�<�H^ؐKd��c�hր��c��((s� \��S�EWƌGi��7H����FP���]�Z��Hc,J!c���WD�y�nm�X���o*E��6LH� ����]u�qˑN�5=�i��'����Z��w	φ|��
oK8�v�$�[��7�_��C��2�;Q[u�
i�	8<����b���ⲝ���Q��v�n9�6�K(��\>���(���Ǭ������;h�ӡT��00�[<�t.�C�P�s�l�ǀ�(��.;��.�.ׂ�f��P��F�_K,a�W���Z����gx;����3�O-!Rl�ݑ��@X�k��L7���Sj��:^"W<�.��A_oŬM���u�S_���I�E{�vI�IyI�����3�I�C��.�-H��R'��/��誧>猎�J�f�ڌ��X�|�)ڛjb&�"�zJǼ�Tm��8"�$6{��E�g$�a___7h1(� Em~�6Qlh�-\v��ǌ��� �ֹ�!n@0��D����B��Rï�0�Z� 34�+J4q�.��s���GjJ���7��6�`}�Ay�>���	;�����^�ʶ��%��bE��&��p�|����J����r�|�܁�*^)We6�!� W��i�S���������/ ��9���I��:���:E� cu=�}�2�;E7��2��/8��PTB_���r)@[����y/����H�vA�6�u��8GnБ�$�5,=m��� ��P�M|��܋�a>��ȗ�d��`!�
���i+�C����z���!���>������R���Ĉ�e	��e,���Q��@\\\Q
�N, .LI���r5ǒ�?h�N����/?�6�5�������glb��p� pp`��;� ��~Ӓ)��/k՜�I���\4J1+��t�>���->C�6�x��qq�3qy�ձ,�GP�Ğ�/?}F䳔O����赎Od��>P>��p�d�E�-i"��t��W��D��7q3sWL��4�
J����S���H0�Y�����RL�FzĻz��P�9�-Xh��sҷ2�L�a}��r$��(����o@�t$:}vVe��v3��̚$����6wn�Z#�Us�����S��bz9�b��rԉ]H�`^C�������n�I\� ez��
����Es���E��3�Ǐ����I��nb�1(��'�W�:4�Q���2��5��5(W5����}���K�	�gn�"ӡ���gj�f
�rW;���ئXˎ+)����@]{�>I�=a=oh��sà��~���D���k�Q��et�&��'M�����ܷHj��߼Ÿ�7�z
�qLIŜV�8��d��f�F����!/�'�v�x�0�9V:�n�0�(y���(R��N_z��i�:7qziV�Eņ;E�D���F�SP���)g���(y�O��ys���;Ґ�= 3��V�a�����26is�J�11ty�٪�NvNl�S��w�	eV����J4x[[������Q�kj[D���}B��T�^v���Z����f�_i{%:�dj�(���,T��D*c�n�{�Vs ��߀s�q& �ɻS:�*��B��iuy_�!3r���Շ��_�^rqZV$+Ж\����7un��M ��@�����E��G��VhE[��-�q\VQ�=[EE���I���������4�d�i�|
ǯ E�sp"M*LzXn6��l߄l�_4��Li��.0�'��_,;�<��7z�ƚ�{�"�f}rFg��F'�/~��" }w��>-%�Y�慽u�9�A����6<�� k~o$/c�:t�@Y��zеԏ5ۉ˪���R]�ۍ�����[�l<I\t{٨V��{3.n��"8���"�d�Q���������$�4��)����%�)��i��z���Y���ϯb�4���+��I���k�JWĺ/p
�X��m��>���3s�XdY��s�"���xן������/��ײ�b律ⴵ&� ��ZB[��_7[��ˉ�'���Q??��������d/(�u�,{{���R�(BHӽaB^GN.�T�������-X�P����Ai���0��6�D�ӭG�dH~�Lfʇ%J��䛬D����`��`�KVQ�w��;��|y�������L�u��1�9��P��P������䀹i[���-s��S����I��������y���C��e.K�tkϓ#"��.�՜O�x���I����]��KPbӜ���#GrCo��.��@�H�~\cZ�� *)Ɩ,��-����^���:sI؟q�UQ��d
�V/�����c�M�V�tc������jv�}��r_�c��Vp��ag�-C�&%?낌�2ΞQחQ4|BD?F�s��ζY.���K?�x��~�$	�MZ�I˧?�I�Fm��y�����Ͷ-�z����\l/�ԁj�J���7�jS�7��_C�F��4�d��֒!��ۜ]?�������|J�5w��A��Ľ���nH 4��/3������ ���	h?/�X?��q�y[�g1�s���+�b���\��R]� �p�_3S4�����|�`��6Y�/�Vp�K��~d+�]O����'�|�VW�d����=×�DU����>G
Y��d�tYsb�I	�OO�V�I4B1�QJ�"߂����}�)����� ��b!����1�/v��"4�3T����dn�7`��"T��kj��ͧ�6dY�V�N�鿇(h�Z���a��P�#���N{��&�X��lL̝�izw��^���g�т5I]���r)P���j�EJ�{8q���O��{���i�Ґ��Ldg�L�!��z9���3I�S�͡�!�Lm���+�V��C��/�zsǩ��H�n���xr��W�44�Ox!���c���P�4�7w�N0�	բ����l#�?��+�[�]������r�:HVXۮ'q��j��#�:���F�����Q�ݽ��g.���8�~)i�Mԅ���{.Od�	�F��ͮ/�� $�
��Z����Cd����I��v�՘�d�P.Rq�n`�����9y���-b!���L�Q2�𬍫7��z�&XL�lҢ���͛-j-s��TfNaaaZ��?]���\�;��VZ����=\��b@d��[���[��O{6p&�3|DJ�$��'C���o��c�8��E\�*-j�}ٶ^�7�)Z�k:�]��G�"{�bּR�6]�w�%�e�F@�~��ږ#�k={e^{��M佃�]�O��b��ݍ���G���xKP����]e�n?�D�v�J-�G*��H޿���C�'��	��F�&kE�wT���5�Q��ӱ�]�Hjz6�<6�ҁHT[/0;�5'����')�i3�ޛDQ��0���i ���"�p��\R�ս1��=a,#�eVw���+�ߑE�U7)�6�Ns.�1M���y��&g�ScHݟxm^�v"�囧c����1�W_�;q���I7�秤 �e�0�. ��!��̀,Ϩo/()�<��o�@$u5��e�=�L��[������3��"������5��hTD���T���[�#���b��R.�6�}����܇C�d*���y2�S�f�b}��F^��g&�_Ify�\���Ə��b�a/(��͏�m�3X�qN��h��w�9?�z+r��$�T�l�&y��ȘP�`ˎ�#�7�Uo�����^��Z= �3�%�ۥ��ѣ�T�H�;��~�M0���?gL���#I5mK�
�h}�c��+�ε�w/������kg��'��h@����h�VE��jW�B���X*9���6̹�^�E^]�GMH5�k���r�<Sg�BRS����\>V5� =������͊���͙
�%�S��������y��EÚ�����4<îs^�sB�;�O]b�i��#����tΌ$կn�����Z��8�39C��\1QrV�F�&���(�D5�	F�̇�{<�I@luK{��RpD���d�C(m��1@��jD5�zq!��q�
wD�~,]U�+���w~Ո�R{�9jο3�3F^�G��_��S	�׌<�T��_*�9W1ƍK�t�l#.���3�%S���]���äΥϳtJ��+�ڟ�fA�9��.��ƶ=�X��a[��b�0��.��1icZv�=4'U��,�&MΪ�\5�����T$iX��齦�II^~�:��	��?�4����������n�܎�JY狐���E������ ��'�_m�)ɓ_�@�&��!��A�w����Zh�m�TzB)\J'EL�*-k"'��ɽ�������kH���(���j���<�'mZ0\oh���?��lI4�����s��&p�O�K�鄅|aW_~�:$�B��=Yfz��c�W{�z&(�݃\妡���c��v�֘��HA�M�E���݊JI��ʧp��f �C��j�z��GoN0��$y���2e_���w�r_(�:�`M���^~��q��u|u�����.���2�;d�v8���D: ��\| pV�x�=qm���'[[�LC��E�Y�ԓ�����9WI�������|�������1��Qf�}�s�1�M��W�B~��n����y��>O�W��{c�h��f"���"=�$U�J��76=`�ѱ�^^<���7���K�jo��p��N���@j_%��R/a����ݤ:�w��=y�ş��;�-��h�F�0��� ^^=i�W� <��_OZlE����Ɠz�o�ym����ɚ�X�o�o�U�u:�E��*�j����2���[v������h&Y�br;}�K��a�?�.�F��F�<)��ꆚOUj�
�T��F`�G��b�X�'RIqX���䥟w���z������|�ΗG��� Vhc8-vo)Y��R�P�C� �Ԏ�����������Tְ�Z�ɢ��e=!,S|��g��|5%��t��c�fr��(������9�?�*���dpKs�4��_R��F>��z|2�2Պ��ɾV���G�����!��m�:����0�C�򷏯���[��,-�W{��垭IQ��ꬨRM�D�wW��6�i����mq_�o[����\30`rt���.��"G��$��w6xl��&�������?a.�,Rk0���Z���)�r|�ț�H�"���5��C��̀��/?���l�GY�al�u?t�=4s��W���7����?B\��'%�D䔶�,$�Ψ��ۘ%��0�"�f�C�P<��~VG��F7������*��oE@��>M��q��R��mR���E\~�Q\ET���q�����`C���RSW���>S ͹#����<59z��#^�e���ڒ���2�SXJK"�6�9L��|=����hH��3�k��%���\^m�>Q��RF�&ҕդ���~?	!���k�?�H�(���/��x¿�mˋ;������ |o�U**���?>���A����nw�s\a���������f ��u�Tqc�����	0�U��Py��6F���Z���ړ�"��R�%�Q����׃���))� >��:��_����A2����n��u��E��|6�����f�.y�����E�ʿ�-�$=V\cmRJA:�U>x:�bɘ�\��UZ�T
ō��;� ޤ%ݸ�<���i*BR�bJ��-�'q���l]d*��;�5C[�D����$�C�ҁ+�o���&�0�1�M򿙙�b�!��8ȝ�_Sd5���^X���)���8���^K�k6����Yb�;7tU3o���Q��1�G����b�i�@��.Ss�`��*���f�B(����>�mX�8M��-r�����,�c6�}���*��MXwJ����9x��7�� � ��7j"�Ú���st��P*n9�B&6�)s8� ��ǧ��
�\]T�%�16f����S�7=����lT�L��h���m�y��ƩfΔ#��U�%�lip�)�S'���o��9��y�����)�z���0-ȥ�W)��[�ѷ2���9ØB!{��t*�HϺ$M��zu�Cv6��=֨����{��J�`c��f�,�'�u|o��6dFv;�y>�5 8�O�-���6=���؋������=�6Rn[#�R��ߥ��t���Ly���7v����=3�9�g��,]�@u4�d�t
��4�g?��K��
Ƚ����?|�P{�
DnD�� U*���0������!ޑX�֪�-�"�v�o�Sy{��B�p�fE��_��K*)����� hej�l���}t���:��j�]����C7��w ���@ͥ��Y fRf��3Mv�K�;[�M	c��6&O��4zaa-�%-��Ĕ^�B�?��N��<cH3�,���'ͼ �������u�b��pE\�����ƺ�����,���|�v�IGn"-xV+h�&�s�.�&Ś,t�B�������L��v@m���o���'��U�oN����~�*�����$}��@�:��7"#�v�����q4q��0.L!�ܖ���tNZ���YI|�̣�PԒ6�����w�}��ݚy�yC1�w/� mP�ܓ�;)��ܙ���t�ӫ���� <+�@�bm<��^sZ8{l('�,��sڧ�p����1a���Q)�踁�-*��K-��,��R��2��b�,h¬��`rAH	��[�ҙ���3�-8���	@߫
!�Q�uv�T����j����B�-�$l5�]GN�$����A���&=s���VD���)wܥ�8���q�;��X
��E����ωEĥ���@Mo!��m9I��1Y��$t�b�o�����E�M�al;P��C";���� U�C�:��|��pa�HB���0��FM=�l ����jF�u�uZ�,��vi���p�9��0�����%z�����4�3��`O��P��g��zL����Qt&�ET�Ĭ2TN*d�I��Y?��	�b!��ͭCW(�K�0��Z-�����~� ֲdyV�:����V(�|�%�~��V8��If�y����������S,�����`�����?M��~0��d$���a� ��4-�9y&���=4a�}N �(d������Nv�^����b�C���񎬟����������	�\���vkŜ������H�Ǆ�=�����~�9�Sh;�V��J����&j?_a��8�Ø�% E��(��`YP��B}L^�NEg&�nc�V��Q\m�R�ŷT���	���E�?����L�(�>L{���R��΄������+m�6���d��ɦ�<dz����Fؐk��
�^��������s�:�Ҟ�+0���z��d-��n�n�Ie��*e�
�K���u$m����.� �q���^7&�����#Y��I\��Z!L��u�5cL�/��]̝��<� ��wi�H}e
e��n��_��+�%!)��[� ��dٍ�SF��Gɿ�9o.�>��c$|٭!/S��]�F��*vC�JI�	�صk�VQS��*����HܸS�p�|oBߨN�P�M.����p�fj����Z����3DP��0����ʓ�w�U��#��V�����B�%�G��+*���,
οπ�O���G%�A^j�׋vb6�H�/9���k}��jna�њ)�9��./#c�5��&M\Lt���96g�QaJ
L��%�^��!8�龘ZB�g���GB�%�9�{��κ�Hբ���8ti��%A�|9=�<��>s�6�ן� 6M�ⴲD���s`�YQ�����c�^��dOk��v�i���&_�OnZ�.SrbᦹFލ�$']��Al�@!���ǡ���봜������FV�'��������0/�w��"o����ڼyϳW|M��5s8m[��ɾPen諔�(&�K;i4L4��L�,������J~���M6��i�֧����}�Y�3�dV1 o���u����]!q�� �j.Tg=���=��d��p���g���1w���?NhU�l�����ќ�L�H����ڌ4�kϡˁ&��7�B�s8�@O��ّFޯ��:� =�-���:�z�$ɼ\��d��D_���B�Ml��%�r�'{�ԣfL�
�Y���K��NHRc#�2�ˡ���0����xtm朖����H�l~�|���p���IQ�r"S���N"�A~���i���oa�8�qz���p�͌���]fZ��1��.���d��gn���)d��Xa\ߤe��&a�L��"A�փFB �[�sda{�k����uЈ q`eG��VM���FQ�Fu��C�b��Έ�VFZή�bw_����e��M�"��e�;PZ�E��j�}��+�'W�-�J��
b1�[5#oK=�,#��*������+1�jzV�G����}��O��,+�%3���fŞu�����1ov���x�x�8p�������nV>��Q7#��89����]cX?eSw}��F�/��l�er']N�\�m������r�	B�7�F��q:EW��͛�]o���06�*Rb��,��iz��=_ZG�G�ٕ���N�޹�Ĝ�I�^�5�(l�a, rK�ø.����о�FZt��j��;%��p���]�ts�27nt�,����
V����:�m��*����F�@,]7����}u�����j;�]���m׆��Ɉrl�QU�����O����o]T
6�j�49Wd6;�Q�J�?�.{�Ű�+�Sjˠ �/�/��?&j,&��W����6i�E���s�X�ŀ�9sg<����S�Ӂ�����F���/���Qc��v��R���}�����g#�8tk�$����f��8"�r@�>'<��;�u�@pC�@�^�
�K�ls�(����$������M�,T��ϰ�zϲ�ȇ��L���ƀ;b���%�g��Y���f�]��[Q�-��1�U�EQL6��(�թfU���T���\kdb��ͻ���LS(J)5�w���J���n����6M!�=��w�#Y����j����^��?�:J�a7���e0�m�H����{�R�����f��;S*���ef�����?��	���75 s�x_c�ݯ���>�G�;Oy#��|F��j�lf�{�ύ���puˉd\�lSwǋ��I�����"RF�/6�F��ps|��d��#i��H��-���DGq�����Q�JN%�L;�S����ڔ�%ǣ�+,6��:���w	��E������?R`����%�c�uĀ��+N6�4��9�T�������7�V�_5Vo>,"���2�ߘ�N�������"�SQ\��N�MV�LrG��/�Ͳ"WS䂀+���by/�T��=;��Ks��m����t�-6z���7?�e$�����/���>E_�k������5���}j@�������A߉E=�X'����j2442�I��I##����a#�<-<M���l��F���'g&�F Q������O.Pi�^�)Mut�A��޾L(_�kV���ylyF�qi���<=-�O�R�/�U)&F�����$u��x��Ɣ,����0��R�v#��CϘ���`�xJщ.��RO_��N��V 0���2��dY��Vj�ڥ��������+��j���R�ȭPYn�'d*S�.�[�R�&���=���P��ص�cOc��dP_Y����e,��93����?^�s���|>�����<�9g2_W�2CB�l8�o �]��b|�9�zŠZ;�'�hͻj/���3�~��^[ ��N��.B���Y6b��̥|�8�S���&ùd
U\�%��bE�D*�c���M?֏ B�X��)-�0���M�Ȭ��;�ڙT�J�d"7����jޯ��S]�w1�GG:���)?�2]�*��������`I@�лf���+[�<��B)���ܢ����Q�r^+j"�𷠹Xm���(��$!�+bI)������(j�k���46w�_�B��A��r�\d�q��Q?&�s �6��n��D4��Q�Ws)1��X'򤨅�+�
8t�[ӫ�SXb���������@UX'5�w0C�p�G А�ZE*F�������a]� ������^��q��p�.���	����6o��D[B�m�掉Y���k���5�z0uM���9eG��H�a��l���ޥ��j����a���'do�R?_���˾T ��韜{�OV���TM%C�(���x�ݰ6�$Ѓ�Z{��8�(�>�ܨ�Li��jP��[}�r�Pڸ���;/�,]��>Fn��
��?����_"��
H�f��?_�~*Ew�fFa�1����L�U�8���I�R=R�1@k������S�׹�?J
Lj-G�������������Z�:���FB�0� ������2TZ�փ�i���s��.KͿ.%fS��\~ig�\� �[���n�Yx��$�3��m�& ��D&C\M����f��|�)wZ;�a�Y\:/����ї��f�x�X�+�i����B����N�z��1{ �_���w�8��0�ެ�#�A�L��g����.�տ4j�oٔ1�u>��|���ɧ�e�?�kdeK	i��֪Ň���0%礴V��P��Ai�:rQ�?��hX-YC~�
Z4b�����2�)	o+(i��|��a�e0�<]��c}U�8o��\c>Wؼ ��oh�t �|�	���O)Fc3瀫�}+���,C�V���]�6pV�Tc�E2o���a�֭Y�$�t���/�l����'�ᗀ�S��ѶoX5Av�����ǒ᪷���?�\�� �F�j5���3r�!����"�#V<�\c�����X�\�gN]�V� ���s�����tpV��Ӫ�%�\շ��[N���(t쿙A,A�y�h>,֣��*4��1
�?����!$-3����xP�~a~�&΢��#����pb��q��3�N��f�����9}��<��DKA��(��]\j�����!��ak�]BL^�z ����CQ9SCg^���<�7�J�H�=��|4��,��d��� ��7�գ�Μ�y�u�J?1�`L�M��=&_F�2����\TV���Z�\Yˀ��A��j�9��9e�"8[�Y �D�M���f��`�:}Z��Wr|lq�$)���s2�φ@�n,���R�$N,sѓ�@�4e�E�??����*
|r*G_mīڇ���꒙�t��	���M���<�ɪ�f�jf��&��Cq�z,#M�0cMd0��P�%�4i���O�	�A+á���@����O�0�@����gA�}�������Z��s�a�$k�'��vJ~c���rݵ����DK�|�]v����d�� ��@���9[�"�0��S�|=�. ˑZ�pM��(szq�.�F:�\�&2��EZR�-�,���$�?H�SǀS�"�M�\��6��!�)�E��5a�L0���u��t�įP6F�
=bw�� �m0�~�-���ڧZ8���v0��w������@i��~z��se���J=Ȇ������, T_җd���Ϝ�MцCndH��#�Cm�V��)�>��dU`x&��{G���g/��E3�f3�D�$�9xڬ���F�Zm貦.O���	�b}
3�km@`��DG[�$x���#$����y�P�E�[8��Z�_�|��b���-
��`}1ZC���aH<������F3�Y�_W^<��rȚ�JK���m?��6�_%_��6��Q,w`o��l���6b�x�:�y(�G�2�q�U�l��u$����|�:Փ�Ű �(��U��$NS��+���]��N�XNX�k��9�d�a�=}���tvB%6C߰�B��0`�9lr��#-��[�b����x�(#g����=�m����k����s�/!��9 p��t'��d�7-�2�6j�!���
�#{5��ĕe����O�G?��4Aƥ޶pF�߲r�3�9�E_���@A��0c�-����(��=����oQ�ɩwJ�{+y'yAAJ�Z�Yz�~��K@�@���{fЄ=&g���3�~��Ф�\5��uk���h�G©>Y'�Ճ�=?&��)�D���.�(-�{�Y�? �2�`����k�3�q��Dӟ��|vs�gx�)|l�� } ��������-]7��,G��G܇�MY ;r�l��כhEb|;�b�\����)!��jKoZ��O?�u(9`�o���w�J{��_���La���CO�r�g���뫺9m�� ���K ���|d�ˈȴ���}����4�ǋ�vEU�FNj�U}S$9�(����Yf��v�_$Y�&����2c�׭?�/ k���:�{�K�k��S	�H��=	�8�w���B  �h����b���'M�*YK}U�B)����z̆�	4@�#Q�M \}�r�غ�]�W��!-�ӥ?9i�	\Gn���s%�X�M�}RV���6#	�)��0�X��Db�M�eΠ�*��� ��xr�����ksx�id�����K�j��;���Aw�i�=��9����^�7+��ٖț��Ҷ#����P�3��B��?_~��4X�;��k�H��D@�q �� �:�UVN �a�M�23�6IS35����ֆ���W��%���\���
�V�Y� �Z��YN���Y�!�l��쫵��D���[@�-V!��H)�J��YZ۷V-��ؐ3l��̩���V�,4�P������0�C>�Ӿ	��$`#wP=�cy���
�-��۰���澯wҦ�?9�S$����p���%jb�У�K�Z�͋����G�{�r�g#X�d!�7��$0�D���KK��]����7�,�� ��<��O]�>�p�`��.9q~e�L�+)��B��O��z�����>${�ݪ��rĦ�}�:�iZ��X5"fK��2�n�oWz^h�Ð�t�
v+��	��9C�{��Z	��	6�/����7:϶d�BGc1'�p.݄Ο�n�]�[���*?A�dx�����8�LT�@<��i����f��H_������$rIx�1��k��Vh��#�<�@��{�8��}�����(S�qp?�(ѕÒJb��}sף�F�8&��E`B>
�i�^1�K���a����S�?8���t�u2�M��"�z@�_�� j7,n�t����$�t)Rq��9";�2��[;Y#����i``��^�<g�R�2K��	�<�y
K�G�E��u��~� ��i��61u��:�v���ם�r�D��[��/l� ����b���+�'���d�n���}H��1)FTׁ��<�FQ?{��i�����g0����� y��f���pW��<�P_C,(_7�·�SY����\���	�{q�}X�
����!�kabͺ���v s�Ь. \�ՙn+�kJ����
���;1��X�vԎ��\�M�4�`?�El�wW-(:��T�?A"�m�������6�ΐ��.�{�y^��d�$m)<���bV�n�����W�t������#R�
zu����,��,���1ޕu0��l[@d4=�h����z���P�i��e)���;G��at��^[m��cW�kq��mZ^蝄�<b��t����\4�G�y�Z��b������*uy[�Y��?K�DS"���P�eM��>.��oV�Ꙁ+�H��i*��@��ϔ=��B�q��<��I�v֗��:g-��y*���U[k>�.�V��̑�]��U{X�> ϱw�.~��ŗ�2����E�.N��Jv\���(��5mn�T?	��b`�&D P����Ta�Ȕ��^��Z8DՂ����^��ΡT����:3LxG��g���Y�~SB�P
��p1��w�sL���i��5�> ����J��/QM}������Mln�-������o��b��D���������Җۄ���J1�91�&/�S
�Y�·[;���j+����C���t�cz� S���.�����Q�%|�z�@WV��~C�œ��!NC��0�GY!�C^��_K�a�]�� ��*��J�3�R)>=�,>�s��a��6��f��ne��0G��(�^� Xc3��Hb=��Nd?��+��"�Z��Sr2���ć�q,xB�!���38�.�R-I�-(���g��4_*R���S�����Ю[��=K$p���eBa�)7�\(n���o�i���hi^�ILN�)@>��z��~k�2�����U/B�4�@.�'��˖8��$]���� �PIt���V�9���~������NΊ�LU��I[*�SN�K��N�C �j��N h#f�FL�Edi9���ޥ
˨:�@��ҭ�j�fj�S���B.����6��ץul������b��76x��r��P~.zL���A+ٛ���/e�_�U�綱p����\9V�Ҝ���4�m'\�%u����'���!o/j\����ÿoy���^My��G_d8h;�o���-���"ʚ8����'�&T�&�MI��9��`�ޡ�%ʸт�S��>��bE��;�C>����1�d2V�=.|4�-f�\� &�xʕ$��D�N|�����*�zj��?l`�~�Z��EȜi�/�� '^�;H��Eќ��/�UZ���7S�S�����{�ظh���Q�����˫1��}���K\��?�,�:*eM��!-R�%�nW2[�!���������B��T�yl� -��e�-��m��瑚Ѷ�UCh�
�3&�Cv~W�E_���ު񱓸��cp��.É�� �b��r�}�,�V�7�~WYխNei�]��ӣ:�lI&�X�J������ǵmЇ��;A��<�.��Q����Yd�:�
�%3��m@�yCغ7��㧱��2��lCC���R`V�w����BB�9�􀇗χ�`���՞�g=��kxn}᪤|t�Y����dAvI���g�ݮ�*h��
�7�>X$�3ະ8P��vi��(�LK�����ھ���W\F8��p�Np#��AwC��sĴ��j����q�I�E��:z�>����FHb�n�GS��y�E�R�t�J����O���Zb����p�Y ��o�7՟���yr�p 8�)�p�$��3���N�a�~z?����K�-��������x�w��V������񌚼�.����f����PK�X* ��0jwA��b��
M�C�J������3ป�*.�Y0oY@�u�٠�4��$X���G'��Y{(⋢:p��3%�^��Nf�v�z�P��A��"�l'lE�;��Jē��|s)��\��9n���_f^$zs�G,߽d�hR�9$�3��Ch���-���-�����gb�a�K�eee���d��ץd`��[�I;��`� �}O� ��HFx{f��\�\-'���k�佷�x��0^�#�ֆB�vtt\���v�x�4�W���F\���j���k"HST�	���\M$���~��vq�+%w?[a��d��%V9w(m;B��/�Q9D���YfU$yi�eX���hP$è����ג⊊�fX$��V:Û򂮜����<P�
�,G�/`q	|�̟��~X�,�JL��rA��چ������J|b
m��H�e���t ��K���?��6��~�K���3�@+)��f��%��G�C{�A���$sd�]f�%]JJ�R�SOi��q�ȇq�!��qP�i�_���ȼ��h���88���-28��z�6b���+�XB �ўJ��͒>�w1��e����q� 7�wZ�e��)P+STTb�����Ҕ� ��.쬝΢0�߈qUڝ�2r ���Ӏ�]��@	�l��\��~�,��k�M�;7db�kZZZػҟ�.Nld+�3r �Y�_�R��>� ��ޗҳ>i���V��Va�1D�E0�kϭ��a�����EC� 4���DE�A#奂v�J�a�ڤ�U�3����x�К"���rに�srk͈����y�P�aH}k3π��S��
���{E'��t��_C�Q�g]9�\J`��G�ť��lL����r%,�9U�����͏����U�M�]��#�1܆ϓ�8���6�:�FM���@�Ȧ��K���>��7,��?Ö�,�1��[OU+VN�)?�$p.�q,��U������P�����,�9�������:��E)�N[��=�K�|��C��uL#,�����z�f� ]�PФI�0�']�ʹ�e�g��z=;�ٸ��Z QhB/i���<{����������hd��0����9�����*辪�j�ӏ�|1���Ɗ��T��� �k�Mi�z9]K��}πG�RR7�	�㭹����ˮC3��άUY�%� ��)���;ef]b�?���2	�����6A�����>*%+�֍�j|�y��Hܣ>)�3�Pf%��JSo�~T� <�=W���j,`�Q��� "E��(˅8�`bb��3޶w��J�6���c`��^?^�);qV`]�;���M�p"�� ��[��@���ʡ!{~�;	�:�/l�{䇟�[�Z���Es=_���{�=�րᯏ�zP?�SA��d�*�>��"[�7�^��%=�<D���k�������"� �[��%�Ƭb[�,�7��U~s
�P2K9[}V�wƛ���+�6�M���+2�|��M�ڵoƊ��4K����IY��X�P�|���Cc|m\��2��5Rzn<1�/:_�(A�AN����K5�r���z�#e��b���\Ȉ�]�fK����a)ω�iLi�Iݦ�Ȩ����Y����n��4?��U�5d���N�W��UĞ��&'�p�+��D�GC� ��q
i�%F���ٰ�z6�'���B5�Ĺ5��W�3԰�,h�w��e�c~'�����"_1��.�'�����	�
�^к��c��d����OQ)Y��sb"��7�Ŏ7���Sn� $���e�yVh���IÔL�����(8l,w��X�ΗF��u
���q@NG�w!�g����l�z��^O�3�{c�<�N}�e!�U"�nZ� �giK��1Il:o��3K���Ok�=C�آ~¼ҾT�8f�:�M�(z�mL�� ��bJ$�$u�`��M���Q�g�k���2�g[��6�ǥ�2��p��[���%&����w~�B{=�&-��N��f���Y�m��s��$a������x]����(z	_���jϙ�:����BM��-n�I��#�G�`�6�z ��f��؜������(��.��1 ���Ng䅣�3G�D��A���'1��Ǔ�'���
iU�YJO@Z�נ�*��,�X.�MR����=6�f/o]P���8K,;�����H���=87ϓ�48��d3�
�\Z��V�E��<���Ѡ.����5SWF�՛�ڋ���oa6ܨ������ނ�ٮ�M���?E��Oʭ��0{o��:A(�O�*[���7_��,X��DȧB�w`H�K�R7ΰ�����m�f�ΐFjir_h��w��.�����=���TjZ���%�)�)١�����kJ]|=v$�"�t�.�B���(�d6�q�ɦ�0�'_��[�X�����k	��S1��n}W�X�֐���>��ڑ�W6��K!H�x�N��|��̰�jf����q�C�`����w8vSQ1]��+J4����:�^� @B��xX�>�O��8,B
89�nS;i���k8V~���[P�GGG�0��Č��a�E�<b=h�$���>E1$�%[��s�S�v���}q�5��܈�J�R�ܐ���$��e"H�-Ѵ�5�!�~����*}~��F��(9RӔ%���!��.�VT)`��_�V�����/I�7�b��a@�;o�?V���<���������l�Ѥm�1&�~`idd$�*iP&�E�cAJ�����U�<����� �`��tZ���z�U�8�Ջ^����/�=�	<˩x��T3 ��N�k���G�^�_kB{z�h�FD ����~��,���A[̈́s��J죀YX�pa�Z���U���d�N-l½a݆���7$�B��'v$����x�!��Hn�If>���Xgs��%o}��"p� �,2=5��s���s�%�)�#�rW��Q�����z��)�b�Y��>x>Z)��7G�y{F�ft��złA���BP2bޒY���& ����@���$Y��r�	���V|��F�n%��B��t��$@#��#-���0���v�?=��c*q7S��=��qR���O ��n�X��ϮZ
 8/���j�k�`��!���Ub�:�ښ��TOϜ��+���SF�.���.�a��(H���+�~�9M�7�Y�BMRRU3�Dce�>�RRcaշ/��봣����N�r4,���D���><�l#��9�Ÿ�]�4���T˘����
y{��T��>���/Q]���F�-B.B�NSKl�DP��`C� �ч@l��ǳGǹ��}��齾3zL����{��>E�}q�,53��y"���3\=���������x�A�}c��?�k{�s�ob�f����
'�#�%���b��7㑟�^>!��PS�j4|^d���Ic�J�@�x�L�����<�0���j�Q��5��^`H�MQ&��4�!����O���"�ow��4���q�e��m=�aV���W��$z��<�.&�UJ"iOVti�/�����8?�1�2�4�j�jW[��lDr�䀈`�1�/���&9%3IX�
簫�X��i�Y�qx��G����.�y`��g�{S�e�
Jr�5�>�#�җ�NƜ��2���'�
�(�u�;d�~����m�ˌ�b�	]}�!� ��t�ϗ9�9�gv28���Jf�r�����c�O���}u蠗t��!3^KH�os0?��*���Z���H�&=9tUFx��mUxj����j��j����kϮ¬����>�)@����Ƅ�s&+XL]�K��Ģ�\ϒ�F�ӏB
@�bN��Y�#e�pR��I'(��fr	ܛ�K��[yثT����d��}�lِ�O�x����3��;����888(�q���^�5��(*Z{�.Q��L��v�������F��@N؁f���\�%�|*v.���rD}�PɌfPH�{�Z�+��,��і�>���Ȱ�mmmOa�3�ᦑ����IGE,8�B�a��c&�ډՂ�:�\�H.�{F��%l�K\O�+���d��ؓ�Q�T�q���SlI����A�!ۤ�u,�"�˓Wr�;�a�^�,H��M�U(��ݰ��:�����F7>���&��ʿ@��L9
j;vBK����͢�cW�|��	���{�_�y��̜=pc��� �8���8o����%�`�f��{�����a܌�T�P�&�u?{����cb];�	�J,�X�����$��	��iry��.+*)�Sҽ�֠Rŉ���DX�7��pQ�J��$(a�-�r�>Q9�o�K��o�����BAk͵�� ���9��~Mj��R�D�S�4����ˬ����G��R��6)� ���5�����ƛ3����`<�V�u<3i,�ڵ�"خ�.�
��-��>W�ڤ�6ň&G�M	�g�M?�C~�U/I����Gy"웽۔i�;��wן�L���Tg+��A������UMu������f/�dH䣝��~�lE�9����d������I��ڧ�N�*�|�;[=c!J��x���	E'*PG��U�}���C%������k�%���j�)#e�SUS�x���y��Cu��'� . �0��;�fĥt���Z|����oR�mU��C��7"H��
X�exݞئ�J7��H����}G�᳣��a>�h��WD���i�@�����@�ދ�	x����kg2c�n���6�q���
z�������n���5?�wǙ�ҍX���W��V)��z�՘
,
���%�U��:���`fcס�l9a�j�5T`?
�W��+R�%�K �N��(]Wr�*W�]�Ӳ�<7�E�Ԝ������ �)�		eNa?�h����M6G��k}� ��n��pn�u��x:-o��ްc���B�d�Uw/�`�'�>#H��Wb�sJT穽sssE111j]���l���ۤղP�'}��������4`�,��{߬7���+m�<u�1��T��q���VH�?jP�̯�;z@�%E~f �V�+-��G���^�zT8��Drf�O��sF���'�D�Ϡ�߻<�}Ɨ&t5��x�I:Y�/�^綆>2�8�;4�i��ſ{����P͝l�\�(�˅�/%�� �
pA<�����p���&j�x��˫�!��&J�q���.o��.t,]Xdu�?�w�*h��Q�[�����3[�N���a��w�w�sm���ܴH�k���4fc����9��Їq��1�S׀㚺��|� s��\BdK<_I̟��F?��r8u?8@.��]]�3����
ٌf��<���ޘ
�k����,�߼�ؙ�}[�e�G��ӗ���B�h��!ޛ���eH���;~R�9�%#A��|[�&q,j�~yр���w�|J�� ��������2
��bJ�u��;���>��=?�{	�oW����
������^�o���G����08K4}M|���UPo �J�נ!cA��g׺Oչ�h��-��|���B�Qܓ�ځ���i������vx��m��I���*f|��D?1W~�W@5�vdr(jW1�E�=�k��s71�` ���D��D�|E��P��d����Q�$�j)�+ӗ�?ÚN>�:�,��H�<��v�w��.N,�H������Z��V�
yNOѽ�z��S�Ntc��x0@<H�J&%wYsEtf2��ۅ����dK�
)!^W�����	^�PF;�?�׳U=���m؏g��v�5�w�|A�����1d�*R_U����<�c8;�vCl�ގ�\�����o�H,M�`ŭH ��RF����:�N�!8reen����;sd/.���a�J�v%��� �w`,>�e�����y�Z�����@�G����N�H�2��Gy�(�
�!��Eu���e���3��0�.@SR���@������Fg��N*���$���}HO%|��W�NʜQc�� )����Ǐ�V�HZ�#�QO�1I��A�� M�M�O*�Y6��?VH��G�Jb� Z_�(J��'����n��G
[� 3/�j����;+	!�
[��B֟�:�%�}U��
�l3�f�*�(�|x�̋�Ê�y^A���'��P�?!�xy�(߁#}ԅ�2-D��c�X����$�>��r!��~ N�҇O�C@x�C�xͿ�g<ƀ�2K�x>�骽�(Yܹ�>��gb�^Y���0Ot6eWm�gس��u��잛\J��@M�1���
�M��д��*.�Uz�@�;Н��ff��pZw26�g�7���[��1�SR���j|B&������/��p"��*������//�g���x�K�+*sK�b{�y8NI)F����W�7��c�v��� н*�u�����r/`tw��;(2���hVkԩ|m��>�?��>E-��<�> �F�Qi�|�
v@�w���P6%2�B����;Mps���N�h���%Ǭ��r�ĆX<�#����\:�𽦀����='�ۄ��~0>E�Ja.�D�W���7��J8������G޲=@�wZjs���N_E�!bC^p��<�5J�L&S�{ei{@H�	�"�*��٫,�KX����h��Ő��̰_�M�Gu��>��1�)��NQ<PNޠ�c�"��y�xuwbt�UP3�ٔ\ӟ	�u C���0�ί[��i�����Rk���Z{�4������G��J��w�~:�f�����%.N$a����l���B$_�,�	XF��	Y�R`����(�� Wq���_�ʡ�K7!��N!����Sv�O�H�]�%,����`�&�xx�����F�B�(Ȅ4)���~��f�A˿Ïa��5ԷCP�S��2P�2`�Yj� ����G��j"�jR�|�ry)�\�"àEA*�,��
�} �����*S �*o�bO��� ��c����\[�߇!ͰS>�,�J�����W��Id�i��u^GH
^��?���$�m����4�՘�斸��N��k���!�5�m��'��81���Q?>4$��p�`��:��6�*!l}7�Qz��t����R����8��9�Y�P[�o�[Y9&I끯g�F�ID�_�SO w7͘������%�p\��!n�=>)���M�L��%�� >����C�����������Ѡ�������(��_��R@��3��r#;FC�gi�#
��P���o�}�j��"R%ol=�Qi��H!<&0ï������I..�h�CH )�֛��c�r��CJ=�luM.	��D�C�l�OL���,����Qw `P�.�ߧ�\v�5?��j?`����E�@�~���O~�ɲ�v4߽��֜eӆI�c��9,�A�7�G�������ܐ���S�Г8���OcE���ܹ��>� #������FA�� �QT���!g�D/h��Z�%�|6�9��6ZYA����K�����X5^���s�>���E׆�C�ۻ�A5�{�m�M:�W^R<:����8�����hE%dz&�%=��B���v2u3�i�TGa�9t"�;��4�L
��4V^�mA=d��п>�cA9t���N���2)��&�|L���y�.T��il[�����t�G1|�����5,]���s��x��b�!�sӻY�Dg��O�!d��E���!��o�烾vJ؆~��f���6ĝ:w�'�n���!����N��@^iL�&���UYޮ�E�/�*΢�ubo��n��Q���H�fd�t2!�8��������4L�.�V�xR����YEI�B.��8��C~3`�̾����R���RD��0�E�sֳ����y�Ri��Xj�mwOO����J�gC�@�؇��}�������i��_������f�׾~£�a����(����q3	� �z�1�l��J;x՞"{�o?1Qv�w�����	�+��8rs�n��+���5Un���M7!k���!<^���ċ��V�t1���,��YB9t�%>�D<|"OPG��s4Z(�PNC�PZ�;1��k��bib�߾�%�f2�����UI����Z[ZZ�:\� �:��4qK�V�-9RZ ��&,�;wN�|�����{�*�bBi�ӳ�=vt.��Sn�Jn_��F���M3N�1��
쏅=�T�����g�������v��u��Z�J�9%�p���	$�c���\������;|o����F���jY[[��?�^���fjb�pʫ*�{E���o��옷g����Y�'���O�.����}��0� �8�t����ɬ�X17��&��Q�,���R((�ɑ����O��eeKx$?4	�W���E;��{��pM��xm?�\����:��>�we܌�*�x��VVO��T0�	8y���\qbbbe.�o�> >��
��I'�;|�[�$�X0ϩ��k��z\JX(�ap�D���M�[��V��jqtҭ�oC��]K����������j��R��D%�4�À�sp`�א�7��\d�]SWw��j�%+�ؕ�q/Y0O	A�HP������OԷǥ���I�Hz�%��5�h���*~L�=�!�,�A��}�;~U���W�?m�
�����)�@��x_ �?=�-!E����'!6JY^A2�	���dX�R��!$��nD�O����a���}��0����ƃf�@Sj��x0Qk}5�QB��%j3kN1�R^\}�"�I�p`�� �*�@\��'���_��-)ᩘKo��$4` ; @&p���.�z��(��@���{���-�7�j���+:���ÇUٽpڜ�M�֜��`�N�-�j���d�Pj8� ��`�/��a̯�&�������fC"���J(w����������*y-����d�'�}y����@}��������7��ڡB���X��'*jI!80h���9�3�l���*��?@���K��*�q>~��0]�ꓭO�w	��΄7J�7<?���eO;����@��)Vu��m߫�[@����NS��U��;�4���%��.9%nO��)��&O2>����j�_�� ��]>�ܕ�M��T�q1����
�$�V �&�Ŝݞ����_<�;�;�)����jN+���M��7z���.N��V~P��哛Vs� %g�#J\���IpI�2�;�֎t��Z��-v;��}	>s��l�nHopXs�_�#�/�~)�����,or�'����m8鋟Y�i�����������y�ж��{�5��?�Nw�Q����-���h�v�p�_�Q��@�M��c��?��Pt+��\��������c�
�/i)ߍ���٥;�&������SJ/�MR�t	�7�WV����s��:��+pf���K��.�8_������|lg0�m����к�_-�7|�R�&�:�ۖ^+�TmSK=���H~��������\\�n+�Y���ĕ}LL;��S�t���]����L1���&V�hM`y�oʙQ�Wb�>˿�Nr��PcS�) ���]�)��s>�&.D���	�����i�.�Ja�4xݸ�Z�۷��o�O������ŷ��ʦܮG�>��0*�U�^g��a��n�:t�6(xk؁b�*�p��z��%��`�2��B���u-}��ZnzyW���O�5o����~��H*���N�s[��C��	
�ޝ�^�뵁���|��p��R������y��Z��o��w4&:z��䭖4�f�<hʣ�'�ݼW��[Fz�餯I����'�!=uHW��[I�c�g�mBI-����b&�/o�4����r�w%�q���w3����t�[`�⎬n��%�VH��N��J�{Y���O��6VD�(@z\���b�f��ү��o��K����@�F�����y8aSgI������R|��)�`�s��G���8�yr��y�9'��t�6���N�Mu^ʅ��;;�k�TYBm����vu���/V�oQ�D"�V��<�P2��4q����io���/-����þ�9���v��w��yn�̬�T�s4K�s���|]g��j��Э�;'�w�0�<Vz��)H7h���/��35��j�de�ZU�/�v8�o�w{$4b%/��i�;ׂyYd��+G:��y��碯��|#}�%�G`���w�v���<V2N���2����Mccc�U.�HV�W�k߱���{��T}�gaч��Q�kd쳯��K�-�����}�RK1�"����XA�D��q������N����|�tb��ܴW������9
�yTn�X���J�q��
k��@�?�pN����;l�h0�M�V��uv'�hQY�>�?�X��iz��%��?m}Bm���}"iT�����\��Y���2��Ƌ�'X������{1�Ҭ��fh��*�y��%�^XYYI}��G4���AX�랿�k;�Z�5޴ggx텈���r:�g�%�1-�e�r+��ǥ����h]xF*�]�4<�.+''�^�������ź�+�������L�W�K����+ߜ������>K�^+���h]���Ja �rr����<-sAeȁ�r���*m��XX�8���}n��%�F9`��c]�l����9�>�3���d2��VV��m� ����׾�nv���o^�M$�0��ٽ�r�L��Y����� �(�Fɱ9��	�륍�����5�=H%E��$ge�|�k��?�; doǏ�1����{�,��ݹs����>n���l5��󵶳��Sͪ����/�)?��>`y)�2~6�{��/�|V"_$��A�r׎)��P��am�yQ�7ͺjTq�䗄�A�w%���@��f��S��!=�N���B-�om�6n~&��Qf��k�w���;�Vs�� ��k����n���@���ҡ|R��o��{����_��]]������E�M�qi}���cx�]}�q[��� ���t��o��쾛���M �\��v�����`dd��������[䵛{}d�o�w���k��Φ�@��]�\c;�>�(TZu�]�j�O{���B�fE���M��7�#^��>�X�qǍNM9�z��������g�o��J�o,H�< w�색�j�b�B�%��P|Kw�gC���B�����	�RI�a�#�<_n���<���"��I�F���\\!�����5]�!�f�|nTh[���-96�Na��nUUT4�v��I�l���p���L%�l�����o�H�i�R�p;��oGt����F��v��wX �[z��'�_z�����)�G`��P?��i�X�x�j��v�f��U̥ٽ����uY�rRT@����V��\,]�t�]�qO�Y\Z(����n49��x�>/�7��y��0E�z�ݟ�?�-��0�~��]x����)@�q�Ϯ���vT8�]W����,�$�84���㲒�^y�h�6kI�ke�p�;o���#���a�4���k�Q�ht�����eSDˆ.����x��G��&�u��B7�P{��,&�[�B���0xpCCdܠ��B��w���#�ϥ�Hy4ix����Z�<옱��?�ˤj@A��GU�@��mHgxvtekG,�^Z�J����DO���׽��`�^F/�$^�T���A�۷�b�M��P5�ɰ���.������
�'�2~�Q<g�b���j�j��]��mz��|�KL7��0��Iކ�
oo<>7�X rɻ=I���{>��W��M���a����T�x��5����j��c0��ݝh $7z������_�-h~l���$];JU��q���6��"d�߁�;ݸ��}t���ڏ02�����O}Q��/���kl'%�;2�1��.F�w!���)��4�`���{aӞ����~�xg�.����`A��ۧ����:lJU��"����B-Л�k�p8�䉮=��ɋD��+r�x.���o���S�\��=���>G�Z��?���@�T�MP��;��]�m�?h�73H�~|����Ŷ�J���Ax�R����N;���7� ��_����r���c��zdjjb�<���a�X�Z�v���I)��{k��e�A#��3!&�
b�l���(���;R@@�`~����9�R �M���J�wנ�
�2�:���:?�N��%�S_�u��9|����U}�����>JL$v��4}��A��c��j�~}c��Yug�ȁ
0�~͵Ϧ�3��_�
cFGh��d�=<<*F�&����휦|�Q��e�[E��ϴ�Z.�*xʼw�����<�s�״�}V:^�D��s�I��'����`�"h-fp��{��c\��O4P���eL���D]�M�*��NM;����]>p����HOʣ~1��nĉ��W���]�J� �@��~�T��7�&P�?��E��͕)ߘ�y�V���A�c�r��#���U'�\CAѮ�^c������Ai��{����@����*@��_� �m��nRD�î�6IZWIX�yE��s�b�Z[U����@O��T�C`R.� � #�|�F�BDg��c���EGs��� ����������~P�&{{{#1�9�@�x�|wbk�m>iӞa��"ݠ)�r%���I�a���-X���4��;�Oϛ��͸�-�8a��3D����|���Lk��X��R։����\MMM?&��$eBr��$][���3bo����d�_-//�z�f�-��ǻ�{���e��K)���|�"\�H���\���5<��� )7n1>�ip��Ӷ�e�1
0��,�䭥����=���ǺUz����D4�v⻤ݜ�Z�	�B=��ȱ�1ء��i)=���(�0��UC�U��C�3���k�����56�"��*s:��+����m�`���EwF�����Ǘg�+W0t�h���E�=��C)����7�N�5>ǧREs��,;4~I��O�TI1y���tM�~����e���G�����%�T�m��P�H2�
�� T2mlIi24)2�d�2l��D���XGE		�mI�2��L�6Ŧ��?k��������w��:�w=�}�ϻ޵��^-BZR�A�LTD�mS;zyМ&,_�)L )�bHQD��I�;�Z�L�
��I�o�ԓ#��}��d�3�([8Jg|Qa~)���3��S��Ī�L&�vtx�b� ��t�D�/��́P|�G\��J�l:\9��>��߫��BJ򗩊_hƋ�����zf�<�P~�5x9��I&�`�#`W.x��,��8?��l�A����լ�p�;-j����u�6i�&n*��O�lL���m'o�)r�L�� �Mc���t�=�=[�t���M�'� �H�ڻ]�ˉ�������֕��$�h_����Ҩ��e�tF1,xc"�E#wH��B͵���i��3	�$�!w�+� ��
;5����o@�S���7㷼�͆G�w�%}y'��ۻr�@�^|��c�k�`���f>���餜����pP�Vvgs�
F������}�V��~�]�p��Z��X�2��/�e�uZT���q39��l�� #.	�'Źԟ>O��?�����hu��)�d��W��������z:\�nͲ�E�x�I$p�dWy��ŀ7�:���]���ng�B�o���=g��^�|Z������=�+7	Ġ���-���IH�����݌��ȓ���ӫ�e�
h5���I�ze�b�u�t����;�����ga��Y�H�����\�*�I�)��_�J�&}U�U=Z���IA���� ��q)"%��5�t��a5t�z���0�F$C��|8����Sy�-�o��*~�A� Ì���N�0t����E���~�Rė/C"�;�8�m�<�-5�vi��y�}��+U�K��3��a\�FkS>����~uA�`���˗��Xw�t��Uw��/���{Q�C�5\�k��Z�+g���&��O=������e1z!s���/������r��S��S��yk�l~ߌ���d��v�-�l��0���,;4��u�O�r{����h۳q
]Gw�����`F�V#/%�4_��!䜢���E&���dݦ�C;As�]$}wtt\�~��}�լ�:P�oϨ����U�y'���w��&�b ��.�1K	r|mQ��
������|�÷!����޾B$}�D�@k[��Н[̞�K�����*9��l��q�n�N�n�iL9�W��˅D���p���C�6�3�Y�OMg��t���5^�|7\\�AO��ݻW�-��jˉ5��_�.���f������u��,����w�x�*�̷fQ&J&K����J��	1�O��WO{s�pn�g����Iߔ5^��M���y:44������m|��c�u&'��Y:�A_����aV�x���i�����ȏ�#�*�m���wOVF��Fۖ����L���;���y;3�+,:�]�5���a����gO"����R��S�\�K��*^ tv"/7�\TL��J� Z�AR*����?n��D�teGU��ג�@�[�P*#�����5�Զ��ȓK��-yj�C�K�J(��	}�����B�����g&��q�NTWx_���pi[$3/���H�̩]WJ�u��?3��Z7��`�Q��3�EPy�x=s;����l���Ձ]J�Y/٩.���K��a�����]!�F
G}(��X���H��7��ţ�GM�VT�|s��ן?c��@�<#n�'������79��=�[I�LLLnCR�>-Ss.�����M�:p-YqH�Q`��v
�8�b�c�]�JMA�&�쒗��ҮO����p�V{G�b��-[����}��9|b~��#�r22���>p�U����H_�@����MW=�z��,�hZ�kr�+��n\��u�O�8��T*�MV��j?�� �+��)��*vsf����r扬hW����-ggix�s탉B9#�{�i��o|��1���-��LS0d��S� ��|��M���)>>~�g1٨�3�:�E�i>�E?=N�x��?4f�͈��㋓�9lV�G�5�P�~��3���E���_��v����šai���1�1}���P��>ע�-}�4w���R}���L�o��(/�S�����|�~�&����3TS �7Z6�@��()*�m��Oݽrѯ���ԣ�����C&�Ĭ_��*�����/�yzz�N�4C/�7�;b]���^_���l�B>qo��;m���De�w:pv?�Ӣ��[b)�y�oHz?��J���=/�V�W�:ǰıv���5Ԗ�C��a"]���Oވ��Q���{�W����w�fR����xs������b3#I�S˹��r	��F��Y�N��j���h�������gB��eGrֈD722Z,@��~�d�jt*���͑LVB��3�b�Ƃ�;�V��� �;�>���)[�;)�XL��o�Ee힡=��[a�V]�%���|��� /���,(��a���_󅃓�J�S>}�+m/����π��k�G_�e6��:�;}>���F��j��s���G)GYi��N#&6
>��{�<"8Į����15���>Y�WTW�%tQ����﴿oM2�-G}�_�Ʃ)��a:ݯL�%2�k{�7����8�����E����dQXg�K�W05��[c�w���S�^��91z">�/j��}��c}�*�������h\/�����>�i�.C��[f�P٩=��?�Jk
�	z]|r!�^I5.W���Z�k�=xBӱy���Ƃ����'R�������>��\��*piJ=,��1qL�o>͈d\�59�G���/SG��p���E�����RT��-��Ȯ��h�?毠h�<��eA��@f��#�����H��%ޢ&8ufo�ay=���%R� HJ��֧�"1���s�(Z�Ow�m�;�{���c)�>N�EGb�?*M�U����1�������+�sWxcb�&������	sƿ��:�m�V&rؐ(��vi��%G�����*�_���¯��&��Cg�>t5�D�R��;;/Cyeg���|�y��S[I3��}�7�Jک!Q�$�X�d�yi{�-�t�M$���+8�!�8�͎N���9��(&��<�k>��,'/oι��*�������䳝����:~Tj�q���<�cv�(2,QϚ�4�5X��M�wJ$Q���M�ԟ1av	'w0l97�æ��Q�~:S����M�+kn���ʧ�R��.���݀�C������ː݉9���0������B�w�[��c���N�_�I~�G'+�l��\��x�r�Ʋ��q�7��{���v�'<�bD��Au;-d�X�n�����7hv	��|_�DI��!F�*�m���T�g9�Q��/�fH ���\Ԩ�m��?����)�-�RW��(���fF}��%ٮH.�&ek�,rg�Of�Nwб�����m��}xC�gH��CR�i��:Y�f,�#�g�'m9��}�^�^P?�=�y*A0K?�5uys`N��
+����jj�0*~���z�Qޓ/�S5np%�ŋ�wJc���q��΁��:��.�ɭ���ԓ��I��!��n��'��ɯ����e�#�?�hs�M�i	����i|�����7o�ddd����@��u(Kڡ�Evj��Ǻ��m
��v��U���tΑs~h/h!�R�:S:5���;�q(����yn�J)Q������s>D��h��X⏬p~2ğg~�|�Ľ��:��i�||x[GGJ4v��d�|u�'���W�1o��xo���FS��ʬ�,�Ƶ���Ԓؓ7����n~���#���i���R=>�z�q���ki�H�������&��boRu�t�+�Ή�&�Y�{e?�m�*P��e����g�T�-�͛�X�L�G �%�;��4�U��].ڙ��YqyiQUs����ii���R��#AKa�X�m`M�$��럾�1<�l���~�ț��Ҁ�@�侕�G����Bl)�]�����-ڋEńɲMؽ:���n0J������S�7��z�%بp�GO�۵�+�%n�?Lic_t�Y��N�$�'l&72�.WǾ�N��K����zdK98b��7�M����t:A1ث�����'��]���B���#��v�W�p��ˇ���t���5Je's쵼���Uu)�\���!�S�D�i� ;O���$��7^T�j�4g���ϼ_��>C��30�6U7D�˾K[��Ȧ�i���1��*�6^��#���4L-���kl=J%�9�  �4>�Hr�R����_���H����Ew���~��	���O������w!:'��"���L�,���U��ɒ��K �$_W�?A�5A�Y�#W�(����$�S<��M�XT�� *���5�.�8�r,�$�p���(�K^9����WA~++Z2��B���tG�+ڻ�9ө��锫#aW����PS/UZ.�,�h���V������OU���Ay�	�P�m�&D��=%�uuw/E�Wt.[�d;,Z��b��9D�y�������V�=T�m�ŋ�[q0\(iJ*y��D���P�E�f��8_���b�vb#kv�v
�xbfױɭ�j�����B��NY��,�$ߠ�^{�]���	�U}�(���>���C^^ L��x��{M�%��ɑJ3��e%���������x}Z���0�O����d�Sbs�DJ_تʮ<YZJ�@I�ݚ�A���^�L�R�M����E~H�W�
�V4���=�	�I���jI��6�_N�_�=M�'�+��:���̣X	U�����
[ZZ��)���½����� ���
���p��Š�d
��r��u`+�M�-YDGM��[TI��ꢷ�0��{�h	+E�/��3�%&&������Dl�K�4�7�q~��̓%� x��P��4�Ou�b�.�
��R���G�<����cK�=�.\�&�>&@ƴ��e�c�za���U۸��aZ��p�@KFu\�vB���3_�׸�ǹ���^���_"����RN ����·���$Z'yˁ4a�����1޶�C�mBgp9�^������p��҄�p�'��+�/_&�X=I�Eos�t�v�%��
Um*
�𱾾�<N�w�ce�ؙ,�}n:����3꾙���P����>��\�U�-��o/ٽ��[q�a�!��<iQKj���#ݽ�G=XLt9%x��$5�ϭ�e��Mid���B������p�,��Q�2y�.Z���K�;!�傴�s�v�=��t\\�J"L��BVJ��N<6�꧀�ɲ�DP�
OTvqy���U�.�?g����7��fCm	��Y	���O��+S������2xD�w���Ic�=��_�\8,���԰Sk��.N�u`��5�[f��,o��Ud�f�Z��I	� �g�2ݙ��3���]�-�4�gw��u=��]k,f����&���n'�	��� s�K���8u�su�B���#����CCC4r���>0J���c9;=9n$��)X���V���hO��=2�"γ֙�޾Ђ���''��M�C� d��xkb�}�,ࠇ"�P��;��=?m�f 6r��MX�J�DlK��֭[y���{o��'ҰV��vn$�]��B#��(�6 sL�^V9��~�������f_1Ά��H�h�{T�_H���o��� �]�܀z�r�����n!���gJX��Ӛ���o)x3��B�e��E�!m�m��4ՁoC��ˊ�(+���@yE�'��ow��=<e��t����ȵ����t�+\��_<k�M`�x���c0lx4�������	`��=ǿ�����`�y��E�������e*2,|�B)��8��p��a�H�雼>����P�%a��]���J��o���ydX��RW���̍��A�����ν��F1�x7<hL	F�Rz���i�:�p��ҹ�9�pt�x�r�0rq�G�\�#,�,��۫�6��I��n/�z�C�da�;M���-�mSCF�5�N�M
���ےdj>�(/M����c�m��D2�@{�!���[��n����;��2P��T����?;��	�|�ˏ-�U�/�4q�t�S�c�ɧ9��-H��u��Ҽ���Gg�u�ۼB�đGU�<�GV���%����Q�n�By��+�,�,��
Q=���>ӕ��y@����s��^����OU��na�V�~�E�Uʖ}�T�UTL��<�Fn�`6��;hοG�|�à��.���1'`حr�~��߄X�Hĩ��n�M��z:+�7/T��6��q�a�{��#)��DU�AP6 u�.qJ0δf?f=��{EQ�2,v�un�,����������x<ӿd��!��c?&F�7�z�*,U�n`W����vѯ�}��"g7���y��,�����~�MbqQ�����F^�;m� ��������VC�F1�����xE��U{A�D�mh�t]�����V�������0�@TΡÙEX}�mY�J�cX�XA��(f�<$���{�gBdIKޠ%³Xȸ��e`����q�N#��ڎN�PWaV'�c��j�Dӯ
�3�;U�W��66@Ex������z��`��*������`H��%���uV��Ug,�:���~���!B$���e��E7��NN�F�� KX�O5��mG70�j[��4��d��A��F*�t�~�h��޳׉��|t�tl�m���^|�XL��:,fZ��\������6c
J�(�ՙ�x����d�B�ϴ��/9}��DAц�aJiQ?�㭞\�A��{�z(R��<E�ր���"���H>��u||<�����@���D�@w���ė���;:�`��DrQ>����_�����ax�"{X��t��!OW�>�%$���/�+7� ��u�sh�����2LQ ;Q.��o�th!�\�$��yE_ۍ���M'tx+���rh�z���)�M��F1�D@���6�k�f]bIAA�r:)�iT*��7P�����X�wߩ��-�|��P3T�r);u^��~SnQ8[Z�����]lq[H��<����<I��%����*Y��^AUxҗ�'�F��R҈���8��&���7�ܼ��7�%�]�:`�����b~DЅ����E�� Pp1z�[�].7�g��#�����l`���i���.)�l��<MJ���ćXg��������[�C��Y*AA����[����}�,i�Z���{�y��ԗ$L����,��h �6	�(�=|iȥ�F Ф�	�HA�~Ɍ�q��eґ�*u��~�����G���'��UB�>�;�Y	��B߄7��a�wSL����ms@�	<�<�<��-%�a����|J��(�5S��X�����hC�U���+e�z�&�=�*�8�PJ��=#EA7Ja�E�~Z�F�0	��x�����7�,�)���N�� n�<��w!���s���W��uuum�+��JΙ&sn��,b�n}I57�_�w4T[�.���C�,|���_�D�+wz�*��Ȝ��R�4:����W�X�� �/�oP����,�i3j��U�;�Uړ	/�=�+W�Jڱs?N�5Ɩ�Z�W�!��I���mD�Y%��,��f�PGL=%�P�oO$(x���m��ᑜ*���9��:��	su��)m�ſ\��i��L��5���� �,�@ �jO�xiq�+�5�;Ɛ�^�(u� ����-	�������(jh�M�C�!7�V<��I"\�r�������I}��z�v�������}d��cVA���|�(��^jb|��H���T�%D�VqeQt·4�|N_2--�N�d�-�'�$y�pF�ʞ��q�nEI)44�@�3�}�4��6|��ڟ�(�T��D橻�m,�4t�w\W��@�!(���b�\Bݣ�t�6��#�Ԕ�W�a��+�0�wa���\�1~Ok^-�}i������ݡ�O)����bE3�>����=��Tʷ�������l���#�[Щ���r�x���{���"*��+dF�}#b@�Q�'���9)GUBLtb���Γw��c�8�JP�$F%�|���PҞ^'4�;̓F�������~\��T���
����R:�?�ڤ���%>#O2,�殍�v���+O��5?�υyh	/��w�_�[�⡛����Ax���(j�@��lP�[X�;=Ĕ.J�n��P!��v9X�u��W���1dh:Ἔ�g�3�[a�u�	`]��_���4)L��3���l#��/��A�m.ɂٸ�P�ɋ��h$�m|�i�v� �Α_�8���0ZQØz��N�9��1������?�1�TX����g�B<ǌ9�Pͤy%�d:`d���C��g4F֖�]3��/;��|n4��z�׽Y~N�]�/�(9��N9a��ԪƁd\���'����kV���J��z���/�$߶�4��"�m��@w�Kt�C�5����Mt$�=�	�Q�edd,_�������6��Ww��T��y�4�� �%޺�k��ш�m�f3q�b5����0��� KЖ�ہ��=С2��GI�,�l���A�w�igl�����}�#�s�D��N��"�M��.�`=��7��x�
|'��S�^	��VF�(���L-�*��}���r$��dJ%�vz=�����b�LZR5�p.�
���E���$�}�����-��O�a�Y���i�,���gf/{.�{2��<J���������R��Q
m�o6����+rؠ���(R�a-����������|�D��nD!��4��j�|!�\y����$P4�ps�p7Z��)�weee؛Pȅ��N�>f�h��M)�vp��Xi>{?���K�^�X����>�]����'�*�o�n�\�AE���K�9�R9f��~�pbG��gj�ccc�}222;�S��R��7h�pv�W�l�`�z ��=�B��(a�:��u�����͵7	�Sk
37��&�!��0��H��۷�Y�t1J{�W!�����ڨ�D�LU_{;	�z.dv.7�ibB�hZ�͛7!����LE�:���E�J���4�[J��w�����5�pvw���4ɐ~�4�b�k���N0�jJHK�e�j�0O}���e��4t�-)���(�d�m���![���s�e��P�uj�Nk��f��A�\{fwO�����T��Ƙ� ?6�c��G<,?	�2���CA��>����]�QMG����"^��
笠n'��������s�v�kz�j�fbb�s��H}$6�h���]�w^|e*ԙF_&�x�W�?�m~R�x�e���!���)������Wmb�F+���b��a3R��=������썞���L�d�$a��M�5�H�pq�v��LvjB$���Z��+��vTVU�>ݝ��>*�f�F����G�),zZ�ѷy.����AkX)�������|�~1�]���ߜE�#�w�,El�i ��<UX�zr:c��M��=i��2�7��!�顫��6m�������3�vF�m��U��5�
������w�X�>�,��&9��t�z�Ӵ3rg����vBfM0!-��i���&����J;�ƆJ�ƅ��;`VЋ���?	ݙ��6��}G�s�F܏�U\94��Z?K}a:#W+��Pu��b�٧����F���A�	s;����XI"�J�,`+�q�PT�d#42��³�&ub¯�?O)]�a�{�Z.�C��T�{��pl�����4� ��z��/M
���~��
���|�ֻ��� �l�)��]�._�Ltwu�NTr�tr���?+a��o��KVR��bҼ�?�z)eO6���V��Z����൫���� ��&i�If��.��C����f\Ϊv�	-��,X��J��XrD��6_@�:�M4�D�/\J2=�����K�u��s����X�6
�����������@=݄�B+0P:�z�R5�pu��c)�s����ˉ��G�m��~f�Ni�v��#S��T�$�zL�6�� �U�7�dfMMM㚫����T�9��Wz�x2�)��]�����V@��%֢K� �ǀB�
���՝�K�ma�b%�}
&��s�0M朡n��| ��>}�777��V�Aq���&��Ǐ~�Y]�n�6�.����BQM��Ho�N��}	]l�@Y�]]��xY��5`N*�-�����e#�� u��A���`K����4v�K���F��*�����D��˂��g}���x��m��@ꈻ���E:�"�'a��S����$�y�8n���Bk�u��1�դg�?̫��%U�}r*��X�ø��Bu��F1!0*���3~c8c��A��=��>::����/qu��X��y:ő��O���? 09.�����<t�����gyB��G��>u����N��,�*�N���KT�g�3T-�g��������W��L&���=4D�}�.����S���0*�A�O����|Y�W��f�Y�C/s��AVEV]Q޺���-̜>)�J{�#��_'�:�uv�nnI��;�hc�����s�'����� M_Q��6G�����2�-"��S�oa�ܽ�'�xP��[]��@��9��W{��LI���&����b��3	���wї�O���۹O��ߝ�{U�R����:�sϰ �7~m�_��n�X���i&�}Qi��R����XD?���y] �g`q$������8�(�>�u��aŬ��F��+�}R��`̍�0Ѕ6O�����իG��*_T2P�S[0�� ��m����vM��g�N�ڗ�����5K�4���r�k�t���6�z ��_�JY���i�)pM���Bۑ�nV�y��e,O�������,�n#z��Dk,�.*��io��̓�'T ��Z�F\�Α�Y��}A���?��5�g�����G���>&?�/y��{I�nC_K�C���m� ��wyys�����@oqIl%Y��'�I,H�w�9V�∪�O�^����\�}���G���t�0��)(�6`o�Em��Y�f����Nx�����4D���
�!�|��F{/*�[A`��+�#
}&��o8�?Ν��܆v;�ura����j C(�1�K�$�$�UzF�7���HF�0�(5�-�%فn4fz�mR��v����C!A��m����`��+�Ϟp'�Jt��
�d�ީ��?�����6
��l��Qj~�'�'�u�>�9��i7��O~-[X|�:b���Lz����7Bm}�J[uu�#�vB�0`��ގm."<A�����E��^��S=N�ߜ�I�fY�$�h�Vb|������j�q�|D������W�&��7��C���U�xX �m���Z�R�q���ŋs���F �o��@g������͍�>\�D|̳�r�v I���/ҷ��h�V�D&��'�B��:>!��G�|��͓�<Y������$'����5p8_�<�Rˁ*Y�lr���©N����^�wd���(�^NoQ�F�$PR"�ϡ_fwk�D>���{������K2G�D�IT/��sh���4D��H9��+/�JH�����"?��Qz��K�fD�1�u��2�����ӸCLN?��{��l�-\� �UʧqvϞ���# �觷���{R�+��_*x{�D9���DnyL ��Y	�\�Л���ԁI,e"�<}�D�����3�����}�=;ru|az`2.)ieapp�=���V蔿=W7��#}��r��h��&�������m����x!���d�&i��&���L��+-��A�O�-�\d�P�-):_x�J��͗�yw,ŕ111���,��d��]/�_���l�#dfe��(���/\�7w�B�=��8(*�I�5�4v-�F�%���#�w�z�ҿ���C�SP�����Ϧ�U���hsb�az��@%��H��Q��Ѷ�"�Zn*r�-��3���n�L�?-v�
��˟��5ꩃrBF����T�����Ν���ݥ�&�w�z#���^�`��2I �n{����ϧ��3�j��Ͱċ�A��K�ɿ��"wZW���!�>�vӌ��p�힁���������뎔�9Ӗ��n��?
*"�.���Ǐ�f�<�����Sq��8X#|K۔)V|47IK�����"�������ù��I���ߊ���<��5b����}��]O�^��QefɊ�ܦ7��,��=b�.�X}�������ɅYi�٫^�r#��H���	�8�jS�!��+!��`m�ddP�mQ��v���{���%'#��ΌI�b�qJy�����׆�}�D?G��n�hf.qu+�W�3���O�<㪢���aޗI ��ɛAk��Uk�a�n��F�x�r��M����? ��,��Lꫣ �b�}rOL��5Ð�aX\oO�G߂N��"��>Y�/�P ��=޴��CZ���xkp1�D,8U=�FR_��������
k�ۯy���¶ˢ�m,^��R������b�>���cy>�얤�=�\Ǯ�r^u���!�I��<]㟐��A�^���;\B�1���rz_SS�ι�%mܾ�	t{[P���gL.�M9��{_dK9g?K��VZ�`w��T�'�,��Va3�' `���龳�Ȉ������y������2rAW��氉H�ݗ6�L�y�>�|�KDF\삤9�nZά��r�roc3� ⋳�aaa7�a�M���"���ߘ9��,��"�;�)����%-O�hmm-IK�@�~VD���$��R8��d�d���3���勝o���"������dB
 �2w�n�6�]�*��@i���_�~9�>}^B��$on�i� Ž�xqVr��+���s����a����!����W���1V/�R��P��)o��s�\IC:��΄\��9�<@���:)4㱕Q�]��i}}R��.wff��"�,8ωv\>4������,�E�i�R�_�,���f~�a@2@�!jsW�VM��C��b	Zr�ut�A���FJ���C�<��B��
�.����ǫi7�۾y9 o��� Tzc��H���Оu*�_������$f�ȩK� ���?@7��>98�Y�6"|�4���
��zn���2�}��YȰ� �f.d�Οkՠ��vy+�>�+�]l#o�F	�
axh��C�Vs�q<��S�F́�.���杌qF+:v�A�jb��4�A����-Dٴ�i$ͧ�P[�D���������g�ك�7�}���J�W��D���jލ���-vsy!9���B��mSoN�!��|�,�~l��ɋ�XEH���ȇ�牙��Q�ǋpmZr0'''����&�+U2��99����O*����m��� K�۝�o7�x;r �����6��ɽB�/8����C���-\J��S&h��(�4uww����(A�y���t�ģ	����)����u���(�"�5�����2�0�zrкw��ŒL�_(C��x�FB�PK�ܹ�Z�����5Q<���T!!!&ox���T��ȃ���s�{�Gq��l,
S���M(�m���%j�ح���Z�oC�Ȣ��'+[�q��L$T�|D� �§�f?��+�)�S�y��Oz���P��rA��g0k����#����g�t���;@�	r��p����ae�I�*��r���
F[*��\G��Oޑ�(2��~ �~?nY��X�AQՓ�����ŴJ�Ae3��\Csss?xhߐ�2Kz�Ei���H��翧������m� �7�X�n�Þ��YK ?*���#�/��.���$*1��Dn�a�	���!�Y�2Ɨ�hJ���(EZ��夰9ҹd0@���c8� �=�Ʉ_�������L ���<99� � �1�m���S3o [�ڈ��y
)w�i4�;A�����y���E���7hIjc4�����B�����u�>��4��a�7�0�Rے_ul2��
����Ͻr��O0�tv~C]��iL�9�p��d��=� |ҎCn�z����ʯ�Ku{	����3ݗ� ݟ/�XU�B�'���n��� U�p��*�]A{�@ݦ��Β�1ǏW��7,`vl1��m�a���S��������f�<�9]}}"H�KLӟ��%�AD<@��҂�e�S����/��w2�?�>q�l�hmm�U?xpV�`�lA�-�
�>��A�}[��ks��-�%�f^�"[����}|����,�d��db��5���Q�"���9�qh�h>'�����7�l��0�yW�M�8=�ʀ����%��q�prDW�%�c�"GV��n�az^�S>c$$$�c-�V4�??E�����ʊ
����J���c �����!}�⹕O�e��=��J�������P�����Ǚe=��_�~��®M�L��~�������`�}�g�!�2G��5�����{�w@�y9:RLѓ�g1�xaD̛@���M�KHH������4������;�|��ۡ|�vd�y�d\h������.�Ԫk��R<� ��A���([�+�f��0餴����w�n0}���K}��<)����)��ME�����{u~%�0�ߴߡ'�=!��e��U���N@o�A��ӷ�Y��
@z �5�M�� Pe|C7��I���D��YB�gqi��{����?K���_ ��C����?��a���0��`�sD�6���I<��F�d�"�ws�����G��>�X����0:���1�芆��6�j��;"��sc��pG�W]��:I��$����<߼LB�m6S` R 
�yϦu����N~]+��J�C4�bv�]�ߎ
��`4x_���%J�4��r��=�����z�Vj�J��"��ʕ��j7 ��=�!��R�}�'����U��y�pqӨ����4���w�0������+�� 1(en(ʙ[�� L�N����z�u1D���w2��n{��*��C�.��a� #����NrH�i,��>�`�2�P���|5�z����K��ECt%�"���9^а�Q̡�������� �"C�����`5�0�9��I��X=$H�yD뚑h�K�M����X���0@%luu����5��C�$��N��=�ʛYWEs��.<�� f3 r�h%�:"��0d�yu~���̪�_@sh��_*�B�������I�!�ܞ�ۃ�<�V����.�C�#ȗ/]Z���}���蝍�"œ3��I��!�쉾ïE�����m�0�P@1��g���<rd�=��c�p���{��+4��K�ݶ*m�'it� 7P�$z�!����L��x����Ƚ�_ׇD���Wٰ*� aZ�O�VeC��˪&0���Z!9��[J�i]]�\`V`V��iG�z�U�ly'S��>�G��I�(��L~Q�^BQ��K.�r�:���B�����M."k�XzK�'-}�b<5t�{��vUt��d~r[�V#mo�_uQV�AJ�bs� �n� ����9HEY�����m�>7��I��.�X��~r��b�������C�9q=g�Tx�n�[�������W瘚!�$Bڜ=���o�B�R�`!� t��s!��Ͻ �΀��2�'�h	�F�Ɓ�MK�âEi��>ri�i�i��3�J.�y��t,M---E2��8�/ �'����xe�Q�z~�.<�
3J��b��P�4l7��jʊ���_��g�o�v��\}kNT\
�JeT{�rM���/m*�TY�o��s� ��@C�P����bt�5��|LXE�
s�e��o90�&��!�H�.�/�\Ho!Ĝ���J��d�rP�467g�;%W���&�Z�X�b�2߼�{g�^�N8��激��[~�NLL6�;�~��Om�'��0�}�^X1˾�p{CQ�Un����m�D����/��?����}}=������6E�Z�@���*@����8�u����TQE!SȈ�O��Ulz*��͍Oo�ܽi]?>@]��]3RD_��pォ)�=V�����pߗ���)W��gmh�Ԩ]u�1wU{�.��T�J�"�P��N�"�Ko)#��(�.~l`��� � %(F$��j�(���h��ס���������9����d�O*�8�D��O��Q	�c�{�����lyPܨ�oU��[�^�Ԭ,27��,��<�w��.Y�dRhb��(u��"6ɻ�%�\��@���K3 �Z��R��SN��q�+�{$'�.k�
�\^�{y����	���:޷�	H�e�rL;��D��3z���N�����x�6�< ß>�6,n�p�ܞ���3288H�%���;Y���I1��r9d�Cz��}�:p~�\Ԓ�5,��
�Ld�	�0%�R��a���9����R_PN{��_0F��U�U�	�jܗ�&|��z�pܳ8��P/u��_��� <Odj�����'%$�5� ���kU�șq{�&���ͱ)��7\�}�p��I� �h���k���P���? �0�U�����}�re�Fa�[�����Ew��Ukp��y�:��0ԯ=3����	�*c;PY@��&d/b�P�/�*/Z@{�?m�Gϟi�;p^ ����0�7����_���-r�k>��Y�u�Kj�Փ��+@�~����C��WZZV�1٘)���G���谂�b<FCbՋ�fEI���C�:�� JM��	�'���w��ע	oG7�K8 &R��*-Q/������1��A�dNI��A`n�o�I����"�.�G��Q���b&�l�=NM?��������>7�:�Z�����l���.rB�[��Cb�P#���#�؎�w�$Ԑ]�J&y��B�ʔo[�u���2�_�+	�W�����~�CcH"��}
/[F�����3ZW̲hT���c��!	L������Χ�8����R�����t�ӎ;v��1�RD?� �r�Sl�����8��x�9�����tP�M�>B���� ����I̒��5���8�[F��`Β�S ;�ZUy�������r�D�ߩ����:)�NxE]�8�ɃB��ݟD����-�����<f��
�ʚ
�#��&�e�8��#�?=q����&���4H�'m4�)Ed�O�gNG	�>%��ٿ@D����Iּ����Q��d<����v�c���E�c���i���ifY?f�C���9XE6�o�R2�Ѩn�M;��s����Y��� )0���=#��9�ʓ�pcS�h-<HgY_o�FU/�A�4�u��i ��w�O�@�5Q<I�vy��0C�2�H���<�g�XL���ܚ<��p��$��m��t�d��u�6��3(&�]�̑	w����Y����b&_��Peؗ�=�Jo��)--�y�����H�Ul�vh�3;��:`��N�|�g�r*g��T��
Ӿ���L* �8'J�O�8[�B�E��
0�� ���N�P!m����
���W"?��D�0�H5)2���@��f�q��О|�nG�D��������$>ޗa��C�\�b�ъ)��0����~�_dmd���D{��cR��^=�D����#�&�����p�[��Ź�� ?�B�`П�����lϣ����]h3@p# ,�sss�����jS��*p
��v�H�ʂ�S�{J������$�Bg�	��1'g�I�3Ψ�%�78�˖�����f."���A8Zan~�z��z��z��Ja0��m�X��џ��^#���}�%�3�Dw���6	���+��m�=Q�q!�(#�S1�}����>>��d��7��l.}>�諸�њ�&�d6V_!�;�P(Scِ��mݐT�4S3�������t��d�B�܈�#�c~�f瀀 "����@���>3���/-*�z���w�_��۳�c:��mr ��)!�lV�����W���F_%$Y��D-��/���t�gE(������{�7�j���ї��������x����)&�U�����1L?|���Q�Q#�2}��ɞ�UvcO��	���{���Ԃ�{Ԣ�����(]���O9Z��=�ɻ ���W�?�ȉ������6�v�ax>i��Z)xQ���0�,없u��G���|J#�:ט�c:�|�ͦ"Uc���ۨ��}���ڙaSy;m�K"3��|@�0/S�.Ϯ��Y������<�V�뗻�f��	L�0�M������L'OG���I\�B!�VFB��a��@ʛ�f㯎�'�߿_�6��x�x�5�&/OX_ut�?�yXSW�6�>�ѶZ1N`E�`�8�d��`�BFdF� �<���jD�(ATh�Id�bEP�� �2
bd����ɉ�~���w��{�?��pv�^ý���>�lQ�i��$��~�a�H�H�r�j�N��$�9,$�D���ɾř����w׬F+o��G�����[3���4{��{�:v`s�Q$z�������f��#m3��I���Źs(J��KJvμ5��;:�����{�!�
�=�I����M�՚���x��Q����m��h��hkp���a���n �peP?�Z���sYYY�.m;?��T��q��b�����;7�����ώ���vF[�8�����:��$���U�
r�9dM����EF�������{�J��/�r�}s:&6��ь��qX�3r��uK_�h�������5=9Z>L8��Ȭ�cT�Dw2����h��������ӗ�]��ëK������;�����6�L}���mY���v������S�no���ǟ�M2L�An�&
���D��dXv�Pk��б��.-��uK�;���ۓ��[6�Q�qͿ��59��a�"xpNN~zT8	~�)�i��U��>CCL'!��G']'���>F�H������/b��}�	��e�͞�7n,M�i�!���j�	(���:��>X.Y<3��a�Q$��R衼������5:�h�ɥ�w�����9��]{�z"���CC��?�ŋ�#e���n��_� �I��X''��߲*ͷ��M�4�����������zFڡbt��-��ԸH���vf�?r��DRg�_O�k�g�#K��	�5Z��_�6�VuY��]n��w�{]��Gl�EEER)���xzg����5q<`�U�SN��4�dt�;����ӟ��6]+7�
��w�\[� �<�xxF��ٻu�ɓ'��#I��L	щ���!~ꭂ�\;/95T�����O~���37�X�"��4吴�����������"���m�K�������OY�����{/�Ժ�^g?*v��p�xy{��Mpy��7gd#����]�hv.,k(�gӹ��Ш�wlP�������'b�R�A���z,�-mw�1�A�{tt��q��=vd��JIh����X^����Hc��c&�T>�5��tS�鳛�|�'�Z� �����\�G�%4لϤ�!���@�{�����8��;�Ҭ�bC�R�$�����-���m�Z(Zy�<^�% 83~�AG���˹�Qf���_|?��l5^a�� }�oJ,��M�$r �7Z}�;9m9��7]�mX6R���9�b&s�a�o�%PQh5y�[�g�H�UG�&�%�C�k|@Q�P��}�j�������};/o��\���^��rG�g��z���(�9"#�V���Z�Mo�y��<���J�m��I��+��2h�h.��f'<�O�>o/�\J�m�D�I�?W�?Z�R��ۺ��U�!�A�./�K{%B�9��æ��(��BÊ� ��_��c&��v>�-��S�jQ�~z��uѕg�`��7`�������Ѳ%�D�� ]�t5�<��L �Ti�2̵ٍ32[��<�#������$�oqm�'�ϫ�Ҫ�P��bmH͕k8�R�S������]�頻��hY�h���ݔ�h�4��"E��q���Z���4/M��`ck� �ޅ���+w��-���L�9���Pv����?��"��뫆jk�e�k�~�GHww��//6D�%Llv*��ah���T	R��� �2%�������!���Y��[e.��^��|
nG9ѿ�H�_�B��N�-B����JhKS���gF�"�ۗH���ۺ5��z�����(�N=����l�x���䌄,hBY��c�":����j���ڮR�d��u�Qc�?�Єb����c?i]���ѹ�����s�g\���Pդ���9 8WS�9��'T���EE)x�?M��z(w�8�edݒ�HT_��4�A��b�n�����,�Ԗ�R���2 ?�+6$X�!`�C���@Q�:���!���w�(��� ���bQE��S�Uo�����.��u�w�A�/��;�F��62ԼLLb�UI�=j>��>Jrrȝ*�F(��j떟�b�y�4Լ��uQ��1o��5J2x��=��Z���J�-Gx1����L7k��k�������D!R]*�9���T�}��C�^�z�<��5ڻC!mbr��PT+��&���\�j��W��n�dZ�v���ˢ��~�(�E�n/)��yad�*���O.i��GC�TԆ��4�Ri�66wՅZ�,���u��=��ak�6Q���@�//��x�Sߜ���*v+��l���ބ�U�W�r�y2>�����/؂ |�?R��a�O6T*�^{VZ�c@s}����j�,�e�)�SPL��������y�L���E
豐�L ޑ\��[e���l�s(uV��=�Ǯ�,]�D�_��PTO�O�����Fw�B��(�
J���Bd�&����P�B9[[ۛ���A�N' 8X�İJՕU�[G����1�r��6��� ��JPX�j�VDC���@�B�9DX�I&''"w�6K�;wN�Mk���2RT�K�p ���䴹��^ͯE��/_�loȰ41v}��A.�&��$-A��:�읃��ӊw��6M���qAY_6P�O���$l��[#���ޕ���,���}|r����uW�=�yEɶ'ߥNl�8�w��Z�w�3��4=o�_����d�o2ɾ5"�e�a��j�g'�&�wn�l~2�>d΍م#=��#,���l$�ܚ�V�Ҡ�U�� c=�N[�p�Q;;���_`�H�:�MQ|��FG;��+�����L���쌹zu1BO�Ug���m�L�:�3H��Ϡ`��_~izzzl���0�:N]R6x��W^Z�U�����2��<�����Qs�w�����Q�|P�q�{�lJJ��P�l����ڊే��;+���w�����؄�| �=��,|�4A�mv8��~��{4��~�j�R���nn?�>s&a]���7��^��D2D����_0���"����7�L��H��B�s�Zą��9P��'���:���J ej=�q���ڳ+U�8'�������㯡ms��,h>�=6#/oEee����t�t��� ��;Y�����	�)����ޘ����ϟ߮;xJ��H���ciAAAFF5ǩ9���J��g����ʃ�"s�Mq�*pt�CCCȈ�N��W�7b2��+�0����X�9E(G��Oc���X&Ky ���� 7��ۗ�0���A��P�����/P� ���5���D�yc���p櫰j��y�P�)@�]�����A)���T
%�.��447�CU^�b��_�j�-��a=��Z&��
����a�4��sؖ�=0�
i�~Nc�m�
33��:c�GP��s_�j�	1$���������ROf���L�vV\V��3��,ok���b,|�~�h0ǅ����ٖ��j�=�H#*:���w��TKZ��>CU*6"�m��2 #��WSm���jpj�k��� ��&�m����^�EO��˄�1�o�y�ˏeeeG]\�Bo��3L�x�@�����PM���:8;���U�˹�G�BQgQV�lls�ȏ"w͝�񿔶:���}}e	�����B�Ag'v��.4e�%A��V%An�/�� �'&%������B
_q=w���>t�6'On;+�=��wGf����?�t��`����|��/�����f��c���3Щ���w�?�JQ�����oٲ�����Q���~MY-g�p�
�S4;�P2`�S���������>/���%%��Q|���n�"�svV��
��
ԅ�#7 �S�Y5zcc���_<��h��!���d.;s挫��"��B�+#����XQc~��֊p��������h�u�sԽ7��}l�ԍp�546�C��
Z�E�LmEQ\��.������R&��i�� ��+W�B�K��C轍��4
��eF�g\=O�w�ȅ��)��^�q(M��CyCP67���!,��{�"˜�U�6�=�G��]�_�����@X�:4��!6`��Wv���54���'��d�fdli���>�|�9�1#'G266�j�����q�q�"����z�C�r�޾+o蜤bY{�Q��k���i����=������#(���Z&!���|��ڈ�2�J ��xj�ʕ+�����]S�TJ������.\� %-��x%i�v 0����G5gfFK���Eb�ő<0�����I
$�/G�� ^[vɒ%[���P�<S�����ii���$CD	(��e�z
>������i�p����88l<}��Qk�c)SrPWI�Z���2�2����i����K�Z�9��ޖ�u�9%ӎh�*�]x4 @ыe��IT���ǐѡÕ��уy��wzM%���99��2x�5x����"��e�%��*��+��F�x+pY�`�%A���������ֶ��ు#���{F&�	�&��I�?}�P,_�rM]vժpD�P��Q P2.�}�d�UH<�DoDDԍz	�Y�cЮ�x{�v�0��-	��NP���B1���%3��I���nY4/D��[�PB�c`@	K���C��P��"N�-~H1.�+Fz&+͋Ԗ/_�ޔ玲���<�s��i���)���wRS'��ii�tx_�b�����s,c��*�j��x���[�n]���Q����ɧ#���{	�Z��`�rd"�Rh�j���u����|����!Zr����_=��s�2��			��R�ԉ����@4LfѢ�`�%�^*�X�W�J�[����yn?����om���)'��bhz�
Z�1��O�b+O�I��j�h��I�i�B*A�EC#`1��D������zFn�v�4k��g��x8�<���x����zFo�Q���uy������ݻ�'N���׷9~|`�S����Le�0�PD N��X*�A��-��1�Wo �@��E/w��M"���K���

������	���~E�|�_}AQ���!�kc1n�(vxG���d�[W�jkˢ�J�٭����<Ӕ�&�uz�nގ>f�����`���_�A@N���e��**o��P��\K�$mG@f��Z�������1m�O����ً��j�]�^�&��q[��K�-�Qύ�=��Fb���&��ޫ@���+{�����F��1әj���rI!��ޔ�1�������-}�wo�B�=iZ��Wz>?i��]u���T{p��cG(��,SD��z�� zN�`���%p�P�B����a�Yש1�x��o�*c���dZh;C����MN�l�ܹ��nZ.�Mٸw��3c� �y��}���f��+��q`2G�ׅ�$�����>����p����
�������!V�_�xQ�_Z2#��>���1��eY-}4O���YV��u��8�*�n��3��b�^6;�,��XҸ�}u�����L���$����3�OK�q������Z�	SN�Kj��͌:X!�]?���r�-�B��,�<w3fS��{+o�;&�z���P�K��d�;kr��S-�̭�{h�\�K�vKz�Wʡɒ�kb-�nh-�ܹs��ڛT���x�%�D ����k�\��bQ�Eu��ES���:f�৫�����n����#�[��M`��m3���Q��VP#��ɼ����f����8�\ӑH�����@���n��!`b���������4���ETg�R�x�<�{��F�v�?�2�h�U�۸{]���t�����/�t<��,�^3�Y�7�0^���x�k�FV)u'���}ҳE��mv� ���{@Z�t���:��4%�X����Co�@/��B�{,z3f�{���L�NF���>�&��m��]�Zp�������AE�c�����$�x�4�����<�kXE��·C̺}�^�RhnԩK�'uܕ�����l���3��?��(Ċ	�f��u5�	��)��]�:�b������
�&hU���,٘��<�Ӆ~'���b��xF�&���"�fb"�ewo�i���on��'k-[��?.Z.��1�>�:�����q`i�!;v�N}�!����k �86����~{����̺��r*����Afݎ�u���EW�\)Ki!�l|���!J�˜�q���~�;$Kzf2Ug˧��\7׈>�:��^S*����M��j�w��JX��� Y���ؘ��ð?����+�$(���v(��g�+B��z�����_.~���○_.~���○�]�l��<�p_.~�����&ǂ?�ƿ
�W��X!�|xQ�W�/��|���˧/��|���˧/��|���˧/��|���˧/��|���SHCސB�`����ݹz��&��w>^��|�-��Wت��N�Ν�=j�V��),�n)��9�t����[�Q�ϩ]_��8,����_5^��=f�M·֡?�^�ݓ�7�v^��r{���oߢ�?Gӄ�����(�{��z�T���/���R�������������I��'� � U�`ݶ�������~�杰�q3���Ʒ�j��g.�Ő���l[��қ�|��!��C]]y�=<F��7�B����B��/�吪*-��"�������$� %i��6������|��-�I��4G��-=�Iڈ�
wʙ{����.O�r:h��9>M� R,�v7Au!���?�e�#𦯵�翺yY�u����?ۺ˫@Qd�σ3tBΘ�>�����_��i{9�&�9�r�5�\^�Q;Z�h��[��:�">��*��C�^R&!+�f@}�E�9B��ϒ����I4�������?��������:�
݁�E����'Hy]Z�uNQ"HqK�O��W����"%�u�h.k>y�Mj�x���;����3;�7���M��`��{��k�T��!��- ��uujτ/!�C�XdZ�<~�vH�=kw	|��E[|��/��Z<�R����b�H�tCbӝ}��1SwA^?���g�l�ӄ�gE���t�]K���N��ލ�ݻW{�*4�_�������~�������^x5��a��b���K�#��FdL3j����N|�w�p��0���z沃������m��y�{M��~b��9�*El]�g v�	|�׊����\O~�.1��S�ߩ	��|��*M�b�M�ޞ]�0#���g1���?44$q۶���z�q�֭[�%`Q��V��
���G���bQ�
�ñg����1RNJJJZ-ŏp�K����!c�I�8%�ڮ��������Еb�|!��^'ш���>48�c����9$���v�Fm����J��w@S|��������鯲����	FEPq1�3(��7e�`M_�6���}�����}�}���>�z�����LjP��hA����2��{Q`��SRS���K7p���job%^Y*��Ou��Q;����o��W/�W�z���c���G�R��Əa�6]A
]��@���+��Ж'� �d6_b�B��8��%��8v옾���(D���]�Y�`36�M��MॶLd��+��wy=+@֖��������sZ%�.��Q���Y�����?�< kS&�!A1sI��7?����mXPI�~&�N�6���_"�'���W��%d�$b�Ow�2�ד�َV�q�*=��p48*������~s� B�["8Z[LL�X�P�����T�kE�I�XZ��K�]��v,P�i�Xd���jv�M_�M._.)��X�^�2#�4h�#.9��z�*�e�_��0��/��E��i}�T���^#�:�ho�X��o��Q|�l�+,�z�C2�WQ����h�~T�q���®��~�:���]��,�M�{/���e;��,�w>|�LصClW��`�0�"96��S_UD�� N�ӂ������Z!�j8 #d��-��8���?�ˏ?ϼ2w�+Ne�֡��TH��h�`�Ka�cc�5�� ^�6y���嫒�nv�B���<wx��Ŭ��\�������-v�;�z���d�.YH6璂a�&�E$�+��w����rW�q�L��ܷ����h�u��2,,��F�Ɠ�s"���k���֑f�M�Y�#1�~�Yݿ�aI�y��n��z����Qm���7�8��p�ޝ
���!z�$�˖&t8!ҡ�v�BJȷَ�g	�m�F{X�
�������m$���ߞw��7~JJ�$�����V2�uw8C��lֻ8&��b���"��CNt���.fu��YU[{�<��������s{웝F��x�ʑAud:�]�(�:�����s9�S�A��%�1x+��ա�x���'�O��u���Ѻ�+:��.\�c�Ĉ�����K�E�:���"���M�w8	�K����L����#�1BH^FC�`��fvcoK.��3B�ޣ"�$���C��������I�C��t���zp�������zSzvI������!GHQ��*����ڔͰlV��%r��*Q����j̠�#�L�r�e*�1O�1OԢ�5�a�U{d���D�\pNd��C��H�+N��9�Yw����"u��	CJ�ur�ѫ�n��B���.{�'����l�(�V���G�p8J��L����c��dait�v]��?ڧ��� >Ml?y��l����v���-�و>�	�NK���Q3f�>b�C�r�`)м6��1=���	��;����K	o���n#}��ź�:m:m��v8;4z�kK�����%}��>��e':6/�������`�DO�B����-L�R8H��k�86D6�jұQK���<)�� ��n�e��M��^�J�������O~�z�c�Q%h܀��W�S�=C�*ۻ��߈>�	�:�&Կ�Ʀ����w�L����V(�L���̞w'bR�%����]0�ӧO7E[x�J�i�.��}ߜ��[��!�߂c���D�s�%���7u��i����(i�ouy��x�X.(����ˣ5�/;�J&���ry���l�qn"��`���5�'�㝰#��Jƻu~s���{_��z�Y�e�LD9Si����Lv�
���W�%��aH֐$�_\}NCz���߰&������հF���N�@��YE��ty$�ꋲK��
�_Z�����nXD�8���M�t S�}��F/5���i<t���*��Y�?L&�6:F)�|�� ؼ��(�� .�t�K 9剚���Oq&��#��"i0�cD�B	,�%*�~s(^6�����6A�)��m��s�<��	Y�����:���)����q�����v �x:m$��$����6�1��<�A'�_�|��ZK~��i�v��R�\UB4�kI������ۍ	��{Ж��9���gn�sA]��-Mٽ�7	����No^�-0�qƏI�KZ�F��
�ۇ�ޢ��Ĳ۳/O��;�&͝i}��S��3駺k��/�*(�<4���P�Zɹy3L��+���0�޺mυ��9����|��,Nյ��3���i�0����4�Y����w�%M�u�1*R�0�0��Ǣ�޽{���!�$Ϝ��@-��nt��I��؊�FJB<¿�h4�ƭC�5N�k.H������	�������b%��ܸrc&�&�q24��� �
s!9fC�s��*��j;4��i��@�����ʊ\���9*�Y
qt��F��%	CJ���N-]���,YB�S��r&��5���ڗ/_jeܿ?����}2���i��I0��������$���4B�yA[��w��p���':ke�\�޼~�>��.��MB��� ű��w3��R+"j�/�{31���{@ӓ��
\3y%��	}�w��j��h'W��+��PN>z�H�`�-"~���?q�]�����w�z��j�"�d��znTpc�8Z��;��L��+�$;cL��ǯAk���H,I6lG�i�C"&�PW�����]	ۯAF��_wx'�q� ���d��j�B�)�eA�h�tZ�d38��Qq#۱�n���4�i���N2�]�Z�}��'�y<A��C8�0=�.�嫞�Ç���Kn�p��F�Q�6?A������Jr����v�~���@��l%n�TE��Ũ�G$�=(�v�CMM�/� |k�E�}|wӻz�L�gR�S�EV${��1�Nл��r~��K�����_ze��ݗi�,dƍ��l�k�	�ȝ����)��i�?@h��4Ӹ��'y�v��MM��ٙ��S�d	h����c���i]���j�ˉ�������A^NɢԘmD���(���D��EZ����>�����X��8�*�ᑀ��ޕ�[i��\v,���`~�~���.����/Bͅ�cmE�QK��Zl��`r�[��5��g?61*��Ba�Yl� 2��<6�ei_g����V˸~d��H���}drz�;�e���G;��&!�<R�{P�y��<��.ȼ��p���N��{Z�d��R�D�(��z�ѻ�f;��poL��G�+���Aiw��Uvo D�R��2&��!L�S[ѓ��p���J*��ǜyZ����urZ]�n!Z̏�d~!�}3�ۊ6���P�-nVb�H��^�`P���FR������ׯW���!�$"��Y+Jۮ��z�����Bi?�=�3}hk٨c��UG;�1�7�2����C��i,�K�» !��!Ӹ�l��&�V�&���T�"����nU�֊rɾ8'�/���9�p�I�yML�삤�tٍ����X\��]y���C� .//��[8���3�Z �4F�DY�29�˨@��R���~�/�v��B$r�Fj％�c{�]{�5���!��0�ג��Mh�&�D���3SLk� ���F�7�3��P�W������8y;O�������n''m62��Ԟh��=�)�Iu�cED���꯳�
��c	��IS������,�U����f|�v�l�;�XG'r>���F�VT-��Y�Cm�J+`����x�G���Zx��x�Q�AsFz�@���H�}��˞,�Xkd6��D���y�E���*�ԑ�'j���J����&��hn�BJX�.�	0RO��M*���uE�i��P�g�:le=r�u�#�ni'g(�1;ژ�Y�~f	bE×�V455=a����N:�Xi���Y�=��pʐPft0333s,���v")�v��iUU�>�r��.[=~amz��tAἁ��Fe��3
Q�F����Y}�t��3�qsP|���k߲֝����c9��}�iWd�qW܋��>ZDV�g�쪯e�k~B;�+�c���d^V	����G;�ʙY��		_��W���Y`d��M��T��T�����*KX�Q��w�3=m�;���.�޼iS�$��Q��mȝg����p�B���r�8��t�A�I�.[(�1��.�GFp�1�3F�o�o��y�����WL[_<V��ڳ�CJu'ù�8-��"�I���p**&�PP�[@Z݈�d�� ��o�?N�z����{�ky�w\����'jV���L.�xد�=�32S�/d���!�#�]�챀�~�ظߡ��"��!#$���%��g�<������hoIl���������+�&�;tZ`aj�&�*}9��N�N��	Z����	Ov�1�I��7^�k�
�Wډ�h�z�wb���n'�˝��^�tZ\�-�^_%����+��r�$����%�����(����v��/�Z��!X����	�r�Q'�*����ۈ,K��_b���d�]����F����lR?R����1e��7]Y��:4�ot��co%|s����<
C��$��܂ſm��������|������B�8����,徖:�煝����������ӃA�p������D�S|�;�D|eψdapSk��I�ȝ:���:M���c��]qP�����	A(�⸲i�@(��s��L�;���ߦ#2D�zڻD'��M��ˮ�y`��{c�Wճ��z�
���(2%S��Jl{g�kE��O��E�+:<��aKC��U��0�l0y�`��y��p�Dfuͽ���s$O�Z��)}�Ԟ:择�\���i�KǇo��0�hTDB}ϴ��9V�������IE��AD�!K�g�j�@�£�r��$�!����cI�|�#NP.�����~��,^)W���̠%r[�[ᔾyx&x�\�Fx-Ӌ�g"�B�ĊZg��v��/<5O��RT����
g��)؋���N��V��0m3L�?����9��:�k����J��~�t��r3w!@w~%�e��x�]1*H<��bv��9��~�o�����q�1N�] �2ΐ�^p�ҟ%����Uuj(�B�DCI:���wF�=��}ѽ�V�*�;_+������?~��-�D~_��_r��޶�♈ C����ُ�5k/��&#�����C��a3vװ(���އ�^�Ȳ���D����)$�y�N=�c��"��cG\k8k�X�\�&�B��K��Ђg�-��c���r��~�K��J<S�g���:Q��Rsz9C�W��SO�#�N-&`y����OD��X��U����e��C��.�)ii��u��Q�^`��<����a��dB���뙰r(�e�C��h.++C�ύ$��4K�u�L�]��vE�!�4gtr:M��]<�mC���bj�%R�s�����8Y�Z����!6����O��q.6޳<�gb:��l�V�2�Lf?�U�<+�����V�q��w碚Nʐ�6j�Xc�x�� -����;LLG�D�{U89�&g�����c�N4�VTT<$"�Rd땐˼uK{��i�s�����a,�yJ��N(��Qv��2-Ea���j�i"�2r{��T�r�RĢRf��z*�:�1�y�!2d֡)@����U�ȼ;M����\�/�
��R�F��0w�[��U<ގ��33�������*�.��bټ�5?��x}��d�!~��=����ZȐUnР�J@����CD�+6G���n�͗N9V��ޗ�1�$�Y�`�U�8�x����gW�Yb����B��QI��.��F ^7i,3�}�t�!��<-с�}[��J��S��#VM��K��2��a�ݑ#o�ހ
�'�����8��]s�ξ�76�gg���N�|��S��K�O ��o�=W�\魼H�U@���y��~y`���F]�L:l%�2V{�$K}��u���P��N�A���+-�����������i������֒�&v��tP	�@�p�M������ڣ��\v���w�<-�/G�$mO�|(u���>�ܟ��3�6�S����w7"���d��i(���/݋������kll,��ZԊ��U�S��p���T�4EU�?j�� J��ѦNv����֦��Y����WeO�i�k;����k�����(�jPI'>�v� i�gh/��w#z	��=x�,]àaH�V�]���_�������T!δ.GI��"���Lt�!�ۡ��y�9��PBKT�I�xZ�6�Ȋ�k�@���`�`���N��%�cl�����C�VrE�����Q�&9��ۼ�	v�Il���{%��q�nk%G�u�ʪu	����#Tc�\K]�h4&��_I~��/�W�ASAN��v('�����oe��~�
1뢭��e��A�H0�=�z���l.\^�� �t�%����@��� ���[2O֧��y�f���t=9�Ξ��h�RgD�1�i\�p��XȌB6�S�.)��x�tK������GԄ�sO=�/6�-��}�+K�"�ڇ��?p��k���̍ı�����?�̑2��~찑�\OUi����d|����c�S��U5�u�]0Wq��|r�,�7�~b�Lò�E�❮��港G4�TE�n���,���/4��~�Z��sӴ=�?S��V|�i�Y �?8C-($k7r��FFFVJH�\!��� �P"�Ÿ^���ר1�I��j��A'��Y�Q ����Ij��?C3���)m�F|�&q���sO%E�間���W�2���b�s��%5�UCS���1�*����}5�&����D�+�Fw(?�^"=���gտ��4F��5���ҽ�N�9��I��m�|II��2%�O�ٍ�;�޽-�Qi��Oΐ���OU��u�p����=����o�!ghH^kL�r��R�%IXp��<�����!�O�+�X�i��Z70`n��Y�66�&Z�	.B�Y�3����*h��0F������ϱ�7�|�[��6�n�4v�y��b�t����Dʡuy�2l�l�K�a�܇����`��>�G�z��k��3 *��-����wN�($�|L�y0�v|�]S����K��X|dH�a~s�j��kbX�Ӫ����C1abĸ�"�o9��_���V`W�:J,I�>�M�$���ơ,m���Lï4N$���z?L��\�X�gv������� �I�SG��H�|���(�쀪ТV9���X'�Ơ�����5挲��Au�Zr�ZR���yv�Y���[�T\v%�	��&�>�e"��ZQ����XY�(������fS��*n�.�"�Eh^*����(=MWptphҒ^���Z�y�7��^���X��CY�X��0��F�C�dp�j�@
��1�=�%�ɒ����gN9���W�c�cIL洛��	rJ���f���U��4��8|�gA�q";uR��M�}���M���{OU.��%�C����uu�q��=%��t�w	��*ӮZxf�|�V;w)5Mj�\m��s�q�d�~i��7�3��[ڊ�~u�����&�v U�E k��9b�@�}��h�����=*g�'e�=�6�4��@�����2�944�oab��Ig���I��i��z�2�b���L�SNkν{�c0����.e@s�5��$(rr�zL��h_LD���z�%�f(M�Eӝw/�c5	���ށ��ÁTW;P�;j,?��VM"o=ȭ��ق:�s�qTbELH���7y�32S��l�3eC��#J���TG�o��CC\����f��#X���m� ��%%��S{Ʊ��Ȧ�Ä�Ɇ$�����W������t�~�z��xW��%J���(�r�8��*h������ͽ�Dy�nN�t?u�q�T�&�Nk�"�P�����!�1377W��a��������}v]]]9f��H�0��G��VV��:M`����u����#4�8���)��3ќ!o�RY��m2��iP#�ac����N�u;��Y%��krVR�����9Tr��;�n�\#�vYd	�X�&�����d��-�H��p(�!�6	|�k��M�4��-���``���D�(۽�"A(�wi����ɳ��<�J=�����	���Y'S�lo��*������;��-]���Yo���Z2��M�+��Kk{FR�ъx�V�H�JN�ݻ��⭜����)�gD�|�@����"����Q�?�+��뷹\n��~����*�`d�`<����&�kG�\P��
�`#"<��yB���sqm�OE4����2�����2TY�r�Ni�B�w��o�J�?�5OFI<��s�˷�O��.���O�eT��"X�ho"��D�:��"�"f�e���L?�\�����䴨��'!qįh�|�?D[������yvc7Q��O)e��)�%�Kշ���g^�q�)A��%�$(3M���-����y�U/�yZZJJs	��XBcf���T$1Je�{d��ܘ���~6j�#(��]����������qq�°jBdI�6!�k�����qI��X�|�$�j����x���555�׎����R���=ȰV�Iy���N�_t���f�s�\���ڟ��l�7<��貖��Vԏ�	ԣw���c�6�F!W$�m����p��]�&�Wj�C���J�tel��DKօd@-q�����C���"����C���$l�b��r��[���L#X%��r9��U`�}�D����`t���(&��[ԥX2�z�CdA���	��W���)��{3�v[ٝoτ�ƃ���3D�ǜ��[����8"d��Qo_�ײ�ں���~�e_���p��8�p|����z=��[��o��}$f�pU�����Qm\��E�6`�ȠK��:�b�u�P�\��K�1G�\GnFĜ���_M(<}A*ݱ
����U��?������&օ.�By�Du����F���:o���֯�����cx�8�O� �[��P�l��C�z'�^�=QJF�D�넢 ��/���0�1�r*�S��S�����>�и������DF�-V�:F}eY�Xx�{�A���-�6:���j�j�p=��Cw�����(�5�<g�&��~�w��V��#ԟ,��n���$�K�Qȥ���{��z '%�+��zZh�d���m��h��n�Ih`��\mHp�#� ��5�O���K��ވ���,��{����r��E��	���
�!A]�H���FZ�<�o�Y�ΘQ[����y�|.��R_���t4!�Y��y��b}���ȑ7#�V��k.��[�"��r��#��%��)�kG���#bioo���^�.�:OM�7�J��DQ@�!�-j�s��%An�(1RjB��7�����$�mK�����eH�͡��lv��O��j�vF)_6˧���>TF��o�y�5�~����ˠN�;;v,���9"����[N������J�t��Ut�v��`|����N�.	�yė�B	i�'�R����̴��t���D�zW>�~�x�P(lՔZ���%!�]RF S��g�щ�ΐ�<	������H�����'��G1;]�!T���')(v��יh�*�tQ���&_��X�O{����過Y�֕2�?�;��r�djC7P5�5�(ʵ��q��?85O� �-Y��M���)�^���xH13�Ǖ�=��������؆�4nS��b8+g�o9�9�)fh#���%�[���_<��gЍ	)@�9g���)Ą� �õ��YE�갅_��Ox^ I(:
�"H�����=�ë�r퇴[��oJÏLf
�{^�^�r������<�!��Ƙ����j�JR��\1�%�~��gup7�A,b�I��K����s/V��#~�~�&p��E�#��;�i�Ԅ���#��~� �.�>��x�׽�@�y B�ie�I�����T��V��<��z9���A8�w�(6�{�ՄSOY��w%��v�=��ۼ�U�g�n��@[�?Zrܾ�"���`֩C-^+w�g�(��8�_?Frn��	�<v�tK��X:a$X=�k+&�"�����LN���Q0~Vk�/�21����5���w�ʵ+�	�7Cb�Df�Lie���'�!�Rpْ��cפ /L�5�Ί�6}��Q�u�%r���NN��萷�8¿>li9�������"�z�憦��z2��g�(kK�]�*��Y��>���H_��'�uے��#��{��S�jB��*,������c.��j��A���P�7�U��c34�_��j�Dp�u�C����@�\Ǵ���~�"THّ]�K�	G�{�����!*����)��ܽjj,�`oo�	 Zǽ��(ĨR-��»y���"�9��������i��n"�%8e�%��"%%%�qJ�o�_������P̢�~b)�9���"ەl��ty<�_i��va�[hÚ�r����~�U��������z6��y욡�˗�n�1��$� �ju� ���֒�\�.���<Ra#n�#Y#D(�I�_�N�Ԑ�N<��X�M��Rt* �ҕjVۡ�<�N���(�qC�k?K��rqee�5fG�Tr*۝��W���h ��tP�zt��x��)���32L/AA��a�[}��ک�P��@n�Q���X�8�s(y��:� ��B��goQ�đ̪d�N+�	��X����l���x�]�܏��5���@F���')>�=�����y���5�"@0�r�A� X@��i:�]�3������(��0��$�!�A�����J�3���[��~�)(&�&�6
'I�r9��<�evM��Q�����e�/_>���K����.�m��ur�U�K�S�����9�__�?\�5!�,�]�r�X�g6P���Vm�߈S�xo-��t�Vvיڍ��^�����D��jFzZ5���j8�uM
���䜈��@�1
ـQ��2��]:S�I�ѱ��ԓf��j��o"*d�\ ~r��q����j�:�s[1iH�x
>�+Q�/��ȿ��G�{(IM� �*�B6\ܻ9������V�vLN�7�������-��M�=~6�}ͳۄ�E��@����.k�*oB	�Y�,,��>�/�	�쯾3A�h� A���Dm�E'�b/g�Sܙ&=$��z�Y�,�>.j�Fn=��Ҥ\e��"�W�kį$�1��:�����)X��"tN� F��f���ꖢ ��:O��>���Z���X�r����/��^s��]��P��\�#��=�{8�i��{�$�~<�λ��7~��<d��۫O�&����e�O�G�{Q��=�u��v���U�{-��7���3��U(�9N9�v����1�"ף��	*�w��|�w�������0k�..�Y끅�!��n%��n, J"%5UKNN�ƽ4��(3'߽�ʸ����u?�u���~H�/X>���	v��N�ՒPns�'�x�;�@�AM�)�ދ 1&S��(-���,�Ă��A��k?���,��i��hg�RL�SV&�_���r��h��"v����F�y���(��i���:���rDkk`�wtoH�8����Ī���&����l�n&��~h���XD����PUy�	������ce�g��:���I��K�@�(����%�a,E̺�G-������ߠ���g��Lf���F9-Slv����yE����A��3����'�̲9Q�����Ch�_e&qZ��V�z�5��/1�����%Z�����ה�.ҍ;��>��Ri��Ҍ?ˮ1���a����>��z�@�I��T�S�+��zk�v�<yc%��3�������Q}_�mv�Rd�w�[t����5Ǩ��(��J ia�Ĭ�2�J-^�:~Q& N��i����8ik�_�֙u'�.�����5a��w��V�1�aw!{�5Hk�]1s���	�S执��?~����g4�`�L�offf�	�C�q�\�bC	�]K]n&�R\����گ�6�&IJiyw~�oyĪHCZ�M�q���:`��w�O��R<w�U�ps����V�9�������b��ݓ�ĠW�������í7.c/!$g��g�C�4���g��w�m�Lz�5W;w�;9̺D>N*$��׫u����j�X:mz,j��ɗ�a�g���Z�_v��IN�v֦\� ��_�����;��v@ʿϮ��O�d$�NNo�ѯ�B�:�s��ū�.�r�ϻGK�&�f��=(6vin{�C���f��ࣜ��M���{�7��g����������i[_�Z6(����!�5�"�E�@D�@�~�}ĉ#��3XQ@�(q4,Q�FQ��o̍>�R�7��{��{���~,���2�Ӕ����w5�j�
}��D��=�!��H��eR�R==�H�Q�/ef�?���nD����|��_Q���<��!���O����u�Ɖ"��~��:v��Α(v�U���&=��j��,\qL��)�4-qJ���`q�:z�␈��� E�
�Q	a[�l;����*\���A2�ˎ�X��N(���u6m���8��bVֈ;xZw���׏����^���θd���p7,s+�5��'%��8�U%b�8�fr33��!+�Q���[&���1���!D��K����#Ʌ�\�o��a+@[�˵�e�da�.Y	���X�ҟ�`ہ'oWh�-T���*ZNNNk��J��9����,\�Dת�(�>U�Y/r��p��4MF�=�?�|-vlԏ�U��J��!'w�J�w�Ĕc+�%��/)»8ΐ{�J  ^ 
�>F��_l;���O��:@�BZU��w��ۋ�Jm*���Օ6Μ<�t-��LƭǞɻ6�YB����X�
�c5�	>�K)�Tff��8��:��4��z���٣��@�o�lNff�K���k�\|�~���Ɓ�V4{R�MI�߸q��''����0���au�K���@�%*f��C���$��������t1�({����3����>����?�Fg#d	9��F_M2������5{y�o� o^� �ݭ{Fă�'df����V��H��Zs�\���ɠs�XK᛿x�~�w�]�C"�N]�G��-��eӣc�7�r�Y�jH�,�^�?�N�͜����!�`M��~��u����~�����Č�Bg5�3_���݇����W �����๳|w<�qi?���Gw��n&���?K�ea��ZW�L��f�k �O���+�Kܔ���sY��wtc��#�1O R�@�[G0�o��A?(��V�g���.I]t�#���[��E���L��v�&��1pk�k�z��	4��Ix�����O��V//�ALL9�
W��q�;_��U^�+M�������l������[���7�KJ�&��+|ޏ�� ���>��AV��ݹ���CD��_��v����"{ֽ�i��j�b�.z��E,��,?��
J�/���.�u�yw�\�?X��!nT�2���{�8ՃD�������D-ӐW����n��AF*�i)��lȝ�ַ�9����<<�$V:�v�JP�x�-��y���?Rec����u�_�RH�dK.Z����7�!I�H�v�����[����l[�N���]�����>���t���\�="׳�J�mҷ�޽یΠq��v�ƃ�6��c�ݤI{���Y���+�H_�u��g7��3)-���mA�J[Jcq��$Դ�k�g�����}Tԍ��Is�Q�E�^��F�e�>?בF==g9��Az2��p;�m	K�Ŗ��糥�7 �lG!���?�2��3<��`���t~����D9������l���|+��X��+�O��)`M<d��<^,�i][��	�RZ �FOP�̟|||�YWH���n�D�5JT��[!Wc��s�&v�%���gpLS__�J�]
������NG�$� �A�S�b�����u����nz�+j����Z��!�~Q(�|-�`�f�6�7�����~xH-�[Q䠦��چ]q��85[$*�I*@<d7��9#����(1����v�$0��DY��[�f6�p�b!��1��� G�M?/{�RÌ�I�Q�)���H��2���N:R���|��e�&q��n���?y�~}Bqa�Ǐn����z^~8G7B���.h��R�uFo;���f0�;"%�}H��:���E�*�����,f$F��U��7��
�u��@����%�N��O�+:21o2M;��7E�����n��n�g�u��r����v����y8��k���4������C��ʬ�&:�[�"��� y:��>� {�b"��n�]nۑ?3.$O�L�~Ȕ�O��xU^Y�c�G9��ƭ$��6���[�-�7���p��9x �U���
�������]���� "�&w�o�<$�`ڜ�����y�Ђh������
��Syi�K
&R'���Č��G+��L�m&c�-+�|�6���̧�F.=���1`���JP��¦�>I�V�av����&�����o	�U�ڎ�R��_�~��<=�@E4&C��i��p��a�j�u�y/����|>��v����iW� �𫦙�d]]4g1�k�Q�ێ���x���4���t,�~�Dq�F�t#�g���%5l�F�-��ִɊ��;T
�����Eާv^��7�x�+4r�P˔��h݅ǑCX�Dt�i$ܘ�Y�����;��j���;�<���J��1ߙ�25�7��hX�����Q�ω,�c��5��|>���G�:��{Ď�Es!�cSe�O�(�d<�]q��{䄋����.���%K�78>n7�61��qW������u���B��3 :��Ш!o�k^�ΦBfے��q�.d�3�M�M�!���ˤ!��I�L�ސ�~XM[�m2W�2�ʳ�	�O�>�F���I��b#`�
H�W����i�*�ã`��8��3].���M�9���MͰ���
��^��a���{x���.:E�;��%�P3�\l���0�I��m�1z��v��jժA�kw�r>C`p�'Y��d�|I<�������D�L��
�ƀ`0�Fz�Zm�I�+v�)����F�O`��YO�2����t5F>j�F=�P�2���(|��?Ě���6\ugG�ye�i���ш��=��"$�a6����� ��5���oY����#`�|޻p�,�oH�0J�VyG�C��sS{<x��(|�P�]:�;��b[[}6o~v%a��IW�q����O���������酹i!M�bz��L�������۰�g8m���]����
�5z�B��%��H�0����A6B���A �Y��k��r�,^=����Si��◔��q�#c1_joAmU3�'������33[V�ܾc$����)���lm�S��[�m�2g1�Qc'Ǽ��44���D���uq[R�c����Sxu�X��b�e���m@u,�m�����t�a�:�DY2�'p}��Qt.�`��J�l$5����� �;<ǅ���L�&<E�p���).���]1����FF��l��E�Y��v�4���f{���GqNGtR'·Z�`yH�-�s?r�X5�h+o*�	
���5xֺ����&���&3i��?Rv���/�����f*J�Tr$�p�E<$���au�v�t�^D�9�3�q�� �e��[�ϔ[uE~�<��(%����3&f�2�}�mSp�v��w�ܙ���9�ʁ�~E<���kܓe"���^$������^[Ϧ"g+9!�_�Z���e�12��`���z��`����6��Tf��0��A�`��P�1S����mY�z�]�$ FNsS��UHa���f�X�:���j����r4���utԫ1s`_���n5l+X|�j/q��߄���2uȣL�͚�F��0����l������q�]�a�b���&P�'~��E[�wq��	�T`��uUl���ׯ��%���R�D@�ϵ��ۖ�Ӏ�1�7&������F�m�
xS��� 8��V���y�zL$��S�0<��I�Fb�33��Uj��1Te4�(�vj�"���+3��c?�J6��W��Axq��H�Wf��Ԅ��]�.ŝ[��_�-��= ���\M%�kyE�Ak�K�������.���������&��:؝�?Lh)i�;U.�}��Y�����'�n�[�D�rO¤��6���.q��vu2.�-(��H��(��=�g�ʹ@��l���� ��L�tt�6f�'�,�~�p}5b��JJ�����tTB�[=g����Ss���Xﺉ�F�b1�`-	�uu�3���2�Z���|6b��� �=��b^�*&�N��B��<�ሒ7#˵���?�%V��ӳ<��T>l�Z|� Hј�e���kF��(em��8v5/�k͎����(y6
�3#v��D
��^͎�#j�yYYY��P�䐑R��s��
S�Ջ�U�7��[М#YmhO��gΌ�c��e� ���:�NDyY��˦MÅ�ù�\\���m��- 7mA�H�4����Yr�y���K������s
D-f��K��6	C1(5��׮�KblFn�n01�|��(%9je�6�������^%!5����X���D�+�����,ᾤ?���`>K�0�m,�s]T�K8'f��\�tZ�H���Bz�%��[�ʶA�n�c"r�< ��D�%6B��`��S��؂5��E����n�^��~�SQ�5(����ŦBC�?#��s��G�����Tnʗ�J���pu����#[�(4��Ex�]��j�D8�>³�lL�+���"�h�D����|�B�������D�X��P�������9a���n|We�F�da��+��AXm������@��_J���=1��]�[?�g��^���� �}�����.�5��=��y�n���"5ݲ/S!��}��m��kD ��}���DL�D���CeuU���kK���;����19ݥ8�@�-�˒�,�aFM�lCi�s^J��Ơ�{xk������O��<�������~4���.�DY(`s���s�Cm;1ziE{��en  v�-WZ�TZcrB�1-��`\9'��hJ������OR<�ƚ9窐����*Y�pb�E�^�z{�J�궉�u�B�9�,�_��\�}^�q�m#eo�$z�>	6PԷN�@ّ�괤��H��j�:�e�J�$X�)h�E0�8ÒF��u��Q��qZKs�xQ壝��5�WC(/OO�4F66��?{�v���N�nlf�a���1�p�4�X��ȇx����$��ppuՌ�z��H0bl�>�Q�),J���ˏ���'�Ho5Y��Bf���`[���z�mG:��D|�َRݏ0��c� �P�>�*�CL�
㊅�$]^a���t�����()��i?�iN�-��c����?~r�.E�K��� `� �$�ϟE��vA!r�2�l������j��e���^�N�M�kE��ҕ��T�YIW78�'��s]����?�-�;mؐ���E�8O[��>�b��7!�o�ݾV��յps4�cmŞ��H�ZQ5��� |!��[�;
��![�c��6PU~�8��u
�U��S��3�Wc�����x9ZZa���k��������e�����8�ۈ9�o��9��h�Y؇��uA��ӯ\�rvس�Ѹ;㳒�Z������~��ne�"f���þa/�œ�*Fg���N�e��:���;G+�����vV��ʟ~�G&8�=���z+Ȟjh�
�m`P�&ƫ��ܧZ\�{B����X�H���s��I��A2��qS�_�ό>Y�'@;S�ѝ�Gh<0�����T�8a�'ħ^�6J,�c�wx���v��n_'h���K�(�O}���aQ����;��ow@��B�D�b�q�+��P�G�޽����E��UbZ������4�z�  �^ 73�3�#�ع�7|x����F�i�`�zM3ng�eБQ�w9�CbdZ�q����~���~I��PΓ��m1��u9g�5���	��R�B�<ؑ�����H�h7��u�w~E�<�� !���$Ƌ����4���l!��jo��GSccT,{x���)O�PV�$����q��}�p�o��nᎧ�!Ğuqv����Z�����s������+�g��f��ƺ�k3w�R�� .5F�������{�"��nK��d�C���5��ëن��Twf�AᑶQ���X�Wz�Z��w�T��`*o������!�#�p`�q@��7B|����ŋ����X��6��T�Ǉ�ʅ�==�/��I�����	R]d5�~�s�S��*G�,մt��Ml,���]��Rn�i���x޻� �@��(xO�$��xC��?�
��+N>����d�F����lݹ�i,fz5�\���_���DBD�f�]����L��|)''�	�JyS	���C�B�
��|a���O&�4�a$�}��^�IQ'����J��͑�b`��GR�>�
wU����wt��p�X���4v��e5Ht��*?II��7�̶?Pz]���ll"�
h
�1oY lTg�"���95ƹ�<`�@�^;kv��^W�M\��A�3n2z�Q$�?�O�*Z�SF��7��4�֕�Sl�8���_�mt�MCv�~��{m��G4?�}�e�O��opPݤ�C�O�e顇��#�Wv��?��昋��	�_�1QD祪��?���dD�fj��t�~8����|��n��q�>���u��ٔ
L!���AGky�QY�ME�e �����砞�k}��0W{�-��XJ>�n:�<�=�p���O�QB � P��d�\��q ��F�J#[�E��P�y���%ާldz1B�.v,�_T鈎�^ɫ�������ZЋd/!�-%D�����T���;+w��&�Ֆ5�D���έ��Q���0��>�v�Þ楩$ܔ0۞�"N�֜(1E �1�ˇ}}}�A>����0T�,�!�@�v�?6��.�N��%*$�2�
���{�2�@V�;�&|�tP�h5�/k�����Բ,�D��N�z3&��������Y�������B���]$�Ի8�@8�\Z�6Q�>.��ZʴH9����Z醡�� 3z����Ӳ�aT�n��ea�..�,���=d�x�߇�_6�#��y�N�����%�5�`4�����1�j��K�=��;7�B6>^�7U����y]q�8��܆�BP��ۻC��3�!�_-@}2�$�ڥ3���&�ɖwJ5WV����7�c=��K}F�j���o�}[�D�w��7� [�r�n��/B���F���d��f���p8�����= 3�σ�o@�	d�#��Y�%�3���7\��O���u�Oָ���^mn�h���YVh/�_�
T122��ɷ��A�f��{�ғ~��m?Y�����Z��+�I,�U=K$��ϴ@c7h�B6}2�&�q;���>��w�קԓ�XZA�f�ɪ��U�ވ�#�"y%8���ぎ���l;���켼<�j��&1�`�2�oh˫��^�k\�Gf	��0h���#o��vY�u�l��3h����U�����V-`��<�_�~��e/�n7g�[�A�\��í�?�]����Y�A���i�?(q����a�d���֭�Gy�4��ڞW%�"�;D��]!�;�Ʈ؎s[E�s���婜e�Rͱe��QdJ<�����ib�f�L6��P"@����b�a���]�3'OP�� ��G�h�c�t���Q�����q&$�R��`ڌ^;�^���&ʕ�@���S<��u!��?���|5��<���5p)�?K&IT���Av�$����o�H�4%�f<�S�[��9ΚU���@����7{�K�^�Q���}��LZ���^���r$��|v�����i�j���4�s��s~��4<�[��^�7��L�>o�(CUC���9:������0\/%;��Ejj� ���0X����>>>swf�!����կxx/�3�;���P2�zHi��Z^�܌f������˗��ə�A�gO�xդ�m�~L�� gr�4�t;x\K[֠X�s�2 �:900���; 37��v�$�9���S�6�վh��+����� ���ՠ7�������2u�-�ϴ�8��a������\�ja���0�_ET��s�%Kzy���<r����R�UM�{�Ǧ�9U\�Z���D(=��q��w��/��I��!y��#�)������Wo���Uq���٢_9��?PK   [��X|�K�?  :  /   images/8210dba9-ab36-4d93-90c5-eeae848c0250.png:��PNG

   IHDR   d   9   ��}   	pHYs  �
  �
܄߉   tEXtSoftware www.inkscape.org��<  �IDATx��\il\�u�ޛ�f�pI����Z�Ց-ٖ�ڲc���I�K\$�Q4��-P (P)P�E�.H
4HlÒ�8v$E�,ʶlY%R�(R�D�����3o�9��g�!9o$[4���{��w�=�|�|��G{~d�KY2�`��)�� �"����P��uݪKƒ�%���̝D`j
��~�u7�I�M�]*�2:;��D�����ї�R��B� *J�v������4N�oCGo�f����.	�ޭ�Kg14>�OT�3^���
)XZ�1�z�U<�3�U�iE����3qT#�V�tb"���,i�D�&.�������E*b�|0��I��	`p���,a]�pg��!����BtC`�m�6`7V����-C�if*�c�bb�\���z!MHhp"�r��H�{��
����� �*��5tNQ0c`�5�^�ċ�P�1(�˚���<-�t��@M׈�;VF�,e,Eq�
^��?��%�y��D�k�aM��i$����JSt�a�2|�q��Pmx���g"״ӿ�[N}��Σ�|k�RL�cMn����4a�]#
&�2�ۥ�R���Il�I�aEg���5�����2^��C���t�{"2�aG.��ae�A��!fϞ��XQ�c�k?�3�}.���g�
�4X&�NI�K�"J���b��t��&�R��;��G�K��v%-�[L��P\�ώ�νF�RV�㟞���������t����`��l&���S��b��!c��)'��<�9H�:����;;�
��'��	���4u"m���������h)OQ-�M��5���^X��*h����Z�[�YL��W9��j�*�P�q�
9jŋ��s�b��l�bN*�P���7N�|�iK'�,^�1�YH�ѻF3c�]1|go[v~k��Bow+j�ޥA�q�ݛ2+I��Ԁ�m�aˎ��E��wI$��#<��KU8N�#]�9�I�jX���vʹ��>�{<fj�2L�<�T�M��dv�h�&H��#A�UB
��۾��i���m�e!`\��cmu�۰������u��`o�E���dn2)ꩨ���_�.� ��mD<Dc�{��U�����=8v��(�g���}^Ϻ�$+������+gttk��ɻ�\��
	M"�c�c��ဒ�����9U&XpzsnR]^���,M{?v|N�PFZ\��T����/?�!1N��D�gRn�E��aB��5'0��"�N�yv34��{���d+ *�
*�3��i�΢���ue؋{z�q����6����7��y����Q���KN`3����ښOBv(�TB�+|��~7�d\�"�o!(2#�))��)!���V�M:B�UJ�	K�-
�П㤐�A5g`�tT��,q@�u첏½ E]����Hn�8r�,ǩ�Se3=�._8�D<J���KU��S�h�&0:m@^D��������*=+
ajj
	� �{4�SGhU�&�I�y�J1S�W'�8lB�h��ب����k���d�v$PS��ehtZ���M������TX���xh@�H�D
�)�G���ĉ>����-��b�ڵ��|���J�m###���C  N!���*z&4L�;���x�xf}?�]+GW�WX�<O��t�_<�]��?���-C(6���BD�d+z����eӕ?�BǗz\�4__�p_�B��HsS��-���|�rlڴ	cccp��ęFQWW'��-f:0E>����m"�Ǉ8�k�o`���	VJ���4�cI+�݄D�mu,�E�ɑ?�(�cm+��Qz0�6\;�{���t�Đ����-�ᩦ�===())���J�Omm-��$�_��r"�_���˧u#Fn�Iq����G��c]d!㷰B��B>�S�ô���+u���"��-�
��;~f��RyL3S�笨��*�"VIȄ˲}Lf��>�-��y,���-��iݺu`ٲe���Fii)z{{��S��W>�ah�1�-4G����:L��2�[˳1�0?�KY!�,�{�yrg�oI3u�1�ߵ��H�ȯ���g
gz�Ǉ��Jh��h���,� EF��Cn��C��P[+#�e�	����x�^7^=��gs���0}��[��h2n�K�� '+�n�O�v�s_F!Iz���d_�w<�zb�}�m�L]�i�N�6�H�{Las�^��� Ɖ��6����k�<(X�a�G[��[��G���J�N�P������V�s��w%�򦞇4��xd�"���a1��N}�2<ͮ0q�0�g�:���uS��o��u+7 4=�}��?H3u*�wm��=�"89�r1�X_:�7^�g��w�OQ֓;��`�|�H~�4MDSl�7o�������8�����ֆ������7���12�+�N�^�"9|�Sز�A���Ng.?���(�k��.�6��dX�]��,n� SO9z�B�Zue��ML��
�Z*k�aG����QgX!l!�HD(�C_�׋���crr��� _f��=A�\��S�jJ�������8�C!Y
�����"|(#���f��1����꼈�k�S�L�cS�<��##=hnj�0��m'qc܃��l��pꜹ�G=@/����[�X0!/��8����Nu�YHj���6b��~�r��5�1�:������
���_i{l'��'����c����'���^���:5��76TkH$����ԯ�8t��^��!S�C^?�6�/�J�I��V�&Z���QL�y��8m�AUd'u݄�2�IHM�9c�sb9�\1���}1���
�Y+���0��j�I���py`Sg���i	)�E&ON4�x(*���[&�$|�a7���/~)���+�[<��':El���Ԭ�v;��/��,`�R��U2q�����~~<���P�c*Z����J-h�YU���c��D	q�x<�Br�z�L�%��ڐ��3�d��������D�NP�rT"��f��g�)+�7�o�:E<$�ȋ�iO�_���}x�)k開9R���W��/�"�W�`[(J��
��y	eqL}v9��CK	��pTGRـ{w,�A┄�R�L�a�(��b�R9��K�	�:�6��J��On(�����GX�@#���rV�
�#N�i{��	P1L1�ojM=�ZS�����L=.c2$�f�	�&Tl��A���B1I�[�DV8I�W]*�NqD�˶�C:]j���F!�n-"i��<^�9_�P��!���{�o��E�4�#�p�e�S��1�ƎSϾ�"��cxv���cYL]��Գ�f���L��HX���������:I8�lI�5�ۚ�輢[V$���"��41,P1l����f���~/3����w>������ԯ�2���'��u/6m���k�ޡN�d�y���b�|F8�L�*��ܚ�+�HQ�dV��n��C�h/�:�HHs�a����k�k2L}3��(9 b�W�0��-�^��.b�!�L�s�8�S�۶4�c�T�d�آVYsNx��2w�|9�n_�L�o��ϑ��\ԁ�ky���p4[T�$�ߖ���`u����~op	Υ���L����i����2�vb���[.���b����=���S��@r@�_CE�,L���
c��7e�}C�K98����:��U�~�>`ny�,}o�v���כ|8�❻�A�v��L}������Ś�ś
��2�O���$I�Sk�t�8h���Z&�ԉ))�F��b%�����u�H-E��l`r�?���@�8��+�x�`΂X���y)�����G�ig.o����b�gM�Zs}�\��X���kK����<�� ���_>�)�����^b�.��6�:��{\ؾ��
Νw���Ҏ0Qt����M~�+6̵�����9#��w�s
���8#���:�S��[T�� /\�A�"��n,%.d�s8�o���^��=��lhY����cSm��0��8��s��FL�� ��E,�k�H�N��hO�����
�Iۻ6D5)��k����pb([eN�����VT#��V	�,�ld���2����sp��㗼�-���n���`.>����d�G��3	9�MvE�[{��1�$�^-��١~����nii��ѩ�HVf���Q����1�ӓB^�3\\)��"8��L�ڶ�Bǲ���&��
�YS������r03���T�����yI�^���C8���ؾm+zk�7�n=�!3�%�
L|g_m��V��"_署�?B��<@L=7��N
#-<'��`�x�dQ���{��j�$|�7���~�%���f�S@�8�ѹ���9�Z[�DK�V�VcR�?�y����~dsO�J`��oaͺ����7��Fp�_IH�);&���cϓغ}?����q�PTVp��`�W�m��ԛ��X�N�!��$��N�ʀ�s׵y�է	��Gb�w����̄�7{?+�0uw�
ce���y���bY�����38�:��L�骚����s�wiy5��F�޻o� �4N� �b�ǋZa�g���c�<r{�����L��X�ײ=���X�ǩ��Ia�l�h:wDN�M��H���oR�
�n��Ŕ+:�t���5��~�!��r�k��@_O�`�-�^�ev����SoaA��X?Z/6����b�|/f���L�$9L����
���� K��u������|A�;/�?�+-�?I�ra�����v���:AVbDFd
E�o�{��8 {���.�z��R|xqQ�9�X������N�q�Y�������ݬ���s*�e�M]�+]N�r�h0c�Wۨ�{�؞r�盜x��4d�W<A�����Z���ɩ�{��EE������4�Cq1��7�xL�9���|�}�W�'/����mI4u[L}z Y�Sg���GW	3u�a_T�Rbq��è_^v[^�dK9r�*Z�F�BBv��SwQ(������a�_>�tSN�1�����0@��TZ��a�t1E�xvb9u�L'jȖ��}t��Р����z�O���d�c��~��_xɉ+n+�o=�sj�۝ضJk �T��^�S�T��Z7�e1���%���2�n�⭋>띚Y��;�j�o�x�rRXH|$U�)l�7�"J� �Й_T0u�2���\Ԯ��"���;(�_�	5���(w�,j	�{�6���k�/�.Y�mw��e�#�Ǩg�-T�^��b���r_��UYb
�R�8�WKڞ    IEND�B`�PK   �<�X�IM��  � /   images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngt�P�M�ED�~�t>��J��"(�= �	�C("�T���B%� ]�=U:�C�Pn�����Ν;���{��s����Gm͗tԬ�  �N�� �
	 ��s�*��!k��u�Wƞ ������r�}  n�ʋgz~ikxH,;1}�p�'���tn)E�EG;��ſm�3��ͦ�+m���0�΢��d�T�O�B���Țq�8n5���t����!1w��?�#��M��έ=��ݟm����gv�CLŻ�32֋J�։4���VV֋� ! l��!m��)_��.�[��]α�S >]O`�_~(BiJl#r��lI�.� �`֗�0W�a��?ư���+OϽ{Q�����1\��yQ�鉄Lc��l~�}�(	=>\8�(��z画~'w?pt&eHCwQ��xJ���'��XHP�F	sI[�ܛTN��n�e_>̎�8iHLv;��+f3�W���i�tU����\� ��L�o�"pUMI��Ol���@Y���;#o�s��Ōحj8���.aS����G�Yײ���6���)�*f�r��`��������_Z��#�a\x�;���������n<��㛪�k��k@a�����v��@��Dy�]d��PUrֻ�����bJ�/���>����k��c=��BV�V���?�N�=g���#�:�|.ƍR���P�t����B$��9EҾv<�4$�On����â�gP�ֈ��U��o줼�ْ֙���W��� Yr�
��U��2�߂DUͿyv��L "�H��+��P�J��.>Bm&���N���&��ff��c�a\V\}w��<��A�����|}",0��K*2�����k滠4��M��7V�E�A�b���W��CH)amR&R����B	���M���3[<(Y�z1]Ǜ���F�,����\R[���J6���2�&T��,��n�]��%`n�w�4fB\�}4G��7۔�+.g�����k��;�˳��!�W���mQ`5���ϟv�f��kTB!�̄�	��Z�QS�e�~�s��8�����e,�3���"�=�G�;����C���1�\��3���7�i@@M�M�	>w��k�or�X�K�0a��-/iB�Kt�	�%ai�J��W� 俗��W��;kTY�<����H�T�g�[��VS<Zeֈ֓*]|q�F
�����������obE�|W�"�wD�Ԙǒ�+�=5{�n$��Y��{7hl���ͺ�-z�N?��3��?�ܰN+H��`i<y(�y��^�R���"�±_?�w9�M+���g�2���Åg x�����ٙ΋v��������k����l�eD]r0�i����z�2���}�&���]�k��zw8[�~�DRa�K022*���M.��:����S|R|�]%��x��8۔UJ�&���(�W�����]���A������
�	���"ͧ_{���m��{�	b��\��999c�$K���vsf��@śN�nX��c	q����U� <�m��S���������FG��ة��iҌ#օ�q>������q���xT�0��SQ����Sc��YԔ����'��ƭ^�8>N��-�rF�_;�F�)?o@|�ڴ�h{S����w�(�.͠�T��񒕀ُ����_߈_�`��?#�#��z}�V/�/b��Z4�A�%�`��OĉU�Z#A]=���Qe(��A{�� {�nu@<����莮v"��2�Kr�x䱶������Ӝ8yoε��V9(L&W�k�M�r&�D�t�����TW�&�"M{w�\v� ������*��Qm<����2�g�i���wS�G N�[{:Ϻ>�yu%N��k���N��V����F]nI��^Ҹ���3ׯ��~R98�l2)���"�u������_%�����˞8�2@hkԒb%ĳ���_$_�yD�\���/(��K����]N��`��M��o_������X�#���k���G�.E�;�Vʠ 3+G���<;m/H�!{�P��I-+�Wפ%k*e�wih��-���	B��;خc�jD���}����?ybbշ��깠"K�u�J54����-��7hpѫ'�Z�ʘ1�ԑp˦�)�T�&+u�/�F�y��
������7����%H���ތ#sD���rC��\�\u&��'�|�����m�?����[����t��kN�f�9%&&z˝&�V�x4i��bT�^����^����>���:w����?��!/K��j8P���㿹?�&b��=u��	[�<=]��T�᳻(�.��n�YA�x9�{��a���,��Rā��/��|ҏ�˻�+�k;O/��|'U���</��h�J��o��Q�Z���B�f��b΍�A�NfF*�4�f����Ir"ݹF��F�.tX�R�>�1(M�J6�QE?^܏����<b>�]-��)���պ4�%9Y�ʤ��?�߾\�4��a[w%�UD��q�)+S�z�~k_9?�I<��a����G��Jᖻ&��q$���L݂�_ªx_f�BW��"��7���i���*��OX�K�,��M����f�3%�#-�:��3�������B�a��Z0�P%&e��8���Q���h�d(ۗ3��2���#�F��#�[:�El~���e�o���L�G����2���+Cp�zP,�>�^u��e����,�Ӽsݭ�X��.3?���Mx\�~������թy���5��]���F܈��U}-Is9;d���I���q��B n>���7:c)�P=�e��_�
�?v�B��K�<�w�����L�M{EN�� +FF%��=h��Ν�]�tN����<r�y���gha<�We������/�ؙ�^n�~&��t��m|,��pך0�[*�zeZ,Јj����ږ�0������`���G��Wx5x
�9�DO�}/�ǥ�S�2~��Sm�����F^��`dpc6���7�m���F��ݘ�j";�£�#��3�֩�oa{�.�|)fe?�I���7�m,�}��,z1�U�i�ľ�����!Kjo-'�j���)�{0�/W1Ex�ğ��}Z璱�^�F�|�����U�,`0�7:33#���E���f��x�T����nKU��т.��!X2ܻ����%�ť����?-� m<x���k��6dJ��!T(�.������u.##=�cXG��A"(W+�F[[ M�����;�����U��/��P�ØWI@"
��#�ݝ\5]���1���#�^65�XZr?u"�OOO	y�^3�W���yZ֚��6+���T��ZT.�Y��X����Xsã��o0�yD7�Ƶ�,��bXȠ�kx�tT̖�<�Qe����]�5��/�U��ܾIr`6JJV��P��s��Hu����k�$���[�
�s��$n�_��r��!^�$	�F"�#r]�V��Jl;���|�2j��zy���]ש��#1�b�!w�3�B��j����븫.%��d�S[��;�����u_��٩�t�'ߚ�4������;���2��^4߇��=Wk�A�Z��4��K�$�<;�&%W�eR��3���>+�@J���SL8 0�0Q�%������Z��L���V��o�9���>Cw[���OOT}E� �I|��p�u1���Z��}5�\�7��y��_0�3��l���Kf�TK�)�����3�����g��ݱ+�'OV�S�����.��QS4!,\����
\�������,��9gʡ�G�͋�?|~��ZT1?�x��=�`xnLKni�<>dbpz����B����{a�[����d�Cv��(��f�O�'�1�؛Ҿ���-ҿ��F�E�/��/��?hU;���QvBP���'=��|���X;���v��I49��J>��d��c<�ݖ0gRgv Cs9���m�E"�������R��Y��-�[�~�/AԒ;��A���~Z|��� 5�[��<HWT�����Dv!�Q]l�_2�?z�=�W�Mu>���4z2��b��元U����g�T�/�X��_��G�˚L���_�ƪf��=˖d]�o�\��?%\B6ʅ�E�@ �$vp0q�g'���?�N�L  ɸ�-��?,j�����P�o��k��QTj�\���'���\]XX��L5@�+�R���u8��/B긋����$G��͚�a�������ԟM=�:�G��Y6�{��.�~N�nd� h��?���҆3r�Ռ���y�LJ�b&}R'«S,����yH��duõD�ń`�l�����!���A��I��)���ߚ���q��@����	IdR����\�-o������y�]Ҟ�zE��Yb��*l���|G��*!=�A�8G��7}�y")`��<���Ɉ�,$�IB.@�
�z�>�:��u��a������w��ﻲMS`ك�l�\M��Kt>G�hŹӼ�"�x� ��ʵ�qbvd�rJ�����żu�hٺ-2�{����	&c�����_���c�cAT@��Q��|e��?y)���憽+������!������b���U���IaȚڑ�9+��E4-��Z\��z�]�E�(E�-i8�r�7�)�+|f���F��^�
\�Ԕ׏�yJ2{�C[���g��-6 ";���s27�;�Xs7xS��[�[�h��O��j���J>��R�'4���dzs��bAomqV�H���ǆm~�ǌX��ӓ)�ceBT+)uS{��ۤ�{	�}�ʱ[kr��f�i�x�cڂ"C(�`3��Iqx�y�%=
Zrh|�ED�����)��o�)���=}�Qr4�ҚSh�T��5�qu�^kF]�H�������6݃+�w͹&W[ME[-�q��s��`��X���܏3Ԋ �}Rn75�7�W#$�8�	;�z�%U�����JO��v��[A�g��]��	���4��l&|(-yɎΐ���'�ޟ�e��*�K�B}d���K(������������q��z6�X�Xv�!����b������İa@O�_`7,`|WϐT���t։�!
)�4V�d���£�>��ߜ��u؃u�	���
��*��X%_uz����KWT2�.�G���f�"��9��.1�COR��z"n���#�����ɕ&����f �Fۀ폠X~8������K��2Tp�y������c]h���n�ʬK5���5=�7����x����1E3�(
�b��]�3�B����B|�N�e�����VRώ{$��h6��!3�:��f���3d�C3�*V9�)���e�Хp���Q�g�>gux	��e'�Dc�An.�����o��~5���.G�a�����/�:�S3
\��	) 3l��]2j?j�H�ُ��XZ]�2xV}�:�=3�b@���	^!�W4�
�˞5#�5��u�����N�!��%^R�ׇ�¹P;@қ�����ۨ���1ͩ���ƾ���JSZJf*	VLI���a�Ѱ��q�J�)_��������C`�\���otú��ho(��#"��n�Jt��T^&��+7ƾ�n���$t����&ER/�>�HO�\�Eh0��淟UI(�I�=��c^[Ð��Dw�{[T!��bk�d�F'��Y`���_5�ҡ����H�"q&a��4�,[�0�a*0��2�htϓ8 �l��������z)¿���K�#辢6��ݚ���.ݜ�+����ևup?��*!�E�R�ˇ�W]��ee���M��{��5�,���3�s���3�[$��8��%�߱�g�5${\��'<��0'Bhel���1���W����L��Cږ�s�����~t�~"_28="W^�k�j×�o���ع$��s��%}�P��/+,�h4�Y�Y$&���� Fn����I]�n:���,-�x4]R�W�5����_�^R����fי}'o6	@D����R�m���y�<�dI?����Ax^Ĕ���i�D�N���|���Jޝ�~�?�/绉U�Vf3I�ݡ^���N!,�yWVo��͖u�N�/v#EA12O�Py-��Z�<�Wb�?ڷ�T�N~������kgD�a��{w�).�������9��E���f��7H��o�R�ݲzt�U��)�ƽ�J�"�������&h1�����O��l���i��Fo����
�{>���ť����X1Z�O��Y�цE����\yΓ�w̰��&.� ��G&�K��ث�@M���bB)]��E0����3f=좓x�,6!ˮu=_��dZgU�s��}���~D�`/ �O�u7J�&pV̊9
�zS�i1cnkf��WU�Y�wt��f=(!999���X먨(�)����i	�zj5�ͩ2�m�t�F�Q�Q�AS�;�斿�A���~���z/ַ�ʻ�1��)J�=vb������Qtp���gq���߾i]m��|��Le��)�TO��ݽ2V�'��~���퍛`��Ŏ�p
��6��3%�yZm��&��u5a^�3H�pZ�L1;*ڻ�Z�������gt�k����n����y˜3��W=���Q�d�^h�!x�����9XA8�$g��S
�adw��m�p�dw�Cy9t�dȥv�T|(i?�3zf�4��KtAW�_���F��B뽏p�G��X_��Ί�F���]������]-�&����\���ҋ��ME>U��Q�`bx.�#��._�$�Q?�ԨC�H�`��zi���za/�7?�ߨ���<2��)��>󊐡A�{��	./��Գ;"����s?A�܌��͌% �ïfntgʷ q��ϟyZz���N����L=��́A��R�e�!6x��ax	C�H������n���K��j
ds&��'�nb����NSa���[�B��䝶���B,�з߯���h���A�Q���d�Q���Z� �̊o�E�|��?��GD��e��Ų�scY���*e�i��ʑ�5�~=���)������Ň��^d��%L���S�^X�]�"�>������0�i*�R��X�h<mG�+5�����uՊA�B'���+̈��Z��$rt˒9Mf��i�ɕ$����]�i��4�H]&L �]R�c��w���d�&qI���2�@U0^�
�yA5�0aF�,��Cn-�w�#g�l
��Z��L�R8����;��T�>�"3�M޶2�����Y7���wwqI��Af���
���f�Enʹ�3`�J�͵�]G�8�HBs��a:��_��_����I*��uO�<��!a�-َ�A�FB����W�q���3:ۯΐ���v3����
�J<��� ��u4�c��	�Q?�,5d�PEHt<|�����*)��Mq���3��ҵa+%+��w��3�=�r�Q���N&!Y9��o�ƾ����5�e|��.��rf�]Yl̻�	k��o��gV�M�սg�Ş�&�(p�fXI��3��  �6!���[��,A�O���G���	��l-���Q��8�v�*iD��ҷ��]:�~��0h�$f���FqCPЬ���.�E�}��YH=D��7����+����|��'��UN��0��˘>B��g�!jyz�jk�{A���QkqĜ�����
�����T������88��ZpHE����1?�����@zU��-r쟛eu4&�\�jF$8�������b�ī��x�k.�Q�E9�y�-ε��<�	l�ϙ�Q�Y��KCƋ!A��7?��� �j�p��,,"޻Sgt�5u�w�LIT,P�P�u�T(��/��c:
�gqEj��֊�����Rr�9�D��|�r��FF{Fp��!MUE���
&)B���W�YG<��cx���q�wYX��2�;3��m\�QmY���b����+�y4dq��3�"�f�e^.�aAX`>
.���g�L�6p�Dh���m�q������^\o��� �s,�EW�=#��K�`(S�b$��2�Bv��VW��n,�����p��Q~����xg��ƴ�T��+��zۃ?Ͽ��(  j�/�r����h�&xC����\y��%��8X�f��+k�H�͇��-�ܘ8��?�R˝��xD�6Km��te>�|�m�T�Dr��?�|1��w3�4�;c���n،"ո���\���	�U��ĕ�>$r��^�&'�<��"֜2��N�G�|֐T������w3F����w����l2s/͇�M���}�'S�79�)�1oi4�i̔o�ۤ@�[�U6�Q�KI�$ܘC+���� w5!\^R�"m�$K�=��:`YY&�����Q�*[���J�8�͉O��T����>Χ,.�ppY6g�ӛͅ�R���B�	l����Br�8>�wR{���(��6���v<�x���H��"_��l � ���"�����֒�|��'p,b�P��D~b_�5��"�=m)��gh�ܪ�1���\^�(�X|f ��t�ʸu�ΊZ�d��a��=�9 }�M:�8��8,���:��8. A�Sg�u�Vuu�Z)�/��u�g�~BekLW��&$����.����kՙ�Ř�̦�H<@�E�S��9���b��l�����A�'�F$��Q�M@��M!X�rt��!}��x&֦���6����+V?�띣/�j{��Ѩ`SQ�g�B�<8(�n_C�d��oe�����Jy��b��3C���Օ�ޅ����mc���45�(p�S�r���κ��4��z��VB�>�����r�r��H�Ԃ.M��������Z$��p�3�H"���%nD�x}��sa�:T��ۻ,��<!��j���&�%��tvvu�z��Ĥa{/���G�-%hRi4�9�s������1�'	��k+J�,�ܩ���*�I�+�:��+i�� ���Ͽ�j�?���k�#�p��R��&s�>�.�l~�=#E��M�vk	��g�X���WL��|VzLE���`�ׄ�ce���#&����i�19od�dUԆG���Uڔ{�L ,��F����^����-��coY���+1�
|��6��A��'q����~��������Ay�֖�Q����҉7�=d��`���h}�wz����Je��>�M3��X_��!'\�c��x�N���E�Ɔ(����wJ�N��)��8�t��vH�Ը��U�}���[ٗ�T��h���	GM��(�	�1�X*Ze!����[[s�i�
�QV.9���?iʂ�� O*��[:|��=DE1���
�	���!��Ϣ>�ۣՂ�+�º��ӛ������v���B�n�u}�%�?`�Xֻq�����i�P	�c���ս<V�܎��ʠ��$x������Od=�S�K���q�Ay�3)89���u��U��?�yO_u	P���;���q�FxeF�N�Ȼ�lb���h����x��I�ܑӇ�KΝ�OW�cU����u6���T��5B/M�V\���e��}��M���i�	}�G;cL�%$0�1��V]X>\�A����o_KP/"�{�ퟎ�%�t�o�mG�9����(v�v/q=t�j[�ˠ�xJlQ��|��ٮ��k�d�9�~�����@��'�/�=�?'S���|gVfo{q���# �d(�H<=��~�V8��u��h�%���Tk��������'����ϑԫ��ň��v�:W�-�}��=~�A�;�aT�"��_��#P#~rdj
;4����FJ���Փ�t)�m�teZ3akl ���'�/�G��;H��}�Ѐ��H���(UF���K>���ŏ.Ԕsu����]1/ž��$[�����A�F�ݳ�����q6F̤����u<�Đ�3`�2_���P��h�3��
 lsõۢۯ���+�f3[1�����x��ČyL���?`�sx�,���$v�erg�l'�$ˈv����[��+D*�6�\�p�KA�c��򯜁�߶�=�S�1�P��w�( �r�K?1Ì�0�o�ū�D�ӟ��}}W�ژG����y������� u�jŻA8���jߙ�NJ���z]�'}����mj�c���颉����s�D&��͎����X/��.=��A]���׶ݳ��w���d�&�c��#�]ȶ�1��<M����o������1�-h&��ۻ�3$���f������2��7��η���pI�9��Zl�E\�����i��KAxp����%��Qw�qE���|*cfZY�k
n``�
^W���@��3�2����&#k����%�Ϩ(����B��KљK���"��B,.n���\娆����c���޹��m1��9ssJ|ͣGZ�������<��N��a���0�.��avz��^#�����ݘ��gdOt'?c��!�H��p��@!@���G��錄ڵb������ۉ��~�l�����Cc��b��
��ӯ쓛��	�v:BqYo�$_���لM���l��'91��u�=[�+���J����{F�(��愂�)�,�Z���/2�(�4�V�	]SX5�f�e����9��EJd�K�S����.���9�*�!�T�:ι}�DX���k�����=��屚!=F]Ї���v|����zv�K ��2D/��� (ة���-���8��yrM��A�r�J7Xʳ���LL*(���ڿ���v9��- �������;�)S?�����/��?�7���q��������"l�@1�� %]�3鷩Xxٙu;�x���>��)��%��l�[.��IQ�E'��������A\	ԗTR쎤 ���ۗ+����\��{����������YZ��5<Sڊ4s�=����^�'���Џ#98f���.|k"VЀ�ZCs��`7zy�"��d2����*��7���ͪR��C����V�I"\�kQ���˩�5L��"�����v^puw��c����&^7�]����.��"\8��o甪u� �������;[�\�cwoeO�{�?�$75aA���q�n4E8���7��u����^�_���Q�$&v�����^.�4�.w������	��B@���ڴf��+�Ϫ0]�9�@�P�
�l�̉�s�ʟ�����n������]���ȕK(�B����>�!�y�w��6!x�8B�{C�,�Z���j��/�W���W-',����"�:��ȼ]쁂*����G�=�{�*�2�?w��b\�3e��^z�#O�o�y���&q�+�%M����gq��W�"]�WW�2P�HF�)��(���1�f�U$X����6��e�Cc#��x��g�������D��*9�����ۼ��ɼlil(qRTrxi�H����<��_7��!�nV�rrT '�Z|#ь<���_�C���V4]���;��Q5�e?A\	��85+ҵ�l�dۊշVp�W���]���ف9����	aX��S�q�	�r���a@@ �#I�;X��ܗ�=Vͣw���r��*��ߑ� ����ܩ����o�ig�*��[�X�5���1�1�I!�Ͻ�*�nt���T��w�u�Kz��T!���G.dͩ�˛�&,T���E��{r.���5��`����1z�l��"wЧ����7g�Iߘ���GC$��̈́�ֵzK�sSG�s3۴�ӧ߯�M��Wn�� �oR2��N�{���&����i�1��L�o=���^i��=@�Z*⎮&P޴���lsK3w���^5uRW@�i�+�hs��|��$]�m���ɂ�>M�"�9�U�U��ֺF�;�p(�*y�!/"B��f���!^0`�m/|9:�W��8i��5�A/��P��l(�rOku)t?���4!�i�HϱiHC
Zc({�sb������F�+čGA�M��y.������}N"�$+��,����:�t����ְ��n��{p��$e@��0eq;���>�j*�F������P� ��A��
��(E�v�+��G���\�?��=n��2�<<4�B��O�N�o%��t�#O)�ޢ^F(������Dd8�=j��s��3����m�c^�6Ͽ�`3��&5]��㫆O��]lqU���M����g��c1@�_�/°�8�5�*�d����M ��0�O\@z�����O$�2�T�V�SΓYKHc䲬����3����=x��6ZN�9�=�ʘ������(�E�R�'�fOE̵�d����\-6Լ���%����6��휀�6�l�ؓ��α�s�GV��7������J}�㯐����Ϛ�=c���S�{:��$���`�|�Y�>v�=� ���ª���ιo�#��n��斫�SBLa��"u�����?N�<��!&C��O��z��dTI�B+��w��W2�jŁ!g-�^}ԫ�
F؛Q
��=���6�K.�0+�*g�;���'�<�f�>�K �7&��!:i�3�K$8G�����(s�I���+��)9h���򯆦��_ ~��&���p'��r��*�g8vn�KR�y6x�j�;�������U�M����.1�nƇ��y�����V뷮�0{x��9撒��rWc2�?m�1B���ۗ��ub�a,� 8���\X �I{\�k#zKU
`���Q�fX�?���o}�^�B���O�@i�sA���MA<���#�W:��=��f���"�mu|r�T䝄���c�{ބn\�*�zE4?����\n�r�5��^m�z������`7�4Dި{g�"���������4����vKy7�FC�N�>s�<ב�*[�H�ɣ�G޻xhXw8�5�naY��ԾŔl��g�fR��{�B*����p]8��vc0�c�I�s�8��%�fG�[⪤6��fi�TJ(?<o�1۷{S���c;S��Z�o��x��2wQd��t��ӏ̯nG�u���E8R3풤�=��ܸ���١�P�n���ц�`i��ԸyfϢà��CxO����ؕT�*�P�D�
NC	|f6ɷ�QR"�
M�`Wg����<����fv���h'}WmMW�Պ����*+�gɐS��B�F��z�}0���v�t����z�o���l��M9��^�����%���������E?����e�g�����6��Z|}�X����3zNQY��vS�a�S������sMGUģ����-������֭������VS똣Mi��A���z	YY6�oPh���Ij@݋���K�����{���{=� 곆	�������fr��;|>�����sm��Q���V����,.	k�ג�%�̩h@��PS?�R���/䀬p_�ؼ%�[�}CԱ�W�N]�)W�"���©��YB�!{��Z �^,:��*㻮W��G��E���LA��<�B��B�ϠUF�WN�NX�z��BUy��]���ƨ\(bբ��T�[�Н�	[��9���[e�cͳ���9=-�FȖ��,C��Iţ�:���qI�g�< ni�L�~�Y�w�y��ʘ�~}��K�R�柁����|�F�y�OU`�aA�fH�A[���	���b���Ծ=���(����m���K��K�g�q~fM���)\�r$
.a������$��ӹyɲ���+M�m=��P.R_U�[�a���v3�է�Fm���T����"x��7����W��&o*���G�zx�o�S�h뽜^8,Ƃ-b�8Y�0�a��H�\;e��lF対��iV�>&��Ÿ��;1���@�?i�+�9���>��#���7h�%-2�[8����SgSk��W���U�Ee��nd�5=B�X䲂Œ�!t�HR�Vab�EI	={X)�-�#<��V�xFC�ڤ=a�E?�X2H��;u��wY���tv����8��!g�˙��Us!���R�OG2U��m�T����u��j�VLƑNX����)/ܧ"��aI���%���^�_ʜRG�1�ʵ�t����=K�"U��h�B�oZ5�6:d���J &-��KF��H�X��ZLY/I%��稱"WA�Ī �G�FQ�I�@z�|�ƔX�üK����>
H!��#��˒�A5�0w� de�?X�:�2v�úueE5��`�R��O���_jFF�Ǐe8��Ԗ�u�b���A���#��z�4ޡZ7"uq��]�l2��#�G�9�W�6d��E�-=�K�TV>��/Ԋn�ܞ��"�#"S���t�����y1��g�k�f�&:��:�H�����h�B��R��w���cg��f|���7?2YQS�\��no7(6z� ��3..R��u�z9g�o�:��Z�<1�|���̱WaGo4�e�P��KN`ro�wC`ɨ��tW�#�J�
T�jC(��
�lH�:݃�uN���L��5GQ/��v���6��{mN�	��EG���;	�ŕ�P���֬TM��U����2Yp	�phiu���Vݩ�GS��Q	�td0"����_����I�xP?d����[��t'�6+E͔�U -��l��2	�ˡ��[�'�'S��了!�}w�/�w�t�����m_��"_����7� 3Y��� !���ʑ�r#P=�~�B�'p��P��/[�	�l��FNM���|)��Y�Uױ�灐�jtr��<@7t+S�Jl2��T�.�z#^}���wsL��O�Z'�8���s�`���<�x�շ羡�UD��V"_~�ʺ:~ӡ��6�I��.�T�'U���\b��b��X�5E��E��ӓ֖xw�jz۵l�0�Á����������,T��TT� m���+@�����E׌2��d��ISW��1>��KKރ*�^��6����h��+V�R�$�p�Q�1d�9�)��)� A)��냁VS���ဇ}��'}��K��^t�g�"t?�w��
�5���#�;��/����Y�@V����{��L�@�NR���u���������W������\�_����y�^��xt��"v�
 �]���/��}��ywl�>*���us��"��f^hi�2�n��5����~%���m��+����;��'.��2 ��^�b�`U�jC{���<��<�<�-�3�ⶵ;I[��u;���C�����Y��e))A2���Li��-<C��ky��b0�9�/Ä)k��vꞱ���'�C� ��YA	�o=��A+h��lK�@"ָaO�j�r�PBg+V�-���? [�w�N�g�� 2c��z�L"��8ӣz<֙B��P����g����#Z=ߩ�]]]�� ��H���K5�&��S�n�g���g���YQ�9ʣն��F��1��tnʰ���.��R��!�\u{��D�KK��-��IЀ5�B�L�������&ʣ2�T���)L2���x�@G��L�?Ϸ�﹐�qXI'tt*-�t��]����wq��*��n��2��d�+��1�%���� �������Â�󼵷@Z`��B���ު����H8�����7t���/eR����T���|�>*��!�W��$�x�@��M��&�4Ҕ痒�[�������g���A'���Ru���2@f�g����^�#dSðS�%W�am�<�
n������ m��b?��|�]�_���{��=���e�����I�V[;��W�8�D��&�e�[-���T�Css���y��G��>6���G�I�B]�]�������/�n��~��Y�¢�h�E�7y� �'Js>���}{U>xٓ-B[*�>�6Z
���D��L��`9�K8�8��&%�Kv���{H�2�l B=3>@.
�M��?ww���. }�I0Y���Ń������Xv~y��l��Ez�j� �9��1-_��ش���K�_��p洯nd�2�#&ί��k��S����ps/�`P��ϩ�E
�\u��3��4�<W����I��gڌ��JU���*!6U�r�K���;t�[T� �]�A%3d(���:���7�w�6{�	Ts�82ݟ�^��7"?�G������X�]p�U�P�<�
؃������2|䘶���k���A�������#Y���ӓ��'�h��ʶGX�g�hHi���d�T��q�(R�W��@W���w�}��?X@��s����bǎ4����vk�է(4	�3����>��/!��O)C�w?���^)�pv9�QT��X�Vg:����H�agqW�UC���)��$�=������R��IE�L��E'���8B��	�D��LjF����1���?-o��>�a�]���"-c� Q��&a7a�,9�H������E=���I� ���͹G�Qc=?���ߙ��O���E�=�Jb�29����h�-,3��<�6�N@!0�Wa�OJuo�5l�d%]��n4��C������|��w�B�8�@�29�mDN\;�������3'�H�*S	�		���d!�2��rk;'�F���!`�/-����^,ϟE@���
�"��[�7+���[%@:/��)L��0s�O�ݧ�,)�b��z�r� ����vi��A�f��Ɨ��ᶉ�\�p����� +Gӵ���9���J� g����X�i%T/��.ɘ���(�?�����f��n��������ao����OJ��B��.��%;yG%�1ٳ�c�k(%$�:$ی}��6D��}7�R��Xg��o�?���|�����������u���:�\#i*WlW�W�ΐ=�Kp��K��:�A+�k�2O�`��Ce�9�_wl�]L
̥^��on��q�f)��J���ԑ)@Od��c��}z�S�F=͑�X���r��s�@m /Ņ�2����ъa�1�F�(�$�V_*�SH������U�987T��A�7�ʋ �5ٽ��K�(*�3%!.��w�d�������ꆝv�����MO�Q�`��Bb�i�M#M����ktfۏke�b�	􄸷�3����=-���i��^u)������_���ǟ�����_��p�ݲ,1ЀM6B���嶱v���gG���^�,��<����`L�3�Y��%��ÎO^>|�K��'�s(�P�������HA,��qZ�-�|m��"�K�b}�\ �M�����	�V�����Ϗ@�A��~���Fn�y<����t���Dk��&bz�$	���!�X��Yi-FZ��R�a���J�
ms���noyt�At��L������,��V�߃������֖_��zv��-9t�g>�<�cr�x�t?R���J�,Ò7l��a �a�c��
�aN�3�0��
��_�j"�V��s�j���D�av�F�J�#;�����n�Rn��k��{���\�� ]��Tζ��W-�w����.}�(�u���6x�,��`�U���w��_�>�$���ΛtD�S����~�t�Y�G�uKԍC��<�uW��d�,]��\��Ϲl�b�������s^$���@�7+�:uMM��f^ߛi�7��1s�_�_�;�Uu�����gb��� /#qyS#ϴj���:����ZS������0���L��L^����Ҩi�YC�n��l�Z���\�nz��އ������,G�^�n�ؒW�0�lC���Ք�c�^��v0��$Ǖ�{6�^��o��F+���xǵ_���A���� ��_΄ e�=O1]�w[��y�QC�O�l�&�_0,)��`Zm�97cW	���o�4�����c�V��L;��_�7��͸{T���f1��?h��<��S���)�WeI!ۢ3+D�R�61�ѷ+����7�/�,����)���'�;�� ����̕P��z�����_s��mY)ȭj={7��Wߣ�N{�����a��'�4��OU�ú�6�L��QQ��3��`�z���`��"�-r����k:�8
F��c�.L�O^*X��u�f�8O�b�[fǓ�r�^Lb2|�ogLx��VIڀ%;��<�rN3�"P���m��O� �x�ZQ��);<OѦ��H�<���S��]�>W���fQ�r�`^�=��N���|Ԁx�ς%V\���cM����'�K�ݢ��f��,����S��t��B�>p�ǻm���~�S]-;&W���DgeЧd&yt^?��������"�g7	�W1��{���z�F$ai��H3����
c351���\�f�������H��þM������kM]�G��Mj�v�Kb�G��8�Zo̻�a���".�U2���yw�MF�Y��^�o�;3�����偛e���bJQAyY���&/M��?�s�؟-�k�S�j�}�r$M�����r�W�p����Q9��}�HM����=�z� LD��*�-��`o?����2����<-MV�{�������z���A�u���I6=yw�z���)�� F3O�(�&||�/)P&�����j���F���,��+�L��}���}�hP�yO� ���d�d�qDo��  ɾ�m�&7ӑI�%.�S�������8m�vN뗨%�./�VT;!��b:�ӻ-fM;c��ȑʜ�ͼ�Ѡ�]�b���pyA��,�����g������ii��L����Δ�p$�?�t8A!���fyw�Lz�����y��Ȼ��H�P��� ��s�J��¿�)�@��ğQ2�MݘZ¶ފ,s`�=g�5��"�� c�*�:��*I���"\A�--,T	����c�L�f>���*9;������Ҹ�y��,N�̷2�� B����)�,N���~S���4�����ʳc�v޶��,t��� N�������U����mjz����ޮ9��[����$�����c���އ�;�4��9���&b��gHf����o���N/�p�Ҿ��i͹�.n�������ԫ<�v������F����&nT�bl�����'G�kQ�϶XW NT
������ެ�'b���\L
�TƄ��X�~�<X�qr���v�����Q�Ą���F<��& *��/S�AMJ���0&٤�k,�T%����cW	�8�&����QU��m�<�85@!�������.�.���D�&<A���~4��I:��˶z�oA�)��>wo�	�r����({SeI͓�>v|U�*�ýa�O��]37w`;���i�������?o� �+@;�îo\��#���*{�}�����f���L�^Gz���-��I7�Q���=p�
#{r�~U��4Ihr��\���^�~�u��Ʌ��w���u~~_�Q�s(���}��M^R��-6?j�\8��8Kƭ@���>:�UeG{:6譙��(.����2Oo�9Ø� �_�`��s�z+g噑�����e��&yQ�c��M����� ��XO%�z��t�ɭ1�E����}S1U��Akd"�������U~7�?��R� _s���n*z�Dא]����si��Z�eZ�y�@�����������e*�/zȉu@;�<��Jh����>u;�ཷ���Ӕ�A��x��rי O��E8�S�z�5��ϱ�K��[��5����p���X�b�}غ���{��5V0�ݎ��sF����u~_��r�eN�h���F��vW�#�d�Ŏ�_>��B��� -���޳.��k�0.&�(q�5��oQα�/����A1�����.Tğ[O��Ĭj|�F?֝����^�?�_��ۖ�<�-���ƫ�%�;k�P%�0�V��9e��"��T�L�8ƴ�4�S�yz�8���!��9oȷS��Ci$�6��{F{��n?�Dy6�A�I�5���"�3��!9m�s$.g����"���-O�1S_��1  �ɼ�+8��|��ѿ��@5�nX̛�NS���p�A�j�7�n��&U��K[�IN��z����[7S��Ÿ��f
wxj���&�W���ɵ����=���~W��B��L`qW�1�u^��̸g*���;���L���N��e����!�~�������e�\%㎼���nv�|�+�_��܁�2KVje~rܮ�-��k���c�O���i0ip�?-~��i  <��97�S�n�����1�tJMƴ0A����؛��6��%�0H��C}�#��f�0M�r�?�n�ؙ�sě}���J�c�����+��b;1� �{?����� g�VF(�<�Xި�&���%�-?�.J�	3 ĸ��vh���z슌X�W�y[�ϪR���U� g�]|����fA��	�.�z6�e[�l=Sa��<���e���3����W�'��$�ׯľRs�D]j�>k#2Zk�T����}�� ���\��3~w��[F��Go��)V��[d1�oo2d��ĈptXr��I�� �$���.�^��{���`z��ڸ*�ePբ_��l�~�x	r�7���h�������� f@&f��i��(>�ĸ�&`�b��ը��lT�cN���yx3��h�A*ǹ�_����I�ݖ����	1�{��01f����t�V%�p���n���\痋���h��[�F<�ty��M7�x-@J/ܼ�{hbUr���o<,����Z2��H2%t
�CeK�7Qw��]��~��&�q­���>C�L��R�|�Y?��{���b�돋���٘�5��>V^/�͑��i�G��M��]���ظ�:�����WoԺ�m@��	�e\^����Kz�܉oɞ��{{K����c�P�9���\���ȉ5�����lb0��GE:j`��?i5+�^��9��wd0)K
��~�&'q>�o��y��F� �_n~�!���M���ה�f���>p&Q狗��P��Mj|T|�?߯n�'�?I;�n��s�f,�ٕິ�Dj�~;?;7�C��*8u>�E��D�����=�B�:O� ��u	Y��H����OuO<NI����҄c�e@;��Ϭdߢ�D�'vrk|nڬo�v��O��^��$!l06FR5�����"#Mȁ�� c?b���	�;�#E��x�=(aa㑤Pqqi�����ȼ,M[^���$҄zU�Q7�Հو38��1�=�4�x��	q:W��ieD�a���εU�/�{����W��N+ߖj-?�ҁ�ؿ6�"�;V����U?��dWvt�
L�1�I�)B�����8r�_�ȬA����mzg]]]/9��O���_���]��Pa��V�ƨ_v�O��ɗE�2�7m��7R�0#�؊���F3 �?*�g�����Z���-��ˬ��l����9�����!9�ӛ�g.����Ο���;a^���G)�'D�@)L"��?��0�=�.1c��G�vԕʾ�� ��Ƈۖ�b|~��6=R5�}��K�;��43:�M�ۏd�����s7Y. @t�Q�y��u��goe+
;5M�X�$әZ�0���B��V�z��-����;fR�<\��3�Y�`ͭHT�����Sr\5�t��+�<�KԸ4�>��I2-��z�9\l�H�tz����Ѿ#�Z�j��[A���1��j}[Jc�LT���į9��w<�/B"6���[������Q��m�6u���X�d
��������4�ٟ�L	��)�l�6S���y�ޑ����zɑi�NR���罏�+�Z~D�.zE�R7j��n��I�~s��g�EcU��a��K Q\{31*�1��&�Ɂe|�{�	��Z���j���^��@4 ��d���1T��0kwD�1�\G�h�v�*�,����O`�t_��9�T�d�8�X�]w e+Nai��p;���wE6iw��O��h�:F��p*lU���"�}?��X^]�s�~`�M��߆c|����:�UMV�`n�.>�y�~3��dB=�'����<���� g�-Q��'J��u��{�ؐ?�Cg=����v';׍�B�j�H���(�i�E��[#8?E���O�Z��9�Fc�t��y�Pa6�1T�_z�׏�/=:t�8�|?Q�57L��P��y�pR�3LN���T�E��B��ş�]FO-g�6#~Tܨ��tF\�t;GuC��h��"$=�5��6��SSO%�"-��t���N/K��Q*Pk�V,E��=xaÖ9"��t�vΒ]�G�n�c�c��]��X+O���P�i��34r�j�}[�M�Vp��2-Zz
�w�*�h`V<݃6rT>�y%���7鈁i�g��r��lM8��������)�r���8j���-��7��V����j��m�V`�G0���W��@���*��=|��ތ�x���j&a�IM��PnW��wQ�CꖊC-�\~���'���~*��1Z�j���&L��1�vS�� �v�~q��)/����nm� ]ǌ��p��4bW���n�m�#�?��d�'WURkdm���TS�
?E3�h�] �D%h���ܽu������
Ʉ'�OϽ5�$-��ob��~�`���Ǉ�aL�J������=��?ˋs��������uwyr(��J��C�l�)h:�k<�Q���P>FbK�^���ƩI���A���-R�Z�n�x-�s̎
���]�	"j��t�2�� q��N/ �|�����#y��mi~���>�	\��UvG6?�˛����9 ��1��v[������C�,�5�L��W��'A����+���hn��}�G/ʮ~�>��'���q�1_�YR��Fk��   V��mD�1�!Ş)�Ũs+\�z�YY(����Oп�a�{'`�Q ��m�7s�#�����T��:�̣]w�$I��>�کv̈I���p��T||Z��h{S���@���R�$�3W26p<�>��[
�x����q�a�t���.æA�T������^Ml�����|b��&����jTOKe�r1��o�
�^�vŎ_��߆&�,��"�n����)�`�~�y�<��"������ڒ���!���ꬹ�4���#��W����Q=���+Mn��$�O0�o�]}e�]2.'� ?ggg�n}C�8��W���X�Y�!����W5�L",����!�� |�٣�KN�T��ѩ��6����؉��N��+��G ��v**G32��f��׮����8Ώ����i���&~�^��;��vE�7��ZI�t�3a۴��HP�!f�σc�ʐ{�У��F�M���������t�u��[1H9�!�O�& �4�`��}���?����I)��Bp7�Yʢ���#�ת��؉V�t�Y���G��w�e�%׈��u��[���
}��k*~�0jķ���Zw��V �b,;�7s@���磿2�-��)@�����⚪֤ޏy�M��$ªg~b����\|8�K^vC�� 3�w
)I% -SԹ\D�Ŕx�O� ���P��Rn(�������h�sg	w��\�V�F:�QT�HB;��NNHo�}�Z&�M��[ �d�p�����N1����%��o���VBe�g��R�C��<\�y���D�(�Y��}|�+ֆ�Yݷ>_.�m�'k��vՌ*�+�.��t�{�nZ�G���?3x'}�U[���L�E��5H�Drr�2�����@���X�zy��6�<��ל4S94�I��9�=����#`sPض����@��K��)�ئQ'��	�§�N��6>��[���`}ѱ����^�V�����6����Q@���o��7��y�rk�
y�r�9`���,�=� �c�{}�3BJmp��;MPvIy"�I���Z%�7���"�L�[��6�]=<ț��R\s3�@m�����$��Ag�}�]��>��Hd�}�6���� ٟ�<}&����.�xYJ�_{k�!��Ӌ��31�׹k�g	���o����E�D 5��[0G�Θ��l�S�h;�\�VeƈL�K�����N��yP���{�,=0�gK����, QE��(��[=�����]��0���7x%�,FTT\=�@>>��\.H�)�Cp}=%' �����h�ľ����"[]��G���Z�}�,M[!J0�&"�5�4-g
�/���z
�˞B��� �I��ɕ"$NŁ�ʃ����\fnz^�v�嫙�oΫv���}�٩(�s�P2^�ٿ2����{��ջ���o��|8{٩#z�ŋ��������I�^���X�d$�+�h�F^+g/4��^pF���j|�����X!
U�?��-	��LZ<yM(��*��e`������Ķ�)`�:+�'-�V���mMLL��=<<neU�4���]$�d:9}^{Sl�DPZy3� o��/�+�~�	p�:��4�Y�]Su��r�ys���I8Y�i�fQ��\�`)r��C-X�=U��;�7|O���M��$ ���>hfO��2��E� ��U�/-3sT���_����V:fw9���ٝ(���x"�"�1�'��n� R����~��I�[~=(������cff���1P^ڻi�8��7FY�^g�(�m�F��dĈ��D���K�߁�qTd:�s�&x����u"ؼ'�U�����ws�x�t�'����A��0RtG���Ɛ%�������J�6�[t��t��>�
��D�~���H���i�g��gg�u��F�������A.�ZT��ӿ���(��
�e�>)k���V�n4L�W�{�hk]a���NA�겆���uh����%F_�0��:,���4ޛ��o�,�r.6	Lqz�y�ީ� �!Y��sUOe�s25=������P��-M�+�\N�����������n��}��?p����iC�d1�����d�t�	����B@�|��m#uuu���?N�窿ƻ�qƋ@��z����&0|E=� �l�������X����ͷ7X3~�U�M~W�\����yn�4׆��LI�!Z=��e�9
*<��E�P�z{�yF�ز�(���/A� 21�	���&���N�c�0���K��eML(����������y�*�%�����dT����1�B(�� �5}�p�-�e�A�`[�c寅����at��C�kjk=�&���UU��L����b8�g���@r�K�o�{��몯�>D�YH�'<(�q�=����^~M������U��E�/�g�<�h���ݙ�ܴ[
�BS�\V���\��s�IO��}�����^��ع����k<�o&JѴ�����U���U������~�qO5��-�`¡�B�(Y�g"�e���x�X�\�iz��Tp�>+@1�`�3���Y��Ƴ��j�h�Q�s[G �oJB��z���n�����yA>u���?ƌ���t/�l|���9`��z�JPI�w�x�󍪢>�K��)����Ѿs5�/L^:�~g���ݞC,t���5o�(�.�h���$$��� �����Ì�"��yT0�ٽjF)ȰK;��D��T�!* 7�q��R@��KG9/^,KII9Iv�r�6�<c��#�f-y�Y�W]% qб1C�\c�:}zls�����gf�;t|��z���^^^�,�tȌ�����h��@}ȃ��>�wۉq�����7��)����=�Y_��h����F��׶����yz���ـ���ɀ��B�dOUT�[yRH���v�Q�Ea���N{9؟���#6��e����6|�2 �S�z��T3j+t���塟m��Pq6S;:@�ΣU�GS�Ffn�
��-<2�LR��'��T��w��詩��Q�Z۫J�	��(�����������*M$n��cjϽ�G_�gh����Q�5;����bO�C�y�#�t�臡�+���^Jy�(����$��������_\{�v�$�����U/hb7�}�|x���2�������'1?���f����uDJͰϗ���fUˤ7�&峣=+��N�R��!c�{���xē1ğ�5���i��ѧ�nC��z�mgŇy�����5�v��tI����Ww$��_����)���t��?��^�0�T�9��kc�ӄ�l��|���g̦�� l�قA�>�����x�}`�s���������AJj��ȳ�v��n)daxz`��4MwW�r����$�n�[&@r��a��7��
���� ���9��&d��B)�M��ɾ�8�ώ	C�ZS)cc\7ve�ןg��q��7�.vv������򷗖��k��e�!E�Ω߹�s�j����g��kHEhP�aX�k�-��&w��?
>:�	�<�m컷�wJ�Q�ݨ��ny��kך�LM����nn�@&$p5?�͛U��(��@
<B����vy���\�nπh��ji��lE Qi0�0Dy�4��V��D��ρ�ٞO��0� V�pQ�~��h�����X��? �����/eo1�w��!�6^+��k
ս+6��N�d)�aMr��M
�X�޹�h�2=C�i;��Z��p z��vI2H�{��uO�\��!S�|���0�옃߯��w��H���8*�h�|�6~�X\���GE��aT}�Cu-Pͅ��JV�a��f�6���kb|F��Hʬ�>�iG,	ڤX�'=��Y5�&8�Pzm[2l�;ܶ�NF���2�a\s��~z�y�B�|.TV־���P�X���P��XAS7��>�n �vNx~�a��ݠ��y�X'<�02�A���A�p0������ey�)Q�|E�W^���ATޡ���has��n�r�TŐD�X�1Ec���k�j6�Vq����SCL�\=Yt���h�y��y5C'��X��g
���-m?2]�������Ct�6�SGyB�	q����O޷H�a����%� �W�A� �/\(��bA�Vh�eʃ���I�z��ax1i.��k�kۍ�nh��'J9�O�]0�?�q�ٴ�+)sy����*��ƹ��w�j"��ȉ�����1Nx	��/�)�
���jVr;jɋ���%KȂk(cB֠]������G w�q�����$�m�ݜ�����Ъ��Y�S_�!��Ň�G�{��P�NŜffA+��@�L�`��8zr���,�3�����O�����w2	�I[d��3E��)�D� |A��|�٨T�א��kp�>P)�3
U3���dg�m12�d�o�z�dG��k���ő��㟉W�C=>�IX �����M`�ǆE�R�
������,T��f,�ؙ
&׬�cFH���̶&��G5

�j���/� ������z��ޝ�ü�)��vv�P���Ȏn��`�����ߐ��+t黱B���eI�e�D���<��=[5z..9�L�A,��G�[���$x�:;�a���M�`R�:b-[��Lt��W�u4b��L�:�\vz���o�=9A����N���F������="az2hr��k|'��)�?����+�N��*����<r�pM'���;�`�$ҩ̤��a�^T�����bD��|�og���#�����ȡ���N>3|��3Qƽ��'?�l^�*�8�4�� ����9�\�c�8��*ٖ7x���d�����#Jv�M�ȿ�6PD�@%��v�?R~�C���^"d��|����]"���iK�ML<��E����c��A5�����G��vݟ�/2��B���^6��� �,������r��x\1b�M���cVυ�ռ�WM�P<��Q+�m�n=��v�t�� ���~�����|ƍ�����eL���cq7�#UH���~U�m,�㫍��!���M��Y�0	�r�X��7��,�ch��~�;�Hy��A���M��a�B�xWb���ұ�/Q��u^�޳&�I��h��`zG�o�m�7Kx����N3�F�W�����
�$~.)�~�+k�9����c-
��o����ڳ��� �`���2��l��Ğ��=��w]ZYҕ� �$R�{ Tō��;d�����i�]QN���^�L �1���
guqt� ��vm>,}�>�5C���w���9<�]3ܹ��6	��^��z#����kb}4����5\"�\>)���_��04�Y��]ܜZ����
��������-�T�h{���&�c���� 	��)��r.��,Ɍ_`X���p�6}��g1!�p8+�h~q~�Pn��G�e�R$������o�]�؀�U���G�\�z(��� ����L�S��%�s.3����~|�?:Ϭ����/6F�����57�	^q<~���yk�ZM%L��UǉB�v�@y����~c*&��a%�r)l���n�*�UbS&r���;bXc��c''�ba��P�}�W|�߂��a�̀�]���Z�kw�i=�,Pf����?�����=s�\��/���NK�@,yPa��^�I�3��5���r;C�Uכ����bX�Se���R�mv�j�ߛ�[��řSk������Ģ�R{�z��b�dO�]E����5�v>��:M�}.�qP{����0��Ă��Ǥ�% J����� <"
��}U?Y�\�b58��q���Q�C(U��3o�~wW�����慑=���~
��n��_-U�O�H�7sC�E��~șM�qD���	
eF2.��y�p�Jr��/�)���/�+�>�d�A�?QI�
%w��Xy)�:�o$���A��8�s�����6���v�ޞ�u9�:[:�n��̸��c��%
҇��3�M�F�~��8�����	�/R������k��H�bVxr�[[?�@7ϰ�zn,%��{��j�ڈ��j�"/�Tv�o�%����e~BSAu�n<|0V,&�RPd�d�K�=q�����l�l�ئ�|��
�LLh�>~N͞�2��cv�o`̶֙�JCo]��~������Gp����
� �+~�q�Ο�^��V��n�x<~��I��b�<�#;���5�6))�h㞼�aV�C̾X����f����C�ׯ_M!�/�K����y��pԐ�S0�?�Q	���/A@��J�	BN���{:�<5����*����+�K򍿹x�pag����o[5�
r|���rS��>/�q�������@�H���c�q<Z����'���ǯ���yo���R]E��>�<�\�p�6?z[���T��!%Ssk����5m������	�5I�zhn���Urr���9����J)u��a�z���iG��D>i��,����s�ߺI��`�x��/K�))��;��ID����D����m��|�4Y��={?��?r=洸�(�Z�!�V�аp���Z���i���nw�`�p�����O��(d�g�"jd5�;�_�84�08�a{ol�
%e�8��Uw�Ƥ�Y��;���7�6�m���O���͍LG-l%;Kuk}T�+��
��Ɨ:�.��N9����]�ƀJ���������D��-�:S�=��FF��K�w��`(b�^��Z�;��;2��fB�#��:D�i��p��nU]Zz��S 
���bbb�MU� �S�\ۛ��B�J��lXnk��^ y��,9&j���9 ���@U4H���u�|�p�<Wʣ���AW��=h+_-�bov�P���c!���7��������z�ˎ�L�ۘ5�^	j	�/�����k��c�f.��N�O8R��kΥt�I�֨ۑ�g�A��M?Ɲ.i�I�?�ň�A�a�.���t^�����%��t�az���B-h	�C����_U�Tu*)cv�v�Zḋ'�~wNu�ݖ���*�dk�-�7g��Ԡ� ��h�ۀ[⇗�R�r�5�(y�c�lk�������K�]vo$����n(�S�&qRSe꩝��:�ȡm�<G�2Lk�w�_���WUTTƟd�*�FM/���6���'7 ��G�\`7*���Qg��҂b��V�a�4�p� �=۱�J��QW��-�-�s�9����T=�Z�ݵ읝���M��*-��p����A��Uz[���Aנ��4$n���:�,呋Yٍ�Թf�oO��QČN��Ի��(|#8g�ylUVh����ƚV�T�!}t����n��]��Op�����gee��%������!����~��>���n-����%��0�������	�<�X1�z|	9��}���Cq	����lq�k�M��9���#ʮ�įCH"���.�>u�����`��EV���SH���p����m���2���&�ƫ��L�e�c)��]��+Q��2k�}����������.I�L������^�~FXXG7�,����k͈��p��h��i����l;��s���\���B^�&~�?�"����?|�"���+W�"b�¨���s
�j72d� .���g�F�/x�W�+�#d�٣����Q���ю�9���iJ��\8�o��	}�fjH�>��A6���J}p#p�>�y<z�5Z �if����a��DI���x��ʘ\�f�t��3ߥ������B���3�O�3����W|(���^ipG�t�T�|y,eK��=�PE�^h�]/$�&F2��@����s$�Ӄ-�\�/�W�-*�=$g,�f��
-Ɗ��P����D��T�sDZ�ax�C�L'�7����ʞ^y'�}`�돑�.�}�j��i?��
�8'����D��a��'k�|��tGVvy�E ם�ƶY �`L����I(�ь�P���Q �v�_�&�-�j&��רapb[���~��D~���}V��N�@w�0�z�8��Uhm�o@QW�l�Hm��q���?�F��#��'Qp��Z<(�p���z��^	We�w�.B�~��9�V�8�T�w_v�Xﻹ􌈕5�.���6g���~�P
��sK��F�-�>��ρ��~��t��֏/H��� o�Cw䴦�T{f}�@.3�m������h��Ғ^E��DV�o-cbJ�k<ږg@�x���`ƍ�}i���˪խ�6jЁ}�(��\a/,��p��鷛�����z�\g�z�y�o�Ӈ��~ !B��g���r$�qyˠ��M�@���xf I�����39���͍�/����	�R�@�� ������s�Bb%
�T��An�OV��u��J �Mx�|j,����AE�aU�,wuv��M0����5��6��A�]�8�h����Q�W��ey�f`�m1��GA(�o�=���N�(ڪ����i�< ����s�z�ss��1��x	���������5� �_���vc	�'cd"�E䋿�1���>$9k�H��U�����R|�*5hi��Z,���p���ަq"(�f����p)���i�����X3���a}�j�D��R�ӆ�Ө�\��Ɨn2�!6�2Z�/2�rh+����<֍�bs�
��5�}8���ӍB���9�����ڱ&�B;D��}
K~2{����i�y������hZW��1cT:t ���2�*�s]���g������O���'PJ��"*�k�v++������0�P#MMM}2�����x�L$�{�s�����5$J�q�%&LZ�08��yb��8-qw(����16��/�W��(���a_2y�'�RҌ����0���Ws6�r���5���ncz�O#+�KH1g�+z��H(���W"�7{ngJ���?(y�- 6�t0u7@��F^��{���P���o�Alw3Z�T�~��n���C�*	�4��4 ���[��u���j��=E�m�9e�T�aT>k��z��7�}�(9T(���&^v���z	��׭�~oz5!9�����*CG����>rV��1>0/�ի�E���D�P8"g����_��1�:}���ݻYOD9nף�!%В�-|�(h&�ٯ}�E�3퉭����������˷�����չa �{a�B�+L ���V����H<�o1@N�&6;%J��U�̃�����t�?�/���'ZKJ����7��M�8��s)���
3�Eu��f���Ń�2�	����8��@��)I"\����ڝ�s՘+k�ZC��Uƣx-���{7��D�-�H6F� ��]9�n/���ވP��ZbFI�����$�~�I�=Jx%8��S�>-�CLn�D�nd�^���Q;�L�X�v�W�5�3��w�oy���)��H4 �i�~�6�a>�
:Iz�AXv�.�qw`W�G/�)QW-X} Q6���oEC�����n�iff���J�~���|k��\8y���Y��L2�z���wD��V��D��/�> 2���y��tXW�q[g��i��E�bJ������P,��[Rmʴ��A�a#�i�CQQ��rI/x���p����ST��}1 𧨧��Cܗ��.����{���ԏ�}}��>��a�?!P���{;4����p�F]L���w%w-h���{��`?"##p��ǟ�$�6�d�d-�$�ppH�\���yH����X�~-L�|�94��DsOO�:T޲	$@Rԋ��믨K��=�#� �L��S7I�_E�5����#)�������1���%6����
iy�B��Aȹ!)+{i�QSi�{-� �[)g���x~5y����H2�M�=�%F�F�.�ǜH����P3+�_���EH�$�-�鲩�B���f�P��HG�xwk?>74v(�RgA�q��C�@s��\��%_�ӿ��\o8b����������#��HEi�c.��;W��R�;wg�w���<��(���-.a����+Z�X'�ď�w������Q�e`>o��VG���@�d�o�7�2��к�?)ciFQM~J��yQ�� _�=ӌ�H�4�%��N�u����V�J(�3洷yth��p�;�s�-��FY��{��}��)�W�E:���\�]���jx*[�� N�����u��ԟ�@�n&��}ȝ޹������&yH��z�Z�����)�M���e}��|���q�e	1�X�+��Mb��^�<�8_%
��K�����
�uL�7l�p$�� <RrG�䫆�nUS�Mm���6�!c�c�mk�o% ;�y���O��-	�o�:e)�������7�����(�Lh�/����'}�0�h#�̇��*.%�-_b��-1,>���[L|ì��>e����Iס�E�F�[�3z�+㮹څ�v���p5RR7M yN�c+��H逅X\%��c/	��h7�a��wU]�#��F0��^LެA�����t�|�/�տ����ᄌ2�šf��Sм[K�h��r�dA����^1@�J�F �4tˈ8�ძ)�n����v�"��tr�4\�6i����B��K���œj`��g����v�!�ߴu�E��j8���l���C��K�=�PU�����c@	��3���+C^+!�<�}��ٜ�D���%�7�ON�hLكg�T*�;�MOMI�%!+���?.��Q��J ���R�Bw�(Y�Ĺ?�-�r�<��k�#��o��f�ع0cȾ �S�K��³�y����6�̑P��5���z���KX�	�zH����;�+&��,�_\z��.�R~�l���,�_yH�|�����4Ld�	�X�J� �jM�����X2�dx���`7=r�<p{k��;b�&�H�G�G.�/�\���k����ƛ�$IӴ<s��Tyc-=��/\��~��g�ʌl��K�Ӧ����(�5oB�^cL5�r���ǀ����+����Yz&�����#��|��a��@��?fuYE[���J��ؑ�ګ�L�5K[{ob��EK�BlboB"�����|�����"ו����\�q��.�Z-�W���LQ�[�,��>~r^̣����Xw�Dj�g�\�6B�����
9`֚D���K���ۡh?{���gx���r��,͋[��|q�z���"��s�2L�?�}�n],>��)�>�&鱐��7�z�a��r����"�uRꗠ6�����
�4G!p�5{�CD�m���,��ӵ�:��(>�X������GZ?	�iP�C-Q���犆^5�O�i�'�ɽ�PmS`�?�&�h�ٷ�ӱ�cx���F5!9-Ox�[#�ޓ�2�k��i��9 ���\���f�^i�F��0=.�~�l? ab�k$ �'3`��S텼�2����.�c���g��W8�}N�.�"1&I��h0LU%?�VK�^Ɯv�h��<�Y�2��]ﰣ&(��E	6��i�4<�G6���z|���0�b��B�f�6n3��`��|��KU8ը�	c���H�gF�^��1.���5|�%a�����E�N��=K}�a��VD}���Z�)D^ P51X]n�P4i������AȄx@�=�eqi��k4®f�"�P�C)��ΏE��$�%
L�U�}�z�Af����{��:��amQ"�=�VS�Ov��{\ױH2
��R�0�K$hM�	L���.P���{��p���C�ɘ��f%޻�c�{cC����C7�)7���C��<������;_�X���b&Kۏ���MSҠ��F&
�捥B����rk�|mt��^��>��x�?O�0x~�=��!�_j8�*X�f(#mA�����c��=.q��Yv+_f�e�����=��Z˾�u6_�&���3 ��M]'��N@�K��.E�[	�&�$Eu�2�2���R�J-7l�7��a��r̅3��\���N�y��w�y��o5�hn�S\�<�$����Ѽ�s�/�I�]T4�����|HM�ݤ��R._�2\\-�<䛐_�/䗃�{#��v��E}�j��ߐ�|��.�C��f9Jq}&LF��C�; #@���<۟������uO�}Yc�µ��rH��w�����To�o�@�(�`�#�lΕx��a����d{w�M?k�4�>Z벪�����0��rXn�?��Ee<*�k�u&臅䓫�T����7�Z������k���O�����Qɱ�n#*9[)V���3A$�]g�/���Yc�����G�3QA�G�#@F#���=�N8%_��1�k�/٪6���#��IH�y��'B�X&`h��K���m�m6!����5�O��|�w� it$��|��o�����A���:ﳗ��.�s`]��̷���hE�\;b��P=��1(z˞���-FO6�?�"�{c��������D*���.]646fL�-�x�M�ˇ;v��~��uz�ZA���8
��6��cE�kD�p
vV�q��H�$�!�'z�R�?6jRω)�,��1K�z�1�z��}�7��lֆ8�A��N&|*�m(w��X"ͣ�/Tlؕ5)��u����I�ƨ`ǵ!lȤk�Ž`�c�vU���o'�q���j�8V[��4�|�5)�zۣR E�ċe�~]�7�8NcB�iw_^��l��p�֧��Y�żv�pB�vuN('4�����90�H��]8l�;�
A#�o�{��A��4�js~��nq���K�"������Q�J2��}�!.GTF~7 �L�P槻Y��go?",q�`k3L�g7b��� �D�q_�x�V%:�oD�6��:�B3 kI����Q �K��B_Rڦl�;V�O�ةB����=�h_.�3�=$������n���Y/�ދ�,sW��E�3�6(��RP�ʟ��Q;�@��$���K|���X(C�����7v�|����C o�m��S���[�zWl�����CUEn�l�i�F�_�'wk��;�)~jjE���]��}UpU��vN�>�w�����H����(Xn5f^�[ԩC�-�z���h�:ܡnU��8/��{b�vs��T�ҭ�9(HJ����$xGѡ`�@1��<��-�&O�B�F��������q�����y�(+�vK��+D��J��U<Y��DBN?�&v��55���/F���!c���� ��Ec�M�iDS����<Qrh�Z��a������GO]W�~]�S��m|���,�^P�o�U�G�g�Ʌ���<?�������5��n� f)�7Q��1C<Q�f�0��t��-�^�6�ނ'k6GSfk��gz-o�5[D��U̲b|Ф4r)�3���{�R	�/��ܸ��w��r�B`��;=�p(�6�	�ޣcTLY�ku�2Z�_�<��=��h�׵~���ha��de�5d�B\\1��GI`vεeQ�󏩨o��x��!poI��1@��]b��^3��8a��4x��Z�����L-�ue����EU�������6i*rtndq���q�`w{?���̇l#�>��bAQ�7r|�vԟ�����8t�����i *���up�W�^�w/~�hp;�s�����E��D�<�Wl�w�����;\>��i�.qE�Ĝz�K���)����O&�Ӥ�:�|-2���e[�ޠ9�2�1�g�����"a�ޠ�2u%�Ύ�!�r���sj��0��^^��@<�R���|Z�y
��������\��s��R:�|��Ռj�Cd��l��d\,%j�u�x
_�$=�s[�Y�g�2W%���M�"���]zl��Ps35«*s/Y-��j'bTYF;�����:��7����j��@��K�:��A#y�;��B[B�W�;7'�5L>`��Am[�q�7�'�w���f�7��gAF��jw0�0S���E����P���4Za5|�g��2��Xw��o��� V�����-w.M����8?���g�b���}b��O1�Ǐ�N��K���K���}��~�s5ϫ)��UI�Q]���u ��1����n��[�6�.ܚ\~�j�Z�8�*r�<��g� B�>��A�.7�!>KÏN�$
��G������}��H-DV�G�J�4=�S�nY{�>���ﳧ����'M�a􆰷�^C�d_��%�W ��\�b�O���Xl�d�ޘ{���. ���d�c�Q#)^a�ibd�������7ɽi?Ԧ�C�@����9�@�h�x�O�s��J\��K_�ƍa�C���/zi���z����c�ө����WVW+>|���ie����mG����-
)ge�vH��H�2&&d��5�S���*#�ER���1T�e���h���+�Q�� #	甝WE�=���G&<����_u�I�{�t0Oo����!#�6ZcD����վ�����Q�^1��E}�W�1����:U�e
h�c�º�Ӎ��ueu���wZ᭦�S����$���3O��Y-��T9S?�[îak� ێV��Dv��e6Wʭ��;����k�˒B�3��6����$.wݽ#Qu��S4���$75��r�{����U�:_+&E��(����f~̸ۀ�ww���Z�΢�VW�����n��;����yyN�ڷ������`5%Y��W&���%�fj{�eA�O�ʇؚXtZ�-�Y4�d�WkV��8x���Z�Jm�mS����y���@U�٠�Kw�O���/qEJ�a4Z@�hs�l��h �<�yJ����K"��Bw�)��I�֖�f�ۊ��z���Q��$&��-��L�r�S{j���ZR��X9q��n"&�qGKP�������#���r<�H���,�j$��ׅ(j��.�U�8k�E MN$H���߅`n��ma�-ʼ熔F�3k.��wx���\de�)ڝ�ȎXf���/�L��$sz��S�pV�k�¬�qc���N�:b�l�����<���ݘ?�(h�u��s�`��������{FWI� ����+c��zHL���XG��F��<C�R�ȵ3h[Iϋ�_,l<e�4�_�9������-Q:���a||��K$5	��ۂ8u�z�B��xX����鷽�Mt�6���]�=�P�ﳞ��V���`���\��5�}QD��P�����IĞ��f�/���jM���q�i�k�F�����F����G�~�	F`wR�Uy��`�ȔLNZ���'�(�mi���7���y��G�p�����܋Q5¹�!����7�����*�pܿG���8�|8�(#pS*�[�l&��*^"�_� uBh>�R��o�\�w�7�j��+ĝ�Z� �t�g6z&��$�n�q�S�/B�������/�����!=��H��n'+~[g��"LY=���x�D�7��d#܈3l ]j1��R�4jM@0�k��ʍ���d+c(��ﭼ?="����O�:E?T�:���[9�Uv3�;AbE5�����_=R��C��]ЁUש��?K��^T* �WI*�S������__M���5<Yf�N�ŗ	잗4E3՚j���?�{��G�N�q�Τ%��Ɲ��:[	��wo]E�~tQ�������U�/������7�`#1'譜��t����X�՝��8$\d�G[�RK��y��~A��Ҩ�	�M,�4~ �ڰ1��tm,+8d���M�>#.��J��}<���b8���϶��cZ���d�J��jj�c��{�}�1U��A�*�ΝrI������`�n�����i�]Q���p�7���(�Rr���<� O��z<kj���og�?s��`�]_q�V�qqIH̎�5�����J�Nw�h�y�����t
���e�Ct�K���m�����cq)Ѭ��:Y��4���:>��@Vs�#�$�� ��@��obn�ܰ�7<Z�-�b	�au.y��9�`~��NȨ7��I��(��4�k+���r�wP?�����Mz�>����9T�yW����͌��3|�ڨ�b���������C�f�j���s�O�An��(na�P31���6?�M>8�ǵ��������hC��N�`&��t�d�`����|���&A�C*���5�7�k1�<�g<���65�������7�k��[�M����K���ui�ƻ�o��:'xh ҉����H\��絺���2�Q�*�8�U3E��A'�v��ߡ�6��6B�-I���)��9��8�X��q8�������t�;k����l|��7�ohn|y��������R�
�5!OTnm�<E7�c��:�E	�㯜µ��5^�b�U"��7 T�Z(F&�x�Ȋi��ebI>8
�/y���vA��*�	�O��¶�K��0��,�
Ė��M738�6  �`�=�b�[�����9/N� a��Rg^lA?Xt3/sʪ�c��ݿ�e"q5FF?����6:�'3'����:��z-�vf��t�q3��g\ e�w$5�k�8ڮ'��q뱇����Z+��i&l�8���O�$f���|���zl++ѽh~p8��� ���>YΔ����VW���9l�O��4/��
�}NLӤ�Ηn��#s��|d��ƍT��3/�� ���G�X%{�C&��lc�~��y����C]�py|�۴G�6�.ɒ�V+{n���NA�E�
� �`���|�^~8{Z�R��������0��3��R
�A�6���pW-E�'��\�b�~0Ԇ�8�n���Z>Z}4^��p5t����$�q��
�M����U0��J-�aJU�i�9�U��`����p�
�I�������}�v#p[�=z,��iק8����oB�����z߀?�B���ʟ&l���A<.�!�0��w*2t�(=��fj08��y�n4�EAe������$�O��捼�򝨉vb�4���*f�8��!J^��p#��)��'����" x���pe�Ğ��6��O���7�<(��rRTB{��;�a�Ǎw��$�~�X��oa��O냠��O�y���&���ĺ+���ib�E����,y뒧P�����f�e�j;�K5�Z鬴�d���deօg���{�^�Y�T�%�ѻ&����x�*���u�}��n��oSG�
�^'��=&Zs;�Oc8Ӹ�C��F� ��G(�{��f8�7��kxs@h1��wk�i@�5��d{��d�.;���GPص�W��6�� ��4�����R���G�[����ݕk�q�YT-ѥT��F�Y�$���5��ëF��r�i^�s9nsm�T?J�5�1��g�2I3�O�9⪾-A�H\��?��?�	�ؑ&BVO ������L����%�6QSRU����t��zR�:�K}�l�����=0�lnhӠ⋖�:�=/�ȶ�������ˆ[�t��Z/��d��/B?�o�	�̐�@�`�q��*U�BȄ�a���>au�3��d|�-��,�h��(P2�P��(�E��$�KUР��X˪lS��B���װ�H�]['дZ�Y���\0^+�bF��(H�A�7�&Z�Gc�}�t�yɐ�6مi�I�����+�������-?�N�괈�
�Jt�c|-��/p�z��Q.0k�B� ��~i�o8z�6��K�f�#���ۑ�R3-?��5��'/�u��y�V�Ք�<riYu'�ܼ�z%n�o�]�%��Q��%h��~��M��,ۻ�l�v�,z�
�Ū�_x�f�7P*�t��\�#��HA �k�K�����&���		ǳ���f�+I�n�ߟ ��%���dm-���v�����ï*1V�i���`�f��������h��@�޺0 �ٴ�W"�B��,��F���Ij�m���*UH�,6���>n���cAe�魼��B������9_֤T��lI�8� �H����ST�=�n�}��X`*xgQG���̷7i j��O�#]�}-�h�B�HEn��+�?7&����0�3���$�"�;d�O:H�&�|���3J��5K<����qԟ�:� g�/�2Wc�S�sX��NC�=��"�vG!�'��d�"�Gk�}�����XÔN�qe�}NiQ�Q�!+�ѳfH`'_^g$7vh@L0:,cd��^o��_:&���d}�&�S��� =��M�K&�ڠ|�Î��iq�,Ү'G�6�ؼ���7��E�X���H�m��fS���z$}}x�����jZK>z�F\\<Z���:yL������Ja ��i<1<8ɣ��h���-�u5Ё�Dn�	�6�IIr��^!�\!�˟�}���&�5��h��W��\�x��ˤ��A��=i��-��������oed�%�@gZ���*��_���+h����k�+]�y�=��`�ˡ�v�-���P/(֫=�)���o��.�'h��o��<��,a���-�o������#�_��\�ypO�	d
��/N�3P�0Ɣ�]������l>cx�q��2�����r���a��>9�R� �RHh���f�` .<�p����Ǹz��Q(�I�h����QAM��,�\>zN�b�@�v�-wY8 pܒ/XR,;��lx��3,��
~�>���ĥ�f�k��\9\��^���7�n�12ɇܸ����?�vY*��yMy�M=:9�\tc ?�1�d�����>�푝X�fsZiJ�
����ԝ�U���:;�a�嫡�.�09�)�m%�(�tx��?�d���C�CQ�RX\���x[�������\;�f��$��{�Z{�SP�ݸʆ ��|x�\�'�3m7vsT�FTxhJ�-n�%~�a/�\9�_i���if�[�_N��˟�� �W˛���@�}Χ���;����=�pcֆqy�C�1�}�$�aZ��<GC���7Y�ymF:��,x&�$��fj k���%��;�����n�1�b,�`�3*�QE�F^� S��z�H$"�����2>����g���b-����l�"p,z���>֦���:��;:u�Y��r�:��Gvz��#��П�]^Eo��Y��A�O���h��1%�����O�2�)Y�F"���,/@ bm�`����؄�;()�GM<�k۾�Y^6���h�eE6��qV������Ҍ/x��q�@�WGf$���U�h���~�s�4�	`w�����G�`�����p6�&��b�c1`V�h���ϱ[ҙO�^&�9��V�	��ܹ�:p�߬�IÅI��3�hDa�k��BQ"��Z�-o�`W���ԨW���:�?&mTr@Q�okF���w��
l4@fC�g�l�����6��e�i_��0O͸#�d��R�>A12f�q��Ք��R�D�8����䩣�D�J����V���
�CclT@]q!���F{�lđ	��n���֌ri �<�9t�V�B��j_P�nX�� ��ѵY��r��$l\�:�7�=��������+I0��+wl���ۦ��{��j��ҭ�!�0��)r�KvY� _�
�ѽp�ts`� <�]i�v׵������ҫdd�Yn�k��Am��S�2�/���ٯ��߅FysW4��}G�~��3��HŜ�pZ�����vu�/QP�
��@�����:Fi�h>��� ���=�5P�`>u����Y���ft��<zR#�O�2�8tL��y(J��y`����|hO t�6ٜ�V�ٱ�=a��"K@)Q�x���v>S)�^��3Sek"�8��5���R����\�B��{Ò��Pd����7�'���yyۓ�z�[;�Y|~�]�|��8���1��!�
�Ҩ3��MV��lw�^�3��sh[�y����`�'�l�5���؆��#X��-��2;恱��n��RyS�G��ּ�iȸ��u�l��R8���53��v^�Ϟ]y�(��(F����S����]39�Q��t��:Ąmm��� '�<�[�������<���U��v��H�ʼ�����Ν(���|ԭG3��zq55�q$޺Τ�Vg�w���2%�[�@[��Y�h%��uL���^�5k��Z�M��E�懽5K���C����$�b�g��ؾ��M������۱��zM��m���=�/��i|�v��DaJ:%�w�ꨉ�ZM˗�k0���}nޘ�"9���q��h7�1�U;#���|�&.�̘��k��.F�pV/��y�lȽQ���K�Wx�Y��x�櫉o���TY��x�{8M$�ϑ/[%G�u ����n6�d�5�����H�˟�9G�bv)v��]��:֒j��u�2��(�g�{����σ�Y���&�x�1���a��Т4��J�]Mh]>�zgW���hi~�CTh;3L��, '��p�qղ"��*90�SW�jd�Rb��;�#�/322x외]��Q�����Q�ҷq������Խ��ĉ�[<�=��L��U�T�R)�V
L��2~�)���B�و�\�44�(le�@6n��o;�Ub��ew�$��"b�Qjl1�C� �^2CS���L�p��	������X��&� ���r��?Ҽ{�c�`D�]�q�>=�r`����>9�)$������!��*�1BH]1|Ȕi�t��E[�>�.�	"�����-R�9'�	�)���0�]>� uI�9E��՘G;�:��LsFO��2J��Z>\мs� 4��,#""&d�0x������7����@vR!��@�7� g�y��bͩ�Y`�&�yxmNYU\�x.ǩ�U�������~;��Vԭ��T����>;ł�\Cc�8�PF�u�x�M���*AW�9��B|S}���z�+Z���.���r�f�wu��]�~��f�)�b��T�b=��F^d���=�{���U�`ү���	A�1D|@�*p���E��S�{�ָ���o�5������'�^�5Q���n��wXf޹�xa����Ӝ(P㻒+��xp�d@#�V�x��{;�-'oȓ�O~�sY�тء=�s�ۻ����+X:�HqZ��e�:��}_���F��k�dB��8�B�����6�9�#�A���Et�8A��0r��ʨǦ�dOHe��l��� ~j���s��K4j��G=	�\���;����SmkϏ,������n��\v�,b�����I'��J�>;��>�����՝�D¬m��۝��#�ή����qq� ��3Oy�����v;][d͹�ڢ?����wü��r���' h�վ���88�q���H/�f{��z�Q�0��ލ�*g�����/�b	�����r�\���}��^�ԧ�Z�W����ϊ~ҥ?���v��q���誔��G�.KL�@�b��>��n�x����gHct��L��a��1q�kV��J�j��޾~Z���_&fx9� �X;�\7X��z�V{�����tGN�$hY�>Ց^�����(}x��cM��N���rn�ݬ�,��=/zV4 (�<y��?����k�e��b�[�k�3�c�AW){�<�dZ�z=�n^��9�ɺ�%��4oo�l������k����3
4������'��*�C��\�?Ӗ�j��r�_����zw��3;�Al��r�=<$-��Po1�ėӒ5�g�w�� e����:��E)��&���
H����u�D�#�`��W�U�НS9SK�k�����P�C!��"w2�ފK�Zv���R
��z��_fv̾F�o(#i���]�1��xh�m��`����A^18]��W��`ژk�{���7�4��(��t��̴{��璟������%��gUA�_E�����?��8/i�sP����~��!5�"�L>�������REZd"�&����PEin��ߤ|�0Wld �>Fɪ�:��p�U1�kͧ��<�潏P}���&��~�$qе�~�U�� ��/t�_����޳�#n��k�5�N����F�\��\�#l�l�_���F����(/s��$��>|��$n��ݝ6���+.�_[�L��&��`5>shT�
(T�}b�\>����q"[� ��2�_$!&ƈu��WS��H��_NF���/�+QmlC�]3��U��h���7�R��w��ws���
T�SW�tJ��!6���Z�9G����1&��r��ŋ�i$���+��3A���ެ;1���]�Cm�<�3*�(pX���b�yq^D�:/�����-U��l�Z����ej�Kc��n�|��F˧ȇ��ؓ�B_�lNk�3�Dūb��u����C�@�1W���;��o�3�Ѯ�4�V7"_SDY���!�J��Cm�����b������S�V�������q'��g�nU�I�2A�d _�a���뎽�.��M���%Q�g��p����?#&������¿�����]���X�^a����b'I�$'s'�oSP��(���B�"2��*:�|ݶ*Ǟw��ܼ�Y�3���Ԇ?�0ӌu���i�	)k�I�}r���z�h��Z�ZsZ��F�s�r_x���v�%���S����1w| w�޹>�Z�r��}� Co$�j6@��;h)�����r�`�Z��$$h: BسO�.�R��R�!(�=GK��Vq�'����q�\�b�꛼���7�T����_���V44z�Ѩ���V����(�{V�O�mcQ�LѶ����	]����~�'�8���_{>_��J[��6���Mjy���GGs��o�&+��?���-}I����;�
ʟaǰ9�ձ�����KT'�#�=d�ڏ�TD��ƤVx!�?���&��9Tu����;B��ɸA��䢟$^���O����dr���/P�q��UI�2Ϲڛ���h�%F�}4��MU�X"8b`v� >j����d����|�B����xM�2:��n�Ql �>eӎ|P4�����Ǧ�/wY_*g�c�]4)����؛w%Ը4@�߻�iߍ'P"	�o��R�/�2�Dc�r{_q�1^��g�M=�^+���P,{�ra�V���	g��b��`�C�K6NA�0P�nk���J�~�$���u_jL��o�Öp���zk�;N��}��.�e�������ܸ`hd@ؙ�üjs��ro|53����xGHl�0�*���5Q�<���+4���F������ep^��x4�ݽ�MM�Ɍ����+��p)���8��if��*d�[_Y�P\1��d��D=��$W�Z�[G���[�Ř���U
ͫW�j�V.����2���C2v{�z;6��s7�-&P2�贿xS6�TbV<oӲ8}5���&���Χ[&ϛ7K����,�y��J���o�R�z\_OF�����sbw�P)�ٔ��N������+�_��/w���5c����5�)�� ��F鞙�ʝ������2}lD��ÐS����P߷[��Äw�?d(~Ƹ��y~X���ce���PKi�`}��
E�>��"D���Q��.��n�)�2e�;�E���)Lj�����2�� �	)���q|�·�W}>�������y�'g,�[q2���v�@�n�`�!?���+ȎOU�w[�����U�#�vqyLP놓����8f�f+���I�ur��J ��5�`���
0&fb��r�`#wE{2�Cy���cń��?�j]HzN˭����������J�.���@��z�z���a���l �XQS	�y�25]o�l}��î�8�L�@����0�'��mT�g���(gv�o�!I�-7��b��CI|���\�s������h���{GOϑ��ǕIPߊ��4�'���8��d�l���:�X ��i׌ǋn��K��h�!��Ρ�r��'��r8��J)�#ȶ���(�6֤����s��Ub��nQ�������ޚ_Š��NJ���8H���/c�ХP�ye�[�Ӏ��J���}�Шֹ�;��˸ⅉǺZ���rOl��� E8IuY���e�zΏ�B���bi��[���y_��]u���}�{��m�=�d,��;�vz��C��o��;O*a*_����f��7��[vdؽ#k3�{�M�S�\:H�Fw�E2(��j�Q�B>��ɓr�^�?z�ܩ=&�]�Iٔ��~������5�r�Dh�F�zĪ�F2��{�!6��F�����	�^��_*��}k��9��Nu��T\O�prl؋�s��~�0������ُT�%��KorS�֜֠���
��D�ӬvUU챷�kC�I�A7��T����k	�,�$��@�4��Ж1=0�P^��3��@����e����(d����-f�śdd�w�Cb�����ߑ�K��v�O�I�I��c��Å<c�\�=�(0�'o��0�8�m>�)Rcv�����K\�������su
����n�@��!�::�f�IT��c�Q�g)K�z�xO��*"<��p�ݹޛ�����l���\�ZF_8�������T
L�[MR�ZJr��;����H�̦�e��"��a�݊�ؐ�!j�2��a/�_ ���K��N������'$�֚'�ڪ��IՕW���L5���/��v�sƁ��~�{T?��|Ϳ�X�Ʊ��#���s���;BמF�w�9V�D�U��N�̕���=�Ew+���B��˨ڥܤ�.��U�4�(4nkk�b�6�+���N��`V�
�$=Q��j�?�!�q3t��������&U W��y��.�+P)�/�F�ҋ����+>��X1�	/����jT�KF�	���#�{���ħ�z�������Wٓ�]�T�������oI~���ȥ2i\�h=�]���f��[�7Ͻ��{o���@�Z���u�m�[CC�=���f����`h�hϳY�Ց+P�+��?I����Ű2�h1pXT,+��Pl9�v�!�c�'���Pֈ��c��Q��מ�qw�S��aj�/ˡ�w��8Wm��<x$�������ÔI'�^�~�Ξ��יq���χ;�:��&��J�zo���|�(�O�V�~�}m�M�����ʅ+~D��L��;<�!�Gu��l�]f�z���z{�L�6�[��O��R�t!"YYY�K���>����h{D��"�R)�\^s7߹��u�9��m2h��M#Ѕm��;C���^�z�����*u����E��m���4��_l�i�8U�6ӵ�Uˉk������D[#$'��莛&�iL��`(��O�ew�n��W �^y�4�sUd�;�o�|z��ʽ�"J�Ƀ|��X8��W�;�5&iW�jkݭ�9����=�:�Bj�_q�����l��1�F�."�B�IMz�s_T�YЛTU�[oD^1����V��4���X&=�i.ϩp�������3��5���m)��ʮ�?�2xf��'� ��[C�R]����՞��"#Dn�=~M�ٞI2n�({-�ó3k?�,�W��a�AC�R:�\�nٸ�}�[D���2x��oEVښ ՝S���r%�< 6�LǾt �-��rM��-1YB����;E�|��;��&�w4դE�/��5�YD�}g��鵐��z&E�r�}���1����K��д}��#��}y/6�����F"lx��(���yMt��׃�[�9�fƦ6��L�t'�tO���J�6�T�� ���-�Z���pڟ�S�'/9��c���9R���0�:2�����w"����#��-[t%݈7��)dP��#�L�<�"}��W^�K��N����wīX0i~ۼ~� �mt ��jGu���Y7��%���f?Rq[]������i�q�=���=�ĹS��KV54br���,�-�W�?�L�Z�~Gw�\��F�����#�i �׭/#��1`���QK�z���4�^y-Kg��q�����3vz8�
7��D	 �|��/|[���g��L�^�cN�#׫���g^��/��V�%�Ⓝ�ά(݂�"�վ
��p
��L��!	*�ǃy2��	c���߾�x+����E�e��;Ť�sNqDȰ"ߔ���0�G�"u��t��k�ӎ�x�j�e�,��R�L�v�~�/�$w�������| �h����t/Tկ2s�F���5|g����g#@��*��p=N�?Gk~��*�Lo��i�����!:Î�x�tIf
v�W3;���G�҃�uݕp�q߲,;�3�����ޭ����()��5K��e����l0�t寛)%�}
��F�Nc�)-������>�<��u�<>������Zդ{Մ7�g&�;q�?�S|��A�r5�	�'[T�EA�/���<�exN��*3�kF>�SL�M5�٪����kye��ɏ�#9���u���߻U;o����?7�G6�v~:��ݰ�n���?Ќ�Wr7���V�C�Ta^
�A�t��Cp�̚��k������jQ��{�ԧ{ޒ�b��kt���Ov��Y�;�6v'�o��Z7Ґ����2���4�k��>���A��t�>!�li�"���"��y��C�\����~4ݑ[U=w�+k�K�7ՙI{��0�/uN1��ŽV�:��9���=���aj,Ӡ���	 �����؀;��{Ey�%�e�U��;	Ǽ=T{�g��ll�Y�ϐv�t�C.KܹЁٮS�Y��d��<r)𶀝� ��*BI����,l�(s4M��]�J��oLn�lG���� ��w�{�ڴ%��F^�]0��������J�~�C�o�fo���~v~�F�ч�z�f��z@`��:9������r�C�s����������t���.�����؅,�����S���̙�s�ԗv��p���.��M��U��o6J�ì�U˜���J3g��4�]���4�[���!�;���E�� *pq�11v�3�����ҥB�/֛��?sd�l�����e�x����6�L^q�$Ȇ���Q��V�ˢ�*Y�H��d (fH���92*}C�w.��W�*����g�X.6{�R3��Ȣb�=��P8C^����C�v�qL�ªh��R)69��U>B�o�����[j ��х~���@����wY��'������_k<�6,��s��V�=� q�"�8����rx����^��|Z�L�4�V^��g�D5���"�x
�0��gI�ρ�(��.����������v������v�?T��䰝yh;\�o+a��9�&Ө�mQ{�˫�OŖ�w^ϻ����2z��+
�=��=�nt5���|E�D�>_Ӳ�,�?�vz^\Kcu"��B=�ɞ�l�v.6�.;��m�H}ŝ�������k;e-���Hs������ő_/�>�%Q��9����R�L-j��*Yt	F�`0|]v�s����i
�eIy�+�[?��\󒞚V�Q�⻱'�)-�0H݊�8o1rn����P�j�v�x�ko�����U"�f;!?.�7��SO	����$ϙ�Q����`sR~'���x�q�/���#�x����ٲ��w����e��윜k�z�d����� G[�n�{�"�5ۙ��7���e��4kҨS~ݠ}�R���c�΋��*������8���?\2�׸���Ιcj�V듥%8���/A������e�af���:�v����o8���]0���[f��^jE�YTo��9��pc��ʾ���b�W32�*�`�6V��NúE��W�[�5�E��3��VB�Bj���F$�$G
�����Jww��KF�����ހ�P߿o<>���׽�u^���sϹ���{b�l`�@����؋��y����k��^f� n�W��-�=p�S5t� \����E���C1R��+�*x�kט�:�}�O ��|^Pz�ܬM�qu��(��;��.Ŭq9�%a��C�m[�;�[q�;����[������M����[���mY��2�<�4!�I̗�o�Ń��r���F�K��=�Lb`L��+�@����j�j�8�0��<�A:���+ڡJ��p|���9��lV����Q u?,���w�̏Ayzf2�����K�9F&T���M�'�wx��Io���G�6h��.	��X3Mz������?�Hñ�~Xc�$�B�m|W;��w�O��xP[^����zW$�9����$K�dX�{2'�s��8�|��>�84���L���Zr�țH�2:t~�ǻxxl2��+ZK^t��P���j�?j���gt��D>me����,SE6w�ЉA��,���uƕ~���X���}+�ߥ�9��o]��+��2+�l��1򶙀�z�O���age"I�"�f�� ?u��B#�G����XWY|p�����P��vH��_g�OFX2����MHS��3?
fȔja��fJƫ�Vm��8gN�4�~a�>����f�i f����KJl淾����?�0�(5��!5F#���']CޭSY��)���ӈb�f�¦̦1�!AQ6�7\�(�=�T�a@���9+	�u�uF�����܇lN4|ڥ���? l7��4YQ�2&8�x��"cQ�'y%<�}\^[Of�i)n�?[��Z�шC���� �R3�i��ڴ�ʏ������eN"P��_�R��R̞l[e��(�PZ1W'Gh��[+��-���s1K<���d��_���I���m<�H5�5T\1L�"�&)TzJ*]H
U�%:��CzM��P��|����z4FƆͨP�x�'���@Dd��JQ�&.�b�h�<��,=��`������T�vE����R-�V:r��ÊL2�_U)��:3�`��,�ZQ�O�~ՑZ����H���*���Bi'q7;1N:�YM�	-%����J���l7���{��X��֙D��Ż#UlA�Lu�F\^���a�UX��ū��5���-�q�9P�������kk��MBY*�3nh���P�ԃ��z�K�Q�FH��JJ/��h!�vn
����R�ψ?�P�p��Ti�M�G�or�_1��-�Ŷ���7����vz��hM+s�����B)k��J��c�q
l��;�f)��R�<n.�W����E���8�E˶�j�	��Iv��:gyPuZ]gMY�pL����,*F��+�A#����j��>fE+�t+0מPζb�~>"h�.cĩfV���|߼�xew0cx��ƪ��E�ז��;�����G=��`�(��^�y~7�{}}S�l.4×ҕ�]�q�����5�Dv���� Z�b?�mt8�T��b�X�����FXw^�.���T����NM*�f4���o�\e���n��(�(8Z��C�~��Tw�J����,|UJ�J��}��g��2�z	"	U���~�CPJ�=7�Íɖ��sC��=� U���\���"�u�Q��FOl���qy��~��Ƶp��{�HG�p��8b��0��Y�oԁ��_�p�&����X�aQc�Ƃ��ǏΧN��W�Z��ȯ���t���>WV>��X���Y��`Ŭ�*s��~އ|��q�8�3٥eTdӖNm�L)��'����m�NX�hr�]7I�����Y���C�}��H�E_���ވ���1�=E2E��	A�0���J��}�-�ePڑq���'�����CM��O���?��&E�LoiD��6a>9[Jw���q�a'�3��.c�y<�<	�����Θ�wa9�����~��yχ��4�藡��g��p٨Q��,LH���*�2FՑ4��]�����5V�l\5�Ͼ
�
�p���	�h=���[c�.J-�����N�|c���x�!�n,�O"o�Ifl�Tm�-�� ^�&!kD�������x�Ȟ{�m}�<�`�5��#G"����b�|ԏ1gW?�$�(������4������&��YHx�S�<<
���Atÿ�2�}��Ⱦ,�S&A�5U������T��-y��ڊq��*��>�> ���!��RϤ�,ݙ�~���N�u,��sD�gt�[|D�۲{�}9�Iu����jֻ�nwµ�BpF"�F��	!YJz��k_��^~ ��6m��Nhr9R�^y�:Oc��b�<�Ps�Bx-<Ur'T���B))B5�V��q�S2���+5�m��-t��C�����ςxn�ܽ�5�b|��Eځ�;)�OB��'� ֊�S��ܸ��I�U<�F@���g�'[[/7Q�Q�3_��w�v"�q�^QЕ�0�'��{^*�T�����c)fV?��*�U���[K��P��띮����;=���^]�7F��� 7�x86hۇ�ǎ�^"�*J���?�F���?�\�eՙ2<[~��x������Ò����� �a �$��2)�0l��E(�/��P���Yfjţ��i ����̻BU�]{�hQ�K�� ��γu��}Ղ�����uƑ�m>y{��ڂ�=iid�v�+ʿ�k�`��Q�j�̚^AQk�N��2m�횕� 1�tQ'~&�U�
j��� ���u|���%V1�$q>5�Z����<N�q۟xZ@B;I��	�
�$���ٜ^}=��5�*Y��@�=Ƕ^`��d�l���C>�-�m��7y	�nR��t=|=�v���۔�7��Ѷ�mL�ɭ��z;�]��N�½����T/7�((4$=��ۭ����d2(O\Hҿ2Ȳ,���=��M�q$+`�/p'�DWk8�D�Y��q�eyU*a���Sp[[[����N�?;o��i*��w��[v����98���v�i��#ބ��}aߒ�7����'ͷ�׸C�^�R�9r�Ql�'�C�zR}�Γ>z�4wm� )b�#�#���RP� ��CwF<͡�Y�W$r�V}R]�T�D���_�b|PH��)h��_�9@0A���ϼ(y�_�,ភ,Y0���{܎9㗝�J(_/�)������x$�7m�z&8�|�� �|/}�酻K��;ٞ���Ӓx�0��u[�5���%�β"���DOx���b��9�H�\�сî�ae�3��3���l���ʔH\B�����}׃r��NsJ��j���O>'$��7�z�G��p璮���nk��/̗��~J�]*���+6���K�B'A�fR��$���������'�8��
��p�<*��S�S�������w��d @xeQP��/���j�M�s�W"�v.���[k�Fμ�R�4h�[�����%`/�pb��b���$0/����(���3c{H0�G/&Y�c����7k���fl{�)��z�vz�1�8��~��<�-��itFKzaj�M���V��hf�A�s���A��\4>�x�|J:qV�
��S��G�$Q�ް�6������s������}>��1�Z���׹�ş!M�������O�k�n��Q0g�*@N��m��y��-}�-�!�vƆz�w�w��&s��ʘ��=�|�+��i�`-��������My��KE� ���$� d�����C�+�ז�Ӎ-�|�l��(��W��:��d]owI.YC��94�D�+OX^kɞy(�S�!�ͷ��G��������U67���Ư:��kխ/ ����Z�T�uG�ۍ�ӫ� r>|h�����P��V>a��+d�+�ҋ�6�fƨ�������v?d��s\��y{_}�E�](�()��4��)����������4������i�ɞ1��n��~*+
�N#义�@T��D"vΊ��@�Y�.�y$����Y�S�����(�Q���*R@�^%�r��s�H^��wb0�"�'����~f#��;k��c�8�,#�]�>���n��E��$7�N�K{��ΐ��r�����˶e�6P�D�Ojon���~x�����?D#�9��[�H:^�`O���%��^K�	npſl�%�0�Gi����&[��`.7�y8��if̙�������>BS�%.7i�gFW-��G�.����-+3�Q�[����@4t�x����o�����Ic��Y5I&o����"vǆ���糿�ܻ�v�6�m������?����v{|��eW�` ����FȬM��g�2�oc:8|\Vy���X��H�T�_L�5�"11l�"���ة��X��t����Qӟ�@��#�ѪbLi�i�g���&.�y�U$�w�:��eP���L�+dј5m�Q�~N���3����2S�O�͏/�M�B��]$GK�.M,g+���m�f��M*�Sb�7+�-wqi�4�U�o�{�G��n��������P���i��h��I��ǎHIheK�.14Q���}>�;_w�2�[�̟�5;c�;�S����m�w`/�'6�:�9H��5sb"�ؓUO%}My�l���35�X�O���i���豈3z�䀅0ywku,j�U��#����ʎ\��懮���7[�^�����������x�/Ǌ�m�B�u��f�Ƅ;���kƱh|�X��]�Z9��+kZ���6��{P��/r)W_אB�3�M]Z!���G�f��� ڒ��h��I�v���"=��NYx|���\i#b*�h��'��2 �n�O[����?5*��֖��*���Z�*��>�^AAӃx���WT.�C���6��2<��m�,4bZ;b���7șϵ\�m-��4Ɋ�ۋ��(�ppY'Jf�ݮm$ߊ�tT����Ѻ'p�1�4�bPa�4��9gK���M�������Ⳕ{ĕZW�J�W�k�"���w���J+c�W������<�"�a�M7�I6TN��z��)~"�����7��X�(&.w'	����"�~j��a��?F��n0�t�|_m��'�23;ݦ*A�~ـ����U�|��Ҋ���+��~)
e���Ee��M~BM��z���5/w���?ol��e�`C���\��6��N_^]��H�:H�;�U�@F��;��%e�=����+Pj��]�D�0��0<�}����d�j*ǅ�^����N�!�F�1�����1��u��A�Ȳ�:�K U��HX\F���5�6�@e�8��4jw��#|�c��d���N���-Tf�,�*�uBT�f���x�\�;[��!�)M�{*|v��j\�:�Km5�ba�jӟ�=}d���;��?|k�O
��I���eY��2i:ZqI��GFF���J���~�ܑKF���9�=���K9�Ǻ_#�os1?�J�x|&j�*���~|�|;��)�H�����V��-	��쪵ǉ.�/�I_"8Dqܿ�0��&ʦC�|;�M�fK�z/�IH4��o�ۓ�?6r&q�^�=ư�������
ֆ��ğ�����9���=hB�H���,��O�����=Ӿ������R��x�cV�����Z��HR�Hy�/�ޑ��+(ڢ�
:�&n���~�oQ�i~�o��j�@O�������n�h�KOu��㕺{d���#�m}��q�Vo9��^��lY�и��{[բ�����K]�#�������������l�+}�t/O<���( ��K_p�o�[��f��)2L4(%BX������8j��S[�a�|/3�Θ42tugm+�߇� N��� �5�=�8�5S�4>±�^�|."�*��=ŞR�2+�[��3�i���A��7�$sK]����N�?�5�n�xc|u��q�g^闕LM����s[��t���s3�W��*�e�wJ)��ha��ʘ������r��S����H�#������z�#<�koI�\�P���h�e���9��L UmS��Yl-~���&�ilq�Б��~}�a"ՙ���� �Ξmi���WǵO՗��Oc�9�q���E��5��*��[R�� ����?����O�#���(�����Y���r�[�%]��r��'��"m��t�ʖ�|�q7��l��u�%�$D^�㛏RTB���$������f��g����tPW����	��yB&æ# �*�L����?S�?������Rl�R��%J���K�}w:&Vm�����<��N����8ߨ�JW���pg�����4S,U�Wn��:�}�����u,��gXWCH�~m<��'�ʹ�Й���Ɣȶް���6Qv7#��i�ǜ^��j5R��`D�^@�5p����2�3m0̈�Y��%�X%�t?�%f��if���1����l��O�ҝ��M1f��=J�S��{�6�n�2
���>�x���7a��ڃC��'�ؗ	�s4�'����,w��f�%�2|�(sT�#7�=+-��E�/&��/*�\��n0i>�%Y�n4֪��]L}��r�\��s�}O{").$�Oڧ��eU}�mʮ6�O�Nߎ$,>(�Cr�6M����[��7	a�ת���\�����25G�Gz��0�>����۱񢺤bL���ӗ��'��^ZW8���:+ZN����lm����	�5R�cɲ�u:Z�~c�w����gZ䰱��cj���:���pҭ�B�_���밓;���Xs܏F#xj�/%q�UZdBǟ�@�J� ��c�@��sV/��'��"��W�Pd����j�n��He�4U���Sꢜ���w�uv��W:kN��>���R�<a�1�nx���#$$�W����S~�zԫ1E�����	*�E��(��v.�#�;Ub�|f�:CZ�y8��i]L���y\eHv(���=�9�x��u�-�B��*:�j(6Dq���̴ۼd�I���,���9�& �)�E�~�0]djj�;RMx1��D��e�'l�Е��;�xF�w��ޣ��m��ڊN��^.�`�ck���#��̻+�Z5��x�l�o<�o-�]Yc3�l��k�m+�p^F��"�T��ɯ��Q:�D�5�^>�M<��M��xn�f�9c���(꧓D�C�V���A�	�5��g5\�/�tb�Ni$���z5gU�~�ܐ��e�m����t�&��y�w(���}n��[d"��}�FH������(����9�mka�ʏ#=�UsPg#xd�R3�ˊk<(���jp��a�<��Ύ%?o&��~D֒�R�ȇ��^���)���>�Y�o�L-�o�{��$���NTf͛v^�Z%Ia��M�ly0+��Ix2A��J�T����i��q-���Q�Ɓ��[O�Ù�`�Y�X��w�f���%՚F���ᡡ� c�Ӥ�:V�￼��X䔎�h�����N5��,�`9AQ<jH�d�>ƛ���5�{�J�R~��.R���S&E�Z%bV�\3�� kW߻s��D͏/�^�}���;u�yd�x����bo2ݠ���V�W���t�/$������5�/{bڝ�Q	̰�O=�c��Yl7�$aV�`P��h;���7f|)�\�y�ta��"�<��P�!�Ea#X]'l*6�2� 7e��b��4��^���Б��b���T�x��CdC�F���%Rvc7I^��k4�I�Hc��L��r*8�=IaѬJt(�<A��&Gl�!ˀ�#]�ᱪiVKGQ.w��F��j	k��}�|Dݣ�r�ݓ���l��~���L�~Y������2eqG��䱿���[�~z��j��j����X�)?r��5�I��\~��1A%�öQ�x쳨����h~Br�Uf�ؼUz��$�i��i0��Ǌ�D� �;7h��i�{��`j��Ng���V_�I~c�RC��/��s%�Y�Şf.������T��=�n�׷��x%��M	Ij=G��3Hb��Z��?��8��=U�
üx����Ӹ���̿�
}�|8��56AY
��K�<�/��V��]l�c(ސ��x������N�^"���.wo-���K��U'%�3���N5������=2�x�\��v�@�a�wT��t��-��`����+W:|���&=������iydy[M�#N��Z+l���%3kVm��? s�E��5�]�[8��p�a$��l�[�7���w��P���.�:�ĵ�"M�Ү#Br_����w�:|��No�"�� )-���U(�/%ѝ�8>M?�vC�>��@���_�Q�t����[��n�㟓�X�m�r*!�ʶ0B��[��H>�y�uvޭX!��!��� S��6ש����B���
�c^�P�Xp��R�}K��w���JW  U�����Gw�P��qg~�q�H�Ȋ�&=���ڝ����nJ���ė��P�����a�4�準��=QUc��T+:�.�3{���d$`3�RX8ۋ�	=�&l��fH��TȢ��y��O��� ���Q`��N��S�Q����i�^�5�w�/�~/7��N`L`Qk���T�����)�����& �ɤ�8�!��Q$a?��R��.��%�g�k}�������V��C�ɭ� ���]�Gf�tb�$`�]~P����]�b��=D���OIK�:�"lش�'K\8�ھ���LѢ�ݎ�g5��Z���`��g
�<�G�bU>�nL��l�fP�ƹ��R�́� ��/�����e��[kw����<�򍫠%��=7ĝ�l���H�b'��[��uڂ@b���7Z��t`Գ+�<K����n�(��Y��k���Ѻa�S�D�v�^���n����Ƣ�H���[49�U�ϊ��L�b�ê2_� +���
�+:��b���uuhKq���rk#h���M)�2$q[�]b�=���徜���4rh�&|a��{lh�]�6"e��M���+3m䅎O:�v��ߧ,��O�e��ȸw5=-�Z���5�u	�d�,�����bO��>2H:B{�&׽���h�xQg���$�~�:��葮���d�����9u��#��dSzŇ�	�-�8>�fe�Mt;�5jJ:�����#�u���Z�R�㧩� �� �f�^A�G�� )Py����4�����x��GH�U@ͭu��;�D�%T�-'�:
%�W�T�<�_��_�hD��;��,���@����Y]��_XN�"�����cf��^O<���&�D�m����ID�V����S�쬐g�P�Ő;RQ�u��5�'�Vb"�S��U�����b�����(O��C�e��<]�|�����.ɼ�V��ռ�F(>�#��X`*ꮱ�	��0���>Mi�g��2�s�(grN(���1��?�"��[��oށ�e^�g`sI�aV�b[)2�zΎm	π5oE����y�w̪�����OU�u N���S1���%�a�뿾.�dM�{֔pel���j�	'h��pN����ޢ��|oYݗw�&.E�Z8I�)į��������[��5{u��,�FR����<�(��H����8e��OT��������d�x�m�{P-Oǈ7�K^���BC���ł�9���)���:d�R9u�ǔ�C���5xIn� h�mD��;r��l�����=�w�ȷP��X&�/����դMx^���T�\��i�E���p.��Ju۫2v	,�ȉnE�mѴ�j�h�[K�g�������[��k������:����K��U�#�w)�c&z��Ǫ$�I���\�Օ*�o��n�ص�(q�"@bͽ�w����_�	���骤M>���ګ�ԟO����:94���Tz��K�>�c���@�P��XCq��h��}Z�=UK�G��S;�,y�3͍&������6;,���}��"����j*|�/�X��Pb�o���\�5Xx�aDc~���X�X�X/���;Z;��.���B���m�;Q�8�\�Ep�����UT�meo4��˫�Oq���A�"�{�~:����k��C�pW��YXq�[�eo0u��.;8ܯ��ϡ[�n��G8�L�e�)��֚?�naee���zK����ȓ�O'm��<�Jg�I{�Z]���{ځ<�u0�G�"M�/�V�Ty���
�ք���9��Sz�R�e�,�-�y�E��r������We~��\�Z�YG��r�D �!�}R��c�s��C�d�rV���Q��:��'E�x�W��!�Ԙ��k�M�'B1G�&>3k�2�#4F��i��=��¥,�aX��������O88�����H�ɐ:E�������N��S�D|g>���+��rیݙ�b�HL#�����:��E��L�/�&�R��>ʼ��M8��2�j�^[�yqF�$�r����#M*��wcL�M?��</RM�@�/c,6snډ�d���x/X��yd�af����S���+:H�(5������ŞR�1��!�u�(�j/yg�����C� ����p�բ�\�.5������(ђI�[�ފ��r��!Y��1�醗l�ɏl���]j~�A����J,�{�W�J�zh��&am�X��ݙ���o���2s)��+4��97Rݧ��9�.�Η��ܢq�ɵ��<��d������TX�I�D��˷��>�D�R�����b��ˍQH���ƩY	r����,0&v�\�
KNH_T��T�2&g�:rj�;��d�G!*s^�uа=�4�2�%��O�g2߰���T�j��q��Frf�CU���D�G�pzS���׻���""��[��,�J��蟅�Ћ}X�z�H�`�(�j�hy��R�<��KIۓ��&�7���ٕ�3r�]��n=F����H�YW
A&$�B��5C�����b]6�����=#��߼���ﲳ��Fk(���:=�L^��x&u��A)�z�hT�J�#�XE�����`?���z������rr�cz��͘���7Ό��y?��u��P��c�Zſ�%/�zg�D�3��.+��0b:�<�������D&P���tZI6�����]p��$?>^H-c�l�[S�M$�`j2��j���%A�4Ӂ��7�})�۪��ϟ_���[�����<���,,�B*��`w*%J�Dx�6V]�I'�X!}�F��9�`�4�H:W�W�I)�'��f���LA�As��I��溻�/�y�?������Xn�N����3������P��/�-u�(�{t��{Պ�C9{
L�.��-X)j���')�� �x ��C�,G7�5��� X��ؒ����!W"W<��P ��r6M�/�ëټ7��h�Q���}�μ�wFᝬ�vt��0�� i��a}�|BM7��O��O�ioo4d���I����WW�	^+��Dk0%����hWp����g���r��Yw�gKo����G5�/�t�~$s/�����<|3�1���0�D K6�����Z����-�R����x`{�:��	CUC-��',�N;9Q�mEq�]�R��[��m(���2���M�\<�&���q��Y����fj{q_�h��{i8�f� p}��[�n>o��o� h>��&?�������O[�+gq�������)�T�����+h��⡿�ͬ��(�uk9��������,|Y��(�h�	�����9�>
������C-t�MЬm*��]1-�%���f;==��p�%f{c������)j���c)��Ei�w6��滔!�d3%R�l7�Ή�-0��v�_�����;w�z�����8kz�Ii^VY �b��G�Ũq�N�d��#O+}���[��n!btܗI��
�&h���4�\�4�Sn��I�1{�VL}#{<��i���䣶{\���
��Q��n��ߚ�:����"b�;E}�	5!}�K|W�Yg3W�Km�I����͐G/�W�d��WE
�O6��&$���V|- ��X�����O����j����;M~4������qHC�o���7����
K_�~�O�X����#��y����N��ȹ�B���O�8�3r���o}	s��N��%��YҼM�72�Լ�'��w0�U�'&���=����?�9"��Hk[�@f��|�_C�T%�÷ǟ��e�Y���
U~�\0B�]�m�����mNL��������38�~���vr��c1��ƃA�ԝ��/�oI�ѐ7�8<*��\#�{of�L$�=���������:���׆����Ί��*H(�#ض��m�!�\a����9J���5
�����Im�DJ�/lQ ��U�R˜��<������	(; �6�t�q.�9�
CZ?8�=tp��+��_�&)������0/��?�4��x��&g.�FY�׶7>O6�U�߼�I���X�������1��_�]�r\ƾ�^��'�\�q9^W�?���7�QI��u�{O�Kw�di���|�S�s���g�o9 M������=���� )��-Q�v齠|������=#
�op���-��F'Չ4��)�r��w��*HS�L����PK   �<�X�� �f  y�  /   images/96fabd4d-0b16-452b-94e2-688cfcbce531.png�	TSW�6~q�i�2*VA �Z*((�'A�0I�PQڊ"��"2�A@D �A���9�s����������f-���s��g�g?���^��ݕ˄�A����F�<�-Y�X�����_>~K��/u��A�����������t;�d��y�����)k�h�>s������mĀ�0m�j�;��k�w27���$[&f���tt��,�ｦ���ݒ�_n�1�`�=��k-]|�!so�O�~oy����B?I��l���K=�w4��؉#�[^����c�}}҂#n%�@�'�M}S�L�d;vg�|\������zƺ�WOڪ��g����VW	@*<�6++KK.��6��{��4紧���;�쇿V=漘5��L������9/U�c��r��;]�[�Ťk)�zj�]i�19I��DU �ƻ�{
!�w(;\Q4�_v��ͪ6��![�V���1���|�;����0�j�t߮9=X0�B.���L�0�C
�17��p�d��ۉ�� �n�=]>�����A�oVtɻ����1�Nj���v�.&F�3T�gČ�iL��S\\|����7=5��SK�����,�2���؟=���/ʖ��k�޻c�ׯX�p�@|TozƬ�N�Q�TcIx��z��j��xd5���:ﭛ�_��cz����5��V���D�Va	-$���E!����Z�����n�\6�^{�-��0~��ߺ*y�MJ��_����s�r���0�Y&Q�wNउLL��V8���@�%]�A�?���z"᫇�\|G�*�ς]��q�����"�"&"/��M>&n{T�=���j;��{#�-���~~~�ѕ��Fd�UD_��a7�rQ�2�ۇ��.M�H��-��y29�H�Wwg!�
��YW� �ѕ�=�QV$_?�l�m��7s���H/ds{W�z���]��Z�w H'z�S%\���4����_$����Lz켣���y����a����vD��WU���u���#0�O�qb�П9���!�������@!����^�}�{�1�sN<rĂbH���Y\n_��e}�NM�*l�1׀w95�����k�;ga�<T#�B_��zu��X���|MPb�[{��O�%ot������$�u�B������)ڛ:�F.P�9����3�4���s���,�D��Y�!I����I���0\��4�����2ښF0�K=83�jLӐ�OV{�;T&���{6��mr���n�9��2�fq'.�ZҜ=�l䣪��5��9/���ԙ�6���y*�w��,+%UF�lr�M2�]y��]4Y�)ˬ�ޅJά�)N9]��� SD�,���.����^��<7��]����))t7����|���e���\I⤌�p�+�4�m�!cE�Tc�ۧ��O�����`���4��BO\9
����NHk��<.Cȝ�#i*�y�YMMMK�,9H�l~}.]�c�����86VY�Q�榆�,���\�Ǉ:$bBU�Y��A�C*�dz�gHp�x��)q�8�;[� 󰱝��l�W����\l�G�.��+wI�l}��v�;��a
�Ӎ�Y�wVA�x�˾�h��&���@{@����ւ񕒜9KF
�-�:�U��]�V�ç�2�ko�sn��z�ah��d)����
��mN��e'*�[�rFXOX6�[�D�ħ�!L�iG����I�P�qT�G�}}���{o0�N��s�x"����Y�f���]�<�RdX��~��cz�Q�t9�H-tRv�H�N��=cn�a�f��fk���[��?��B�eΉ N�]{��&D������!]��Z�=q��o��e�~�8'Os�{'������r2�p;�CD�zݽ'i������܁�---�=���>�|� �"��5�͎�7B�=[��_�K��΋7�d������f=N��s�����0-]K�S\sXˁP\uz�����UЉ���4Y���xM=�yp�A�s	-b��wn�ϻ^n�34W�pc��Y2rEA�.��`�{C^���;UaG6hsl��)h�(�Є��G7U���d]266樫m��ކ������=6z������-�Xw�a�z�Rt7� �$�](�B���-��s�G8��YhU�� p��r��v!(e21���R0��~��z��F���VnYM����љ9�tM6{�9��iͿ��*�&#A�o�g}�Ɲ�q#6VL�┘ds_��$J`����y:o `��/wti1c��?r��m'^$m #����K Q;����ֱ{��1;J�uC0�0�{��v��h'a��a̧QJSp��W���=���{ ������q��"-�l6ȗ�2  H��f9V���
�K�ȋ@�h�
 �d�W.��5r3�{k�Ó�p'u_�"\��F�V��F�nz���CF�����}zvNMu��x4��<�5b����Ҩ�,ض,���R��˗/�2^��o�a)�\�X烠,��O�\	�����*�W��KJ���a'��d����H�4�%�U�Y_��DgK�TlB�m��E���iÅ]�Hٶ�h]�� �T/^$R� �d����X��\����^9ɪu�uM9�![%� a���M0fJ�3�:a�f��A�8,d��h&���X���dե�fҔ#ybvz V)��R!;����2G��[�'0B#Y4͛s��ϺC��@��l����N�.���� A�b��(��g�H����\U�r��ٺhONl�Y����K:�
��g��ӱ��X��G�Qn�Q���Vu�ƾ��0�CzL$�%�j�M��tG:��|�2g��_�����~z����' ���p�R��X%V7D|f��fx@^�
Ev�9�jN1���v�Td紊(pO�#���sl�T��c5��B���Uy(��&�)S��&�\�$Mw�s�zn>�	ZjêkG)��=]��wX��JQǖ��������nE�?@j�����}sa�
?ᘗ�i"H��	T7o��+�6����(g�׶s%[����圀����DS��Z��\���y(Nz�DO1hXaD�J8�\�����;w��������,É��6W�i�����e���|�>�@�	��6��M���WC9ɵ�o�3L�@a,,͠D}*I}��4c�r7Ǖ��cNZAn�Ct�ׯ��}��u��9i��
�R�B���qW����Y|��i�κ"��ۦ �]p�o��	HJ�;=ҳ��8��1�*Q�t������p��q�^9ȕ�6]����Ɯֺ�'�1tqV���"(}��H��l�0��h�0�5.�RO�_#�#��gPrgpH�f�z��`��زT�c�T��$1.��Y�( �(�t+AzvI���)?�hD|I��Q( �
++��9G��G�g[F+~����&�К��f��1���g0���G�D�t�jDG�����E0��p�S�}�]��-oQ��=BPbӥ$]�n����E�x�E�.�R?�Y�CN��k��l	
X�É" �XM6�����q&;�Z�`�������D�~w	4��<q���J�����uϩ2!���E�5��(�8vu_�q�qL��5���V-; �+
��cb��03�E��w@ˇ���1�̠�&5og�;8��9��=�N�Q��(�q������H��9 �)��|����ŵ�#r��Ǉ�z���s;�EͿ��-�PN[���Q�۶�:xF9Ҁ�
��D�x<ݲlf�9�W ��xމ��=)�<ǀU�_p"��0T8foZ����Ć8�' �U����3�ј]s" /|ŵ���6��i��F�Y�h�֊���n7a9������l����52�X����zw�0�T� ��ӳ���K`���/9����
�N����
/ւ]q~�4�ڠ���I��R�zU�R�%>�`K�e��@%UI����_������FI#��o[�z#9oҽ��w4h5�o,$�K��úW3=^0��b��'��պ9��՛���'��A��[8�����֒P���\��
q:*��WO�����5�Hl+К���<u��l@vyV��B�(��A)�ưi6���WC�����6)^�� <�]�T��:�E�y�K��DϬ�ǽ��5��;��_�ѳ��)�N�Ɗ�`�p�Ig�(y�n ����|+v�S��J U��)�q���g�H��} `��\n��;�C�<�����Xxt���,1��;eJ,��-����ӢI���^�%ڍ�j�oŵ0�mn�$�ܩ��(����wS��QʨfĘ%uf�t�a�ujR2�H�tz�W9*3XSQZ9�7A��W�1!�?#����Z=� T��'_���vd6��`����Y1��y'��;�'C����r�[΂̉FrD�:�(дTm�ZUcBgᓽtV��%�Ŗ���m�����55����mQ2�����sYuM���~B+�u?���=��}"xl�7i�#������I<=��.)�{�z'�[Us@��a�q�Ғ��Y[Q����I3Rr��D�O�ƺ�61�LZ�<|E�Z�C���2������<F�`���F��֚��N5خ&�^�w�	U���:��٠�Żkw�ZE�\�ʐ��w�����)}�	�j)��Vs�ۊ��X�ЗFRfӱ�3-���{�zb���Zw��=���͠���(:�w��v��qqX�M��|���-;������K��֖K��I��YV� Zi�q����c�|0q�l������Uº����4@�5D8�i�����6纜�B����pŮ�D�שr����錩�<�B�Qf1t���Hm�޴j�e� XUL�b�'\X}��O�
L����i��olA��(�2�~$Bc)�-�9#P�����{3��r�t��mS�#������Ps���D�΂��h6���ޓ��y��Zzv/�(��^Lb�^����0؝F�Q5�3�r�ӏY�)��S_���ꝰ�m�sCcb>`:^�Lc�b�7:ekK���=Un#/�
�zk<\Yv(F����X!�{J�����zW ��t�s����\ˎPF�/�&�(�&Oh�w��a�<��6��B�1/�'��ş	�~�rl]���0�����oA/i8��lz�E%na^T���dd
Ut^q(���M�����-�̸Q:bA	z�[C���;D��89�0�zq�!�4g��gf|uw�4�4$��.�I 4�?;[�Y��[8���9S�'�BHjH����b�pؚ�����T��1.�`5f���KI�YWԹ}�2{�~b#A�h����2�\<� �20�VۖA"v�?7�ۃ4�"��������iP�p�"@�a$;�����}�*n��� ���d��-��'���|�漾����u��ɬVKJ*�I"ܾ�Jr= �v!n�r�!�Zܸ�Q���D��3+'KnII�����(Зc'��1�"����e�
�o��0�p������d�.�)� m͟��H��#�K�9�%��zO�nS���Ld=2�1�?���<k� \�������y�����%����p��� �U��[%��g�V,�¢��m�Ŏ�Vg�E�:f�W�<ȭ,"Qs����ÑFk�څRh����9h\�*3����������p��t��|�ۛNZ�.S~;+��p���bkc*��|F!�=*O�M��nM_�B�����󲹎���[W���tC�t5@���d ��P0������
*<�L�;U��M5���q`}�/C�p[�ji��kd؛yy�C���`��$�S�[25����	��c�Q>�h���\��	�t�	j�{�Y�5]�<�y����5����� l.P���,�䠔�f������+�\8-�p�-�e?A�b��d�"�(ǫ��{u��#�J6]���pݵ�}Z�� չ.��8<�b[�,�&�K�`G�+i�ۍU۱��&�'�-lϗr8iP>�A���P軜"��Cl�-�ध))��+�A�͢�;����,��tfm!��Ť.@ڲA���y��w	p?|&��PG�&���ښ��)5�Pɴ0��&��r��}λ e6)5f ѪYط�� �0Z����p{}��v��!���[гVШ�y!�;hY���lȲ1���y���������"e~����Bз�M��:K��������էxJ�3�Y��G�WB�@��P�IF��L83�cq
�֜�.*&����0�lH��Y/l� m!hi~mry�nZ�����iƞ�2s�{�[8#]����&��2{C��y
j���h9
�I��!�f�6�O��	�=��(T��^7Y�X��i�sQ		�:��AW�ú��d��t�v�%姶9�B��ŗ�}����4�~��s�) �K�,B�_�U�?������qnv�m`��ڠ⎱c:�+�u�&���&^k�MP�z S1�w��jȇT'�A��m���|vw�jD7�@O'n��o�VE&�8Fy�+k>{�84�Z��~����������?9�l���;��^�����џ�X��	?�M�!Yǿi�㭗�s���2���Xq�R���Z�^u� �hB�}z~)��14~��F(b3�\�e�M��W�p~z-`|�&��َ%�X8W�a���9�'@�?m��9���Ț��{H�A �-���7�PkVw+ڤ�O���oHӒe=��v�%�5|F�CŬ�ڒ���-Z�l���=�A,���ه`��S�X��<�ۛm:���G��}�ټ��=]8� ��N�e`IU�l.��c�hp�{����e�d�Ѽ�A)p��[rΕ_X��W!�����W���V�
o�ɖW'r�n�r22�Z_�o����<ӣ�ـ㇭�(ہ�ey��.�>aN�J����3S36t������cT�8�d��j����$P/1�P�Sߩ�4-v�'sȮ�CB�PMj?(�0'�����*e�R�a�l�O��=�l=���I���
FYb�)K�sO��t��؜�/?���d��G�il��ϒ���䲟Ӓ9�2u����,�E��s���6\ÏR�9���}S�{/��w	(���cЎbG,��/猋��s9�+9��W�c|�{�B�D�N)��>@���:9�T���s���J�ka= G�P,(�8�����^��~�I��f��ps{��w�����RR���0&y77�n��亨D�iE��7�C�i���&��@u �:%I�� 2>ݸ-=-w>���I�0ψ$�^����LX��x�3��M��(I���@+�J�>����Է
�Y�}��wKj�9���z�Ϧ��x�շ�2�Bt���
}�����ث+
j6�6��!�#�c7��ى�YΏ=��څM��*�s�������[R��쎇�:�Ŏ8'���|O�w��ʋ?���z�H�<9�:r�1*��ͫ�Z���K��&�{���~���bK���Ǣ���o���t��}��I���~���r1��M��BC� ]����z�s���4�� ��z蜝��J�L�}H�5I\p�N]e�U4CZ�f1��cvGv�4��c��B]�i���p�->o.��fWT7Թ]�vmfˏp��.�����I��qHPCj����HS�'�zqv�.ǷAj�}aF���J��DχzAW���n��j��9���d/����;3�j�H����<QA@��m^�΍�M�H3`�}��I��̦��ר@�J���ũ'XW��Y{��f�|`�=ˠ��t���-�2�r�`�0���F0ڌTz�Qs&�9����T*���A�i���=�$��P�ej�������|dl��qkAzzd�>�tU�4(Mk�48I�4o�Y��y/�GWg�]�Vp�I���P�c��%_��Ž���&���$��N:�ň��T�f��x0.�b�َ�m�Bo?||�l��Lv�fsj���q&j�2gaFeNP.�3-=E�PSS[Lu��el�x�U�G��}������e �؃�<w�r{g�-�op�q�����p��н�|R�*k��܉�Re}�n~�.](�b���"�7��΋���?��.�A�n�ºu��Gkf��0�ys$�ʻqL�UEa:��^_,(b���`D�ǰ�@^�M��\6�V4�xyqJ�!��Wp�R9i#����%��Ka���?�q�{��� ��魷�4�[����LQr5rb!�gÀ�n��n7���RDӅ=�,*㤪Ho3�7wgL�|.�(�0���!7U��`@|�e/[@'bz3/��2�Ҧ��ϑ��Nn��������j�R�c��p��>q��#c�hE�=��_�@�Ϊ�Jbe�?YPn�R���K��Ka�$W���­�I@90=pYP�+z���ƹ$Q�����J̪�Y�Kf��Fֲ^�dj[J�fC�K�+-�����:r�=P�r����Ĭ�E�=A[�eZ�P����]��4�pJWH���4LS9�49���5)5W>E#~W�A�M��ܡN�׻7UMM&�>�P-��X�0�q*��~��k�'��)��^Ajj~�D����TMu)Y04��4�`�aq����Lſ�D���R*���rnQ��	z&P,�=�������{�#���H�$b�@���&gS������1S-gf�Dʞ�	���]����	�������=�d���\�?�n�����������������������������}�.&F�?i��]��@��=�ֽ�Q���u�e�˙а�K�S�={����L�ym<�8�+!��B�qO:�;)����C�#�7j4G�$�I}f�M�K���`eb�Z,�G����#G2���F�&��뭣�X���!q�挽�~(��F˭�	�k�*�����Oss����N��9�6�����V�xa痼�����h%��Ω�FM�P���ƐK�ǐ����hh��Y�Sk��Sr{�ݛ{wwe~�c܏�n��d|P�b�Ӓv��2g�<��}�NIL���=PlK:�tAe�@��"
�>�u��3,�,�9)�QnsN)"rʧ������gML���ه�:��z��?��r�������q�/�i΁�w������[��ឍ�>���q��7�{�_ޘǬϊnR	PX��P�;��ҕ�5��+*�eC�N��]��Uי�{Ϸ�^�s6�]��M��-R&�:�7��5%;�F��q�2�e����%>����}��,�#Ci�}���K�����K��@C�i-�)�c�=�T�;��DȐ�9�aR���G�a��C!�M�N��f]�+�\�Dy�vf�BH��$�B���ֶ?�2�);]Nz�KIj��A�N�ZagF�r�B�i>4��?zo��Ջɋ��v'�F������
�Yu�+�ϔ۴�T�MLu��qvf���ʨؤ���x�>�Ŭ��
���{&�Ns�������� yG�@�|\\�����sg	��mf�ŏ��Ë����@Hq�G(��άoqs�e���h2G1����K��GK�Zf:�h�9��b�r_�ϫ����l�a1��!�8�}gggBL��p]�&��o����dd��O��o!�����	����@>6��M9�l+�R�r���t�����5�gI�Jc��������[S�\���X�i��
�M���*؜����
ͬ����
��DV�2��Z���di�(Qa��|��+�_�ϑ���b����:���w�����
c]����'��`��8-D+1���D�l�Gu���t������Kjy�ZӃ�}G{jz�C��`{Q`��%��x�.o�l� DX�r���	�%kwӠ����?���͇�z(��N�2�A���j��~�]�r�o��SU(/�'̤�ncA��:�O�Մ��?�*[_����G�we������o�v�X'�
�p�W�d��[\ބ
�( m���:��g�c
y�Ajq���%��M<��'�D����@PzJsV�:�^M5َ󯣃U	"ZZ��*h#��"���V����+)Dg�!��h3�	|˸����0V�2����*~����KJ
���R�k�7݅w/&��W���!������);!����
�z�_�m6�H�Z_+��n���λ>"c�|�.T��~.�kV�
���Sn�ŤƗ1�m+�Gsn/_d-7�R~9�O���m6����� B[�W]��-P�a�"�ٯ�η�a9y�u��-��6�\
Av���< ڴ�)WZ[F�y��4�T�o��b�_���	��#���ԻF��I���_�M�v3�k+ hծ�ry�ҽ[ѓ������n"Q5����ȷ���`�5�Q5���*��� [1�?j߻�Y��'���%���m!�91)	9����k+�P�"\�[!�{Q�������󡽚��MX�5��4��y2�G�������شC4E%��'�W��dM��J�Mc����׈ VΡP�W� �y�J�G�,fm���W��M����u������9���+���NP~�
A�G�w�$B$���)�������\�OW,�p~�8_⓯��_������_S�(T*�� (�%o!W� #.�R���s���t� �����s�x_����A�'`!���L�U0f]��`���J����H+㚗��w���S��.�<m��$�L@��J�t���L�"3��Oa����(*�Ȋ�����&����Z~��p	Xi��1 ��o�C�_q&���tij"h*[P}��FezO����X��r�K�׾_|�ja]���ѻq�YOц���.�:�A2N%�hVs��}�]����C��T:�˯*��O�7\�3E �(�ׯ����c�������t@�D<�^J'�9�Ci �<���V�G���ݹ7��U��X�������j@y���`<�!\��^� �C��'�'L���,�OM޺f�B~Ś��?~h�s�\{��|1��,�������pqۨ�H��0N�/@�t��H
=v��������d�"���[�������߉�K�|ʎ�?��Ż�F �EF��o��q��0���x�����5H�2�}n��Qa{/��R2�Ex3�>�+76�{��͡FC��ٜ�����2�U�?�/�����Ĭ��aS	��mF�N@�vgtEL���7��B��������� �]����߽�;����Y_��qtnػ���@�j6,�&�cU�ߋ�'^�k7�s�u_OO?�s�����Z�C!Z�Q(/n?���ۡF�w�&�nE͗M��F �J�Hg�{��G�@{� �ٺ�3��2�c�V����$�T���~c��@���>�6%%�0^W�r��k����ZS��8�oK"��NI0�`�ay�g��Ъ��o�}�n�\�6~Ϸ�M�!����Um΋i�3�+K�c���ʓ���������T��K
�廇\Y�;�����3��-��X��쒁��ݠ��������� K��ļF��l�H[�vgj���;-�(�Z��˩��wF��b�O��t�(\�14~9�z0񋔆�`���hW#�LQD�y�����N��
���o��maN�,5������6�@Z��ֶ������F>r�?;v�I�՚��|�#̛�M��J�
yvƆ� Z����L�]�l��i� �{��z�v�����V�N�U`@j�������s�d���J`���L�[Q�\��Z����3�B���嵴�g_\Ӻ��������hÞ�وЪ�H��+Y�<ˣ����$A��{�ױ��ة4l ���Q~��I0)z��#˿V��n!�����d̚���4�G�k�>��Ą�ؼCQ<8ǅ�����k��	�P�v�p���FLL<mwww���
�L!VXQF��-���1���L�]�r�H��5�3-h����0�.�5Qr��~D��Ԯ���դ��2<~8'9�����d���qu�� f�y��WA"fH*����w�&��.����s��!���ҒJh���ҝ/Ȼ���nnktuu�g^�#��_/**:ii�y�E$�Uxb�S�V�M����
�� edd0��>uq^���`�S���0�1!1������G�L�ə=[5��笉�/�_�bl+�<�=ݥa��h�F쐕��W9�p`pql��
㔞]݅T��6A���cD�HL�e��f@Qnb/�콙���i�)�!�(+RE%����^���%��4Co��j�cZ�OƓ �͒ͯY6W5�V�vy�G�?�Lu"�֎�y*��-4ճ�32���W����H����Ļ��&�����Ӵ4���w�?o�`PA��;:ć9(�#{wz?f��h~���
#�j�/��a������mll��!�~��.c��[RɕA�Lv��v_]���jޔ�������y�ӓ�!#<<���f�u�N��ț&Ԛ�e�g�P����X�)��4�_�!a�F���>�J`NS]���79*'Zd�	����Y���b4Pv>����������Π��(88�د]Y����v�l���.��LF~�g�_�g"��]L\�Um�	��������L��7=�Z[]]���zݲl/ě"I�I:4����W�^��[=��X���'E�b��3�+ ��V�T�j�_���N?)���c}���p��H)"��x�ԩ��1�'���J����Qߏ�۠P��
��l��ɧ����Jt�2rժU�Zr%V��°�����'m e�>�s���:�C�{��wQ���]N��	i��W�H�x_JE{J�f v����������>��Y�)fć<a��(�3�n� i��6�b0���-*_Z�����L��kaD��lR6DP?<B��mI��5C���xQ#=���. RGc07I#���*��̞���-�Q���>��(
u�А���^&&5����3^���Ky4@����D���c��@���=k�/_�4=��[v�����Q���Rw�Naˁ�,Đ�^wf����&S�<�.^L&���i�ɼ�� 0�$Z_e��]���]tfp��;�HT���5�t�>�[���Ei��#��.���(/+��~� �w>�Ԗ��Hۜ9�@R�]:^� {�d	X��4�1И�B�5��I'�������X{G��\��Gܲ��+
[e)})J�|~t�p�ATDdd�|�,m1L̕�N�j����d�j9,C
3��[�̙b�SB����]/^�8mo��^��99]�(�F92�%8 ��T���]�� ����ʾ��m�+<��`�U���3S�/F7 ���?`hU ��ddWWW(S��C�2�6e���dV���T ���Yb(TQ�=�Au7����툧�e�ff��U�ώD7�{�	����j�5xO����pU���(��熝�K h�v>�lc3u��G��`2ГYY�1�K�SBR�P���xt_Qs����P���� 1�Ԏi�=B+����x'���
��#�1�]u9��b�mB�s�$m���@m��'OΧ5Tv����NH茏�$�s��Q<}�Jk Fh����L�u�2��1\MD?'���m>$�2P��<sr'yy��϶Q��4�@S` �*�"�s���'��3�)�M���Qvt���r3��K�ݵ~�I���m�,��cH���㴭����{�D"�B5�l��)2qqq���7 ��D�@|R�V�]�l>;ҥ��W�*4B������J�B��R�v1I �j�ʌ0����H��%˭ꦬ&GE�$�#����c0+�<��%+}�w}��{|e���T#�Eu���������⎺����I	X�?
�	�����5]�'��0��y889��O�i*( ��Ў�	�5�kIꝌ�+C:�Lʹ�z�e�ڟ��@@� �XP\��)�A���T���Mh��l�� e P<����#0�?m)�(,Wn��0s"��̍<���l9�BT���p;��A�&SR�y�f2����������u���!��S�"�\"Q<3��,���A'��:б�o����M�(7ZМ�6�цdp�L@��Nar�9���BR�I$��xG��1��,��i�^7 vy@:R8h�7s �:Wr����cE��y�e�>q�y��S.��5�;/+ �OĹ���j���a�n;�]�����qfgh�v�� @�%d�Aѹ	���$��E�]<I�����'oe&2�^�d�=I��T��x�g���Hs�pQ�该21��xV�i6f�E�����ˍD��"a=���Ǡ-�*uo��BG�,1�_PP���~󚠄N���!"B�Fjr��N�|���Pt0p7�u+�$E^Aa5`)�]P;�aeb�RS���u^�}Ro&�i���EBi����s�+8X��+B�l9��:�:�'OI$����J%8SZ&	E5۹�?ाLBL(�e��i8��#c� 0|�4�[��� ��
����n[�-�ߣ�0�@��Q���R�*�ng2�i ��=�|�_ ����1A_Q�O�'�,-M0\�������ݻA�Y����M��D����쎕���&��清���/��F+���L��N�N�Nk�,--����G}í��O�4�=P��~�W����b����ک��z������9�&}}�����ޢ��;���;F��23�{�XR�fW�ׄf$xN�:��ȶ�ZO�	�#\��5�5�Zx�$�F��Z�Ύ&E�\8��/�ٔD ��ڀP֍��XP�����^��B�-�>u����A:��ҁe��I����EnG�b7���HH����h���G���roNLL|���r�`������_��i�SQ��K��u�{�,�<�LN��&��&��=�O�@��>^��3~Ƞ����quD�z���ji���O�y~�hr���;��&Xao�篵��C:*�u�}��$a��<���/_���y!�6QX����ud�&m��REEE���M����?7M }w0O8��,���mx�>d��a��W��;
��O����jۣ�XC������8��sF�u���Z\'��E�4қm�9IF�Տ�@3I�o�G�����#-3^y�GQew�p,?�$)�\�?�R��f.��F��J�:L� �_d�7\�ag��|��u�C��l �<�a��k���ƺ������5�6�ު�ݱ'J�.���U���?�AxC� t��m?mrǋ�u����(˓�^gl5UIA�mf���	�?b�)��`g&{��t,����1*�
ᎎ�! 2��I�Ɩ��&�l�̤�V�v�!b��l1�+K�2�<����6�0ةP�8��l>6��>4$/.!��h���r���9�"ch��a>L�`X�񾊢t�gq���4�l�ι��Nͅ�	�YK��h�V,oHC�pe1�v�C�ձ�m��A�w�����o�\��ݛ%<Q���5Ђ��/��-E�K�x����CԧMJ� ݵ�ӫ5w�W��,:��>o]xw_��"���މY�V�s�BS6�$oe�w����{=�'�n^z���\`��T��O������K\a>$���K����S�6�*�yVI�w�����z;�	��[���I��_�w�o��_�^���;+.��m��χ��R{��@�%��!���=<��7�@�%��&�D�'�Hֶ�6�F�M^��u����:��c��&�/?�ٶ�f�N��p(؆����<�p��M?��]]j��}Pr��dYQ�|]�L��3|9r9��>p�0�A��7X�]���o�y���V�q�+%��ٽPr,��!m��v-�;�+[y��~��}}�K�1���hyz��H�8^[#dd������@�ٻS��9�`��;��Xx��K�hn#��_�� �;��ut����g@���ŗ/�o����n���o������?yA�)�
`%<�j5kk^�١9㣹�-�ʧ�o�����@�������y��e:_�(S���H�O6>�9���Q�{�o
�l|Qt�n`�����0����7��pk��n߫5
��}�a���l J�������,d�8H�����AQ�V6Bz�������p�͍�]B
��y�������̳�� �̹G��_��S���>�_� �D�η����T����I\�u��
�S<^9���|�`:ߏ���D<�}{��.��W�����t���n�Z��l����*`xy���!6�_�:����.GȼxiΦX�6P�&D��� �� �V>쇜ݬ�y���0ʻ�kUa�p� �R��v�ڐ׺�K���E�������${������zo��m�|N^����9�	�9%�����d����ޡ8b�f(�[��{>�<���90������r��i%������_�q"��}1Du���'�]yf�[�K ��;ͣ���8�2�]f����jcF�c>���������m���"����W�8�Ւy�ڈ8�=�5� ��Ȃ�)J���_L��y�N�l�S�۵�l�w��+��ϠA��Cbu�^&@�':���qq>�G��?jȤ�W,){]6�4��Y� *��V��&N����J�q��:=��?���'�x[DӏM�z��������Sޔ�{H]}j��"��_�DxG�O��7W}���I�Mkxt��Z���ew7�a��eu�M�dRݟ[k���H�o��}V>e֡��#��>6�>���ҩ�oӾ�<=�b�J$�M�K�\�Z���?�-z�]a��I�(�y37��{ץT�d�����W�/y3�
s%N�4b����t��<t�|�v]
�����F���TxA*������'X�=x�ܛ,�k�ª�yi+��$����a�û@1_AVm�~ H`�O��N�C]����G@���+@��%ށ�>AX���ޯ��OQ 9�Lɲr0�ｚM�_j\>S�k��9�|�h�I�d�����C.Z��2����]�{���E;��}�e\��L��x�!�BGy�h��s�T�'/7C*�G��Nyx��ٞ5 !�/��|Z�Ma�B����ޏ|�anT�2k��	`��_kƹOk6���n��G�V�/��7��b�~Ee�E����BC�WD�����^�ֲ�����6��{���5�������ξ��(��ln��	�D�1�)t�Kl;i�� �n���#`�Y�dz��?g�����
�
c�ྔ�/�0��/;�?�$��l	۟������ѱ��F��:�WF��6O='�k
l7��>�d h�ꗐڕ}��_l��f�����>���F�<�����u���S)�ˤ�ӝ��!��Dj
PsC醹��x��E���A�;�8�v�%�JA�d��R��
�9zy��ҳ�]���s6�������r�B�~�<�q�~����O�QV��7��9��&@���%g*����kW��]���4.��a�`N|�;�H����~��$���?�R��ħܠ��k���̗��ؿ�� �`!�,���aF.�ka@�#������O�#> f��Z�|E)�t0�%��o��k5�8��y|(�{�<��I@�w
�-X�wun�������X�c3�e�[�~��蚮��� �u�����`�ξI�d6�?)楝����@kp�Rz��Z9��a���p�n=���u�m�I�<��|J�<�fėg_��{��F���&h�=�hp�L�.�6i1�d�%$�X��_8���k^,��ټ��4wp��#�D�R�~#ZkK_Sӯ�T�!jx�@��x���N�n�j���7���OF%Y��ɛ}�����n��Y�I�z��/;tm~����ͳ��̻��:=�҅�j�oI�� J�L;$7Bc�$�"9� ����ePF���������/�i/K��x��}��ॷ��yn�,t�H�BEb��%^d�m+Ux�6�$��>Il�>㳑�`d�ʁ���Ep˩���v������`Lm�Mf�P��p�|_�/ ���\ܓ��a��jcjƼ�!tK:�,vh^Ŷ�f��E��렬-<�yp⣐m��˙�C�3ߟ��yK��лe��������c��릿Y�=@)�;����E��N��'��^��h�)�g�~#�Ʉ�yG����u�0�^i�؃���ޟ��y�zA�YS�����S!�ao�M��"g�`���P��= ��2?��o�f�f'[�m_!/a�T!>�@�Ύ�y���d�O!���yq��Tw;�W�Z�my���������%�E�ƍ��;V���^�I[^_�{��7�"�4?��K���͇5��W1.]�[�x����0�##F� <{������i[>�v2��G�8�jp%����+��L����?� ��\�>���W%owT�j���/���[x@��h��(�X��J���|^�_�P��%g���(���3��?����"��`^��~��:�� x��ڌ�}�}��ʁ�+x���A����ὭÈD��b�4�[�<��e_l��ح��^u�oc�a,�3�u�N����	�$~�XO����!/ю!��
��x_,P��.����Vrb]+&u��)�Iv�/�\���E����rd�A�L����ѕo�w}�3=Q�44���dU��F�
�8/b-��$�<��p��[�����d�=������9��^�� �n�)�R��(�Aޤ)A.o�8`v��|q�fq��{[�D���$F������Xc��O���e��߁�F-(�G}-(��	�-���hM�{]�����Q���F��4@G)�2��*?�(,��ur��Ҁq��h^�&����+~wk48uރB��{�|x5
�0�6D�݀<�Z���){�oY��DW4����6p�{z�^�y"������*EVkw��/Qhƥ9\H���xx5ۅz�.���3L��r�ǝ���1
��n	����:�n�Z])��������<��X��Xq���!͉I/����R]�mGA۠�1�j�^�	#=e��Ս���>�I��8e鰵�b����L�2���<����R��dHJ�.�^�Kʐ�/D�e��8V��x�8�j<��{q�����<�/�E��T��I}�A?���YE}���G&�ߴ".�DW1��4+�dm�>��+��ÚJ�}csm�ሂ2�� ����r���$�"�� (�
���Ƞ�AeN2�`��9B�H		����>�{�}�{�����^��?ػ���Uk�֯*U��!�K�|�>���u�O|����^������Z��OE�8&-q�g����`�$/��UJj�L��I��X���/r��
�3�Cف�[ �6�m�F�.J�(P*�;�Y��h�R5�W�\">p"���-�0MEɜ"������K��݊����R�1����&��S[s�#w�GB��w�z��p�߶�ZYZ(y��q�q�8�eu��9Y`1�w����p2Q��`C#""���1����o�#>ǳ�D��Rֳ�9l���r;�*P9� q:4�i˥L������5%��@![�}9�&����Xÿ���}Lx����<Hv�)_N���6N�7�(��^ڑM�.ܵ��뉫dĤ��ޏ���q�<9���=��)��Q��&��K*�|#�i�S�c����%����_�R��9�k��M���Y���礪�+L�� D��7��+ֱx�s���%�������	�m	7Ʈ�~@^����D�$!����0��7%�3*"܌�����Y� .�a����~E�M��`^L�G7�� ���)ϛ&(��t��|{�1�#[�,�6��4e�����z*���lI�����V֚�=��V��
�Z���K@E�u	X@�oR�&[Q7�(�V���+u�P�5�<]�����J��=�Z}턆5d������9r6����b{t�AM_;�߿��i��V�Ujxyɸ�S������ֻ������w����>�I�AG�����;l���$��`�)0b�ʘ��ϗ�T�M��2T���@��W�p���D�]T'�'�T�}����M]V�|�*L�^oj��$�Q��=��7�U�1�r�=���!�����ʈ�2��[����I�'Na���-��Ũ���٤xg�z�����g��U�7o>��Rf��j�Eǃֶ�k�y�'E���`���/_'R$��f�A8(XhX�L��Vg[� ]��%/�Lꥬ̮�T��7x禍�i�/��b��~U}���0p�&'~����q�Ĥ$�TI����@�c �c���P�_*��3���B��*vtx��X�WK����b��a�j]z�������vk�u�2��yy�k�I[ 9ΧW0�`1G{=巽�o�K�.��Z-j��U��`*�`�*ʠ�ƛ�yܰ:i %����L���]:�%�ɐ��J?
S�E	��f����,�l��M�'��7e�Ol���>m���)l������N�eׯ�N��W�Lкk�ޜ�?}�����4��Ջ����tf��!5~Csssg�����2����@p��7o�H�D*�n����B����|�1��=�o5�I�M����%���QdT�ߺ�`$��볘��$)�> �׺�q�+K֋�L���*L�ș�Q���,�[a�p?zt�Mxa�J_���6�`��m:�P���"�A���Q���{�/��L�J~�?pa��5�s?�A-���G�'MB�`��(�r���`=�C�%�I��~�q}���I��58�����In���
��I�=��c�2�;66V;C:�箏~�FV	��E��*/\�/�h�(!����	��N���( ��R�^h8m�V�Zu5ֻ���?����=Xuwa��z}o���q����ʻ3�X	�FN6�N�q�n��(����3��*��'G))'??M��7ٞ�:b�J��������\�n�u��Q�Ԕ$K����+�-/�RR����sM�� t)m�`շ�r��įC;�S����K�%�g�'=�OYs*P�U�o�Ye�n�cw��s*	@kq������G
��V�I�A�k�wDM��%��0�B�ׄu۶��:���!�#:��J�_���>Nqʦ�I\�'>H^���#�7&���t{�>����c,���MMMSA����=����f��x�Q�%����P�Z��2B%��e����6#�l�hnz�p]:p�����s�-^'�%�g̸|e�v�R&�`�t����z�� 6 �o>�Z�����ܻ _I]�5�z~q	>�C"߮l(}F��v��{%�M>Y���= �W^�t~r )^%7�֑/	�}����m��b08{�=��>������Ѫ)�:8���*�D��Dݵ:	��'���_�I�|q�̊i��q�1��$Z���� %�D���5���lRMpP�	Z�_�	
{�}gǴD4�l1�=�3�(U`��OB����S�,e�4�T��	�jev�y�����O~|���(��c�5��.�S���#p2<�s1�[�!ǎ���D�� ��~�[�!sC?K���Џ1��Y����2�E1�PU�����`" -#�]?���a��G�ېW�� E���7�_����L�� )FE�m���V�޸�)��X�:EC,�߃-���ץA'���8�4F2*Q(˴|�?��#�M4�x��|Q&zௌ�P�N�Q��~����ba--n�ys'��*}	�|��ězg����vY	�(�@'�1���eC�����8/�j .�q9�������ݤ�AIh�(��(WG0杳�Z�A�g/����.�d	�$��1�.��ԡz��@�s2�`ʳ/*�5���V;fQ~�:Z�"��{����kP�� V�ea��a�ꞿ�̿����~����Q#ӡ��򺓐b)p`�`�P�fЂl8�ֱCPV9G(���hM�eX�[@T�G8ȫB/�A�Yd���}������o4fL���4&Y�f47x�ɑb���H��A|��(˳�f���{����luEb��(�b��*�ΏP��
��=CN,����+���b��RF�+ �d�I�i�r��q1�x�4gQog���{��S�l�'�;��8<,&.}��4P&�S�.w������I�X'��ʼt�-?
Y�ܯa�?���^.b�F`b�;qaf �o=
)�x�a	j�`��� ���5�����_�	�3���u�2��SR���L������/KY�����ԪP�\�P\D[�@�{���;?�׈l��������W �zc� �جm��2�kGA�g�wy~tkG�ڭ�G�[�Y���.q�r��zv�a�:��-�:J^����On��{��n��8u�Q�a�����L�����%��V5��ѡ��/v�Y^��"hSa�Y�#�x�e�g��D.K��/�����	��Ē(Ŭ��&�Θp�s�/JpM���Ж�^�ho���R�sGǑ'�!�A�����#�=J�����c�OR}e����+��ݹ��F#Z��%g�����wkoƄ7ekdtU��q�2�*����9qC���N�M��@0u����ʯs����JY���=�B}[w���??w$ԧ?�S�iA���y;�0�����bL}�>��+K�>󄹹��%��O��<0�Z��)��~�#���dۚ��V`��R{�����jT�za>��n���l�n�-��Ź��=t��[ny���|j!�?\g�v9u���ߤ�z��V�\h��%�ۻ�љ����i_)n���^��]˧��۝���l7 ��}"_��t��7�]����mK�8P��60'S �eೲ<و�#��(!��3��u]�Yn�l�v;��U�S�"q�N�[���NKd�(P:ҥ�����n�{�\���>B�����۟5�Bޤ�+��E!������'[����y�e�O͕�,M�;Yj�GFa�vlp�U\t�(S_0�r�.r�b/\_�\i5�ф�§ϫ�''a�~x�;�E�͠���龧gTc��t����с�n��B��2���oܫy&m���#���4����z�y�W�����s�����x�@���<x��R��y��CJ�	��s^�h,��P�%���sQ[���&��G�ܡL�*tV��ǫ���ݚ�:d`�~���ߒ��d�6l�Y��L%<��������v>^��������|�~�ͱ	xw_�����D�IYz0����X�=ٷgg+)�{M�P�)�qL��A{���Dn�*���=/�caFH��J��~Xٴ�����ħ#�"~ﮪƾ�%%j��[�@'`�^����D2^��d[c��@Ѽf�e��SS�������`�n)�:&�[͹������XI��҃���vS�^�g�� BH�����j]�Ε�N�N�c~t��^E�R(O]�^�΋��G���,7@�t7��1�"��}Q�j��z����5�Qx��$��Tp�K^ań��J0��_�'ʑ~�A�j�8N�F�z�d��e�G�y�ȧ����HǌS*OZ�;�W\������"�vnTۥ�f1������=�� ܋��c�V��S�(-�2Y1�%a�/Mt���jl�JĘ?�|���J
S�e\3y�Q�,�TQ��K���@jq�=�����]��&v䒾����鞯�������8v}��P�[U�ߣ(�=">k��f�߂Ѫ2�͝����N������ݮrB`�/1Һϝ`��w���	�(K��5���h!����β�X�D�5φ#�푫�r�3Γ����>S��"
�P����`�n�[XJ�d�ݍ�Q�+�	>�8NF9�|��H�qMۅBX�:?�D����%U�V����V�Ǖ��T���Ow.��x�\�����-o"��ӎ��Np�"��h�/�mz�a�+��Ƙy�f9	��o0WR����c0�	BwV�$�]���V�*��m�=��~���|s�j�/aV���+�h�͂�R�w���w"���,�|�Z*�c������\K����Fy��yZ@1����]6GU)ڨ�!-�#�Մ/"��������?�����ZU�ܞk�P�?�hmח%�TN���7��1J��/,,��'⸾�KK{�!�/�vZb�����5s�@�W� �������C������g��w}�ϝ?O���IY��J�����/�,?wH�ym����{B��#�[δ�d��kM3�gΕ+W��xw}~��d�G())��\5��֋pL���p*;��9��Ɯ�,�7�Y���&C�lt��p���s]�X/��H�rS.�a����%���$	���@uD��T|5����gn��OC�׎U�jp�Oݭ�΂;D"����%zy��6���z}'���"l0�n�^���|L��	��o���R�܉΂�߱E�-�}�l��3G$�;�w{�݀��c[��K��b���ӥr���p��Oa%u����'{RRR�	�$��mwf�B��<�P���Ca�����au
���Ȑ�A�ڋ�i|f�P�ѵ�Ę����|����H��T@��E�{��jk;̽��E�D/R��H�b�xOk�w�|81ϋZD�Aj�� ѣ=7\_O�L�=�'�)l<?�wTC\N�:r�1��7�`{��ɓ'�[�����E���f��3�-[���bC�k�����	&�(�|ľ�3��O�$IzQZJ�@�-��Oii���!D$��W�G�����a��偺:RC����OpZ	 7�ؠ��H�Ș�؊O�=�~���	��(���"�j
�=m��|���+�
�϶�M"��	߁�d��$	)f��������S�q���i\�~��-�`�r��y��ڍ����].L���r�(k{{�&X;�#��`��-u�0r�X0(�N��������e�P�(����lœuTu��oAh�R�����f]z�L���$� ZG���U#�kݽ��=>=�l�5�L���f��/���D566�h��ބ�g"Q���=����ݣ��ޚ�����EN���jp�77���J���`�+a�@�m�3�������G���Eq���d5k��UH�<H��s�v6��|�S�-s�w�ퟥ:Gͮq�дLX+ru<^�#m|��s�	��75&*��;��[�=�o�kD�����ve�$�]ײ f���9�6)�U�^��e��U����Il�>������t$]ۣ3�bb%�Z"k&�?�2�����g��X*A7�	'D9��

bY_���)Y���%�� Yx_A|!��;�� !GwSJ����������D�Ae�e��@
�:9C?�)�ޖ��������.]�e�p�,,,h���َ�@��Q�h[*p>7����-�b{�g���Ucŉ�/kdtv��1���a(*��PfFZu�R}���A�d闓����U���!�=ؙ��E���v��3��a��q�0#�Y����?�$	v���g7h�ٓ�D�5|>_` ��d1&'��}m����H$R���Ç �|��
''';�-�7��F�^��K�Iutuu�2��L]`l�O����eH���G���ˋVy�zb����W���k
��O���Tuh�k��i����]y1r��g�s�E�JIH���)��?�jS5�Z%��M�g�52$��;�o�E*4�����Rw�rLLL� 4Wfz;::bhA�,�1Mob^��[����?�ژ�pSo	*zC(�Z�kq����@=Ka�ь4=�2�R�ޗۊ�o��	
rd��ױx
�z�9⼟*R+�Zx)q���o���}���I���PK   �<�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   k?�X��$W� >� /   images/a253aba3-74e0-4776-8a4f-66dded74c7a7.png�USL��{��Ipww��q׍���	����]�����]���9�T}]��gf�u�Z�J���! A@@|��W�����_ ����X���߁� ���:���L�C%�����Qs�:3;��^�fkjNkr����!~C�L���#����"�o����8G���#2��0g�\�.j(C�ZxT_����w5��}�U���z~�p��-nn������������g��H"y�?�L5�� ��O���:fQ��=3B4�c�`�"l��B)������A�r��w���#�?��#�?��#��Q������
<��N(w� I�r��WT]�ܳ�h��=v�4������
�� �FM(b��5ӎ�Z��:a{�9Z4���8��Y��O�7�xY#S�HC'Tu�h�����)8ݿ:��C~��r�K��4��u��B�w�m����V��B����y}��gG�{�R
���f��O�<2�����{N�i�����T$O��D��Z� ���������<���:� 1� u.�=�w*�k�*��u����	}�Pm�\=֒Fk��3��$��z�]E��u��%�*�ųG�X��b�y!����L�� �����$�.mf~���-2f~�o��%���_:�BW�!��	%Q��En�&�]p����zy_�L��/m�����J������tl,{a�2՘A��z�jx<���|�z�N�]4���mZ���s4b����%��LJ�]Z���֗K�1�/\a�K¦U�A���Ѷ��:�]U��k�����dv����G���b�G��ޢ^(� �2]9ݭ���Z�Go-�;,�$�O�������됛���� �ڤ��	�:�e$g]>���?��rL�(C�;3:�	utm��qO�:+��D]���J���ls��CȲ����3���Q����%/������n�=���V���S��f��4�֫�j��x�4m�NK`�]���m����6��0�m,��c���=�������ڝ�Q�(?{���T2���E�U�2:��$L��B%��V�4L���}w���O����>�Z�Tf+u�Ŋ?cUK��"9�����;Ñ�e�o(�$��-�ΟA��d5�	��&cS�dao�4+�{h�9�c��9&:]��Q64m=5,�`?D_}1�t�a��Hg^��h��;9�H!W����&����;($�j�Y	�^�v�v��1�=��fib��[.�aHy�)-��Fm�8
�P�y�q����X��N��A7Mh,���S��������������w� �&i�4�f�O�G��~���<EV��9/���	xo|�W�=���s{S��o�e�a��Ӌ��im�����J�=«5$�ԜJol}�������\~Ȭ?�8�E�R�G���iψrZiF� IG���+~���h;��i�^P�օ�5p�L������gZ�Q�����T�+�.�+]AY��|�4j�����MB�DƘ �Z��0���5���F�t��)�H�-�=Ty��jD��a.����C?�]�x�Tx� �	����;R�}Y�<2�1�!q�\�+�~� ���A�?��L��e�l�:�k���ǂr�7����h͑L&I:X�~lOzUug�]5b��Ɂ|Sl��ʃ
�=����worn�q��h)�s��o<��\2Y.',���	ٌ ��~t��#�jg.[�b�Y�/J~�OǙd��~��g��H��¥g�.z�:\1L.�׻��s��~ȳ��)�칁������ۓ���]��ߖ��F+�û+���/�V�n�����bLl�ubW������ ��0i��f��c���,. 5��tU�x�@)�T���v�i�R���t�c���!��{]�,�:2�|�
�I�MKn����09�w��7;���O�/��.�RQ'�Y���%��gF��d��_��k=wi��F��i�)�g�l�KQǅ��\&�l���������Sʠ��y��zYjF"�l�JQF������T�TБƠ�~���h��O?$8�ѷz����a��PUJb�������}1�me�4xfw�S����^��m| ���kW��S��s��s�l ����W)�7�8➪ۢ��έ�[�; ��!h��}�>�7^��[�=��P�b�M4�m�	�G����M��M���@��~�bZ�&3ڬ5I��u��q������N��]�,ڃ��X3 ��9��:�ܳR�9b����G�$�\�#K"e�ÕI͈��f�/X�2������\Î�l���ޕ��Bt�����n�¥z'��� ��~#�YC���1�	�L#A���ݻ���|�KK,�D�[Da���V�����
��M�j��Z��(D?�DDKZ���E����D��!�9ʚ7��'��=16�V�Y3������������J�� �G.B$B&1���j.'�رm^S�4�x��ھ��-֖o���=����"AusPNؿ^�$�Nϒʁ����f OW�
ǐo���8h+y,�wѤ�'z )ކ�?"����b�!��;FS��d;?��1V���9M���?�}���;c��(�xը�Bj#hA�K�iJ<<���`�k�J��=����N$��! �iE�R�@���R:eO�&c\uF\�T�=�@�_�k�Rbo�N�Zõ��	y�_o37�7Y�� �D����ew��_as�6L��uE"1�2�����1����ս��Ș���+m8̹��&��]i��e�4���G,v� �K."�P�ȟ������c7�9!���<p8��$��&Ձ���Gl�[�l2	�?��+Ual�LW������q�\����?�;�J�YS(o����S��m��r�uI��ʰy����Zְk̦|r�?�f���BE���/�ƛh���/��޵��Ӝ�5s3��y�m?|�;���/o���o-ܰ�E)���:fbUj����
VK�,݌J	����FPٰ��^�.]�<�2��Ж��wa*��� �<����K��EZ��#.S�uR�n][�T�I�%'gg��0cH!����|4����0zNw�ې���N�� %2�k��k2�

��9F��A����I�>��N�|CbH�cф�^���i��ˇ%u��o�:�7�L
@
�	��G	z8��
�@�l���'��l��^��Q넠��L]�^��u�	Hۖ�dDQ�MKY�^ต=� �����$�^���|T�Q�0���9i�C�I['C��l�l�#S�_)/A|�snx���<������=G�q��\���B�z� a�,���'Q���2������D�ƙ�}\ô�������)��YJ?�5���Y�"E�E�(OOO0�'�#?0V4�!Pb�_I)4������>����A?�y�&�b�6���@6ᰉ܇@���m�����Ai�Zy��N_A,?,ϡ�g]��H��?Ux��c2�&pro����#W:��y��Ij�ʵ���y���N
�âD����`1`��+��#k���6���Y02C��u����׶�z�ԯ4��ڙL���/�����/%c�Ǵ��x&���"SL���/�Yr���~�3Q1�0�9�B�~()�+.��%$g�l6}�4��:ZG��+�����1��'�ݥC�	(N+�9�m2%G��t�;�n-uʒ��� ���z�j����z��s�����6��]P�YTd��4�>oϹ{���-�;1]�I���H��y�"ܥ��{s�)p.А����ٗ��}rzo��y�7E	 ����]�!���z�8���*�*��������g�.�	eI�j�W�a��2��߂�ըe��;R-��@-�f$���-��YEAJ�(��N�c��++�����.�l�,
�V��7[�MH�C��+K_�}��O�B�A��H��`��G�'I����		��鍖5"v���J�x{K�_&7�g��>�1RFg�)ߔC�!�;�s����2���l��U�0`;���ԅ���(V2���U�-��C�%M�G�M����*=y&���\Ҭw��"���e7|��r^u��kNY9)�b�Eb�.!��Hڊd��v�Ҹ�'��c[���Q�Rv4���%p|;q�
G_�B5,{�M�����QN0����T�T8ұ���_ɔQ ���j8���=\��h���\�U�$?��w튡Z��Ϊ[a�Pw�:�!s�UQ�{F�	;��3)��t@�j㣦�H��d�����7����҃��xo�� ���4?����d|E��y8q�aec���Q�8���#8`���<p�u�7�?]�
FN��x�T
����2��j�nK�P��1e��&�k��:Qֿhޏ!���J�_�%V7�ҩ� ���GjU+8]�"ް^�v�2u�6��:� ��/�b��i%Rs�r}U�f�9EK��oW�1�F�d%��]��JsGf��:�t��N�?9��͙-k~�$7myb�à���
�%��:��s,]����ܬ��SG�2xo�W�n�ا�r:f�_����E�~>@u��@�ы{2]�>��*�YJ�2��#���!�E�F��(F`39d��7��+��n�[�L����@��K))�% Ob�A��ҡ� ?���/��� k�%}.T��!}�:T#bz2� $��j�i|�o���m}N�r���y���)
)9p�A��SMU��Y�Z���e�H���o�
�s���4��B��Q�k��Y��щ�g�6�C��	�@꧖<�5E��5��$!�:�+Vm�O�B��lx����Ɠ`�̟L��tA�S7�O��n�c��?����d3�tY����V!���m(K-�!C�Ei��C��*t�21oa�;].Vp�T@B��:����S��&{jPЯo�S�_$5|<�����JV�޻�:�eG^I���(��l���!�)<���g�<�ŃX�K��o�D
T#�$��f|rFѿJ�������WW�Ph��È���@�*ys!cG���OxH��`�Obb#A���5%��ތ�~���d���x����_��;���Y��W��ע���,U�jgj}��6[��_�cӌ⽝��ؑu�B>�x���Z��A@+��
�P��;}��@�}^�e|m��"��_X���Ҡ!����y_�X�_}L�K�`ZA
�Y��i7�H�y��[��O�YtC���z���SC������ff����-���^S?���i��^��n	�Vs�LQo��ý�ڏ��H�&3�C�JI�t�k|��ȿ��i�
������*�>1��^�Eu�%ԭ�oHO���jJ����/�I�tr�R�s�(E=�l���<��";z�;V~Q��~��tL����-�r'��ܯp7H��$Rqr#�ª� f��w��Q$�cN"X'����O��k��`M�=%���_�:���/�(�hTx�Ѧv?�4�O�`�,ꨟ��YΛy��j�p5�E7�����Cw+���A��"!9F4̨|���y��ܣ��`����F���q)m	)Q���Yb'd/���\���9�sj���5��:ZU�B�~4z�M$?��ᴚ�R��/"|�ft1nҏ�i��&C�<���ۊ���"
�����b@��0�?ٺï0[==�����!V��(��\����ڡ	k�����MM���e�.����c1��7v�ʯ�(/	��$R5����N&�L���L@3v�p�WI�����T�,o\��!����29��[:Y��WqΪ����[�L�En0�Ag�Sy֨�]�����M<=��KyLe�I��H_�DJ�ԑ��0y- C�v���p�i�I𭬪�%5V$Yo�[��2ɦy�����?�I�T��p
~�G�n�)yP��7��D���Mb��LH��;��y#�ޟI� %�o�u�/���� |a|�QgE�LcC��jU���Q��X�o��D��,����-�g1i��x$2�B(a^p����n��N�@��i��Ο��-�e��y#�sd�O���L��H���h*�gߛ�i��Q.�p`y5t��vn�T?��0m�_7P�姢�-�r����G��,O���ܸ�h;��|���]ḯ`m�T����CNw���}�`��>O`�Xe��򑯒=ħFI�]/`;����l�y�{?� �����%!|��n���yIۣ��[�a.&CFO֌�%�#�H�V�P��p��R��m�`���>���H���f��������A�>�������C��5�3p�g몍^���W��7��o��Iu�?����{"�XJi!�'J
?S<=d�A�D�8�R�``�m�ǃ'�~[�q�p�\�n�"z�%����%66�!�Y_����BL��Aow�F��N
@c"�X��V'�A�J�Sz���G�6�Q��zqy�sIP"a�e�+	�v����Eq����Qo���noƄ�fxz\���~.�W�k�a�;|�x8�%-Q0W.e
u%ȕ;�\!��3c)�͜�����ZuW��Ue��=h�=Ts*mfMB�o�g��]�+����h�*X�E%�k�5HF$LN\�L#��(*���j\���?�pJ�O�i���lCo��o��ۻA�#���a����b���DR�B��y�#ф/&�L�T�W`Rnͬ���q����▄+�p{4hc}NC,��tN'6:�a|��D��hA1m�V�2e��"��9
��˗�ePכo\�G�$5�"��"q��`<k�z�-�-]n*���-oȬ���|����V��b�.����.�XT~��t�x�nY��I�c�.����/����-�W����V4�rt1cV�>ǋ�M	�T�!��)Ǖre�L�Irh(��@/��n6�g��^�u2Ut%q�I�Pp ��
yǴ���+�g}�1��{����{�g�(;Q�(Eq�#?���gY��p��DC9�C_�R�?��5�@ho��FtoHN۸�S���$�����c��9�[7C	��z�ֈj�����0-�:r'���guڡ�B�u1�I����H�-�ְS�_;�M-Yv�[C�V3�`M탅���yz}���@@�/��3�����f��{h�h��Ә�V��rS���^(�(�k�:�m�����,�+��	�*W���dt���(�X������f}M����}5]�_F�D������)'lIF���I�?����82����Y�i%}�J�\�q���I_ĝ���K*eL�̑!⊻���>9�§�)NSz{�U�	�g���	Qm�0ŵ�Ƃ[�/9�F����0���H��]E�
M7�t��c�;sdJ"����%lTb��+D�>^��	����Qk��V��׎�Yg�)T�9�L\�O0r���ڨz�p���5��C�"%[�V�
�ܷ
5졭����Ԟg+
ʨP &E����;�aq����g���ֻ:O�w#�|S����+_��.R���jW�� Qgֲe�B�P�:���|���q�T�C���KIц=������ͫ�n�n��snFy���Y,ٹ�F>�S4J����P۰d]�_�@?����6:i�M畓�ⵉa��m{�6UӶ�����@U^��#�$�
���;8ւ:��.�j�t���2��tޣ9yNg����I�c�ײGꆝ�N��PV�ajbO<�.�f���jSl��ͫŮ%�Y:Rb �n� ��o=�Y�*��	��9�����
�$�#����I��L��2�r*��0+��/����
p��9��mkU���-�&��Vj%K����,6��pteZ�����	f�`��2�=a^bw��A`N�-�YXZc�ăԭ%hT��F\J�\H�Of:���z��L�����h��rݽ���~~V���q��o����Vd6%�>���Y�
J�%MHd�-W+]Mp��r���l�*�J��Z�)Vw����x�C3��>d��1-��%K��jYčTLz
�o�@B�]���xC;�W=��@���f��[��O83�ר�.�B�p*"a�FL�O�EȰ5}��ui�e��K��=F�Af��LB"R7�����/j�����9�oRb�*˲0�1�)��e-n�g�S`��k���u0e!�z��ϛWC�h:KN�Ή������刾U7����m��X�+�����No�k��jy���wԼ�El2E��?�'zn�>��[|]������1u?��u31�<�t���1l`r���ӧw�C���Ũ���}�Β
�zY�~�l� �Ç=O=�]���*x����[D�e]O�/�|+�z��fΞ8Cd�l)�ei�Z4�|*1fҗ�eà	�%L�K*;�y0� a[9�-Sig�O�������/�mv"�������,�"�S����|�i�*��wG����[�" ��mŭ^�l���ֺ����f�����۩A��{j	+px���@�@9���#s�0���G �y3�|j�ũ���]K7�#�0����#��N��~}�)_����ʿ�WQ�Ds��Xvz��ʍL7MZR��Lz�|v�Z�S�nP�ojBVpL[nɁk8$e�@'��H����cט��"v��ރE�ȯ�M/6�4D-����ܙ������)I$b��A�3��V7��\?Ⱦ�XR�����I��p����?M1��?��Qk��cE0���J?�>*�X��6���<%��]\��6��'�&�%�UJ,:�f�:��h1^�fʸ��:�aR&�t"��e�]�3�CaU��F�s ����c�44b�72*���pnn�jk;i�P&ze�Ex(q`5R��V�>HaB��<B�;��2��P�?ԋ�[�U:�w��ם�+݌�<=���8�M'[ˑm�:,0�}�H�&�к����ٺ�F�{yA�,ge͌1�*ΐ�+�-���G63qK��Ao�+�E0	�Q�\�9Vf�"e�K�����I�hH�&���S��Ū��*ok?z�
<?4��� 5SX�S�Ȕ�����}M����$z�<�B��������ά8��UFy��b8�WcwtC�T@�ʫY��t�q��tkc-k�r����p�k��x'<������h���e>V�Oi��,A|u�#�8g=i0ۇ�r'���"t�� OG����� � �#6!�tǞ���6���qɝ']N!�L����I|C��F�w�{x+��1%���;jl�f~�����=��v��F���J�Ԛ̮��f�qNCG^�G+x�8��f��vgO���/E:7�ф����7g]�%���oYگG�8�R4�"븲�@����2(>��_��J�5Ya�3㠰N��^O[xl�WLh$�3��a~��
	��U�ɗ?��dQJ���U6>L���E��m�_��8..���bP�m�!?�_��O�#�8�/k���9�YT��S�C�����؉�S4G`W�R�>G$xiy:��B"�-Ǣ,ŝ���H3�0�2l��$�����ѡ��I�,7�bz�Q�Ob�!��,�93����"��S{��B�z���Fuay�w���u4E��(�a/XK�A�8��IG:�S>\#�O�Ϊ �.��(|b�W������
�����(*�U�Y�v-�n��r�����]W�oX]}���<�胈��S?X��,��P�����:��m��z��H��p�a���8�_�pF���+EK�}� �M�iFP��I��i�{��A�p7��~m�����Q#�;�T|��Ѽ���s'݄��8��&{3����Z����1H���[�Z��#U��ћq�F	�I]��H$i/�&�N�|���t��"[�䰑��ъ_�TC,$Ӵ��^f�I��Ծ�l�/���A�퐂�$`����4��4Ll��f�� �k. j:��4;��T�}]�
ߕ��G�e���ie��j��!��K�߸L/�h�we*E��*��,Ddf����U���.e�!	�ыR��<����i'�u4����~��j�9sۥ�΂�~pf����L\�-��8�Fc�^@���w�O���,{�DD���[Y����вb�]�V�egp�|���l*�\���ʌ�e]�
�W0�7�a���|���Q\;�R�&#�)�0�:a1�v�`Ԕh蝨��5+`�)8��$^� K.��+����'Y�7�掦���qRz�nCe����H���L��|��[�w�UK��\��N�̢"�e>`�c�`g4��G�?G��UլeE�vŐ��Gg�Qk�R0�$����iY�?I�ZN;�������8$���4�V(T�z��Z�_�R��'�C�1<Ye"�SmjX@��`!�0eNF�f�H���j�t�oY�^���as��)!�UV�� mI1�~��0>:��BzvQ�Gs�V����� �C��w*K-����fd@,5M.k���*��*ɴx$+P��AosE1o�����2��B�`�J/��
~����'����$�	^�Rl���%Ǐ^���i���e�������ԝ�7�}�g�!
�����tu�Wh�XS H5&����af��K��Ө�5��k"������tZe#<v昕N��Ɍ�Q�z>�Ӎ�(`��eτKqQ���;���-	.��֕XWo�ѕY��g�������JNi�Y��&����!s8dX�Ēu87Dp����q�7q��f_�Q�c�)#������ 1 Q�>��O�\u�ڜ܆+����O^c�V�$�,���߈�"��M�D�D���u+�Fa�6�1���A���������B)�8+��;����[�3j�
�\�ߕ�����;2�)nT�Z�HM�Թ�T�T��Jud!�ϋN�A�C3��_�y��C)��?����_�PjOP�Ե��<��[�ד���:
ӏ�2��;R�VB�E��E[�H���Y|�h�U�[�n]�4U��7�d���BQ+,5("ue��)=�ct�ٸ~�É���H�����aӹ��9��9��H~ڎM��8k#yC�eQΚ�������-������=j1����r_��{�3BZ�:�P٭H&�a��G %�w	����,Vm3���PZ��*ܮ'��%�ڿlu̧>H�죀�S<V��V�|��1&���Jݗ�I�(	����G���"#�U�00f�A�)�^1/��Te@�c�g�k�m�Ŀ��g���8{��P�p2�gx�4׫m��Jܔ��u�����/jܔ����.,�AF�*o��N..ycf�5r�M���p���=L����g�)!	޺
�������6���7z�:�_��JH�Z�1`�m텊Jb ���������SgZ������mb.��R���l���KCV�gf1[:��]:�gy��s��1 x+�p6�S�8���"7�����g%��F����4��R:vL�]��\�F1���K ],����|���̙hv�Nv_\�n���'�NϏ8ơQ~vZ�����5�@�B���K/v���v�bekD�٣l}#8�9���X�Y^#�>�����D�9��:�"��ǐr���B�m��n��c��])-� �"�\(O]���BA<�u\e����.3a�/'d�5�L�sKy�B�ģh�=4$�Vօ���	�$�<ip��nG����Usz���6���?6���E����-��L�"d#�.,i���v /�ɔ�o��*�լ,K�e2�N�TeЫ 1kB�%e�ʚ�#���H/'�`���2�n���DH�K^��kیdX��rr[}l��E�ECr�0=A>n�r�بtzږfPII�}X�v�~U�x��}i�Ғ3�,_r��g�|����[\�u᫑�z)���5����ȵ���y߰��#�Phj+Ƌ����G@�OW��^�uy�|E����Iۓnr΄�6��}9�>����:��N��/��++�;Nx���9��x�8$�,��+�������A1a��e�b�@ �ڙ�?T��#�E(o�H�l+b�n���|���t�� S�d�V�0��=4̣�r�r�Rfܡ+�@v�Շux긋��w������a�}��P�&d_�
9=�s�؈���35޺�ߵh��
��� 4+֌ݿel�z��."�y�����w��G�%�,?0VfqLڅ���էep�����pmy���y��9�z�D�1}�6V����
�kA<��VD�|JN�.#;ΕqƬueM������0x(Ӵ$��c���B�������qSu��?�2W��ॢ���'!�^����B��k�;���zۖŬ���U
s8F���Kh����c���/Kn=��N�#e�S{�%��{a=N,jG��]�`���\Y1��~T��.4�}'�T <]W����~B\t�3�1%�kԃ��1Z�l1]^��isu1N�+"-���q���} 24.�~��KE�X���8d�Ӭo	����fn��� �;��;z �+�P�kf>9:J��ɔI�
/fV�Q�7m���٘,�,3-�XlL�@��b�+���S�y7��1w�#�H����Ex��	���ƴZQ����saM���v)��ەɪ!�Yo/L �3W3T�3��dL[��p/�Ec��&s:��T�N�R��k�ҁ�P�PX��)��F��$Qs$�-H��~R�&�����3�Թ�N��F����J�g��M.��פ�[�hː�K����Zr`����YJp8�T���ʰz(�����XO�tcg�d�JD�9t2�ͽ���<u�`eq1��fKO�aV�^��1qT:�|R�i��ު���d9��Yaȑ3ۚX�-�<#%z0�t��#�(��h_���"���㯼cO��z�ߢ�	�C��f�d�gC�No��+�oNd����tt�B�qՊ���-	V�B+a�?J���%�HX�j�F�O�`%+�@	{J��R�D�k0�*�,�ax�ǈ�����GGIB�f��b�}��,�!����)ΎQ"^��Vp����zzFI��a�f�aT�`���w�A�H�H'"�X��j��/-y;��8q�(H�j]ت�F��t�@�eg;��	��n:���B�B��f�?<N&��{&:��;�g��ͨ�_��tq����ʡ�{:H�~�x��5�{uo�^��W5]ZE���2�/���;�?��p�J�݉�9�d{=��@n�mC�6a�g`�9Z����x��I��ß�Z$P�Y�Vt����KsN���A4�w9��am����tzx�yer��c!�7�m_��3�3���6L�I��T��k�:C'	�N���g��ہ���,·���%�f�̂��צ܃�g!�y�H+U�)�p~�)�Iw�=D�q����)��D��$W%��w����������4�`����	/5��e	W����H+#���E_�wf5����+�-f1�>ncI_O=P���F�����6��F��="!&��De�(��U{ca��u!{xȭ}!�x����Jvf�|M�B���{�J�5�{�[Yjw�E�F'B��eI6Gě���i���CS���b?r��z����p�
����|Rg�8��ː7�Ub�Ù�&tо��ǂ�i��S��H�v����(�7�-v�p)bn�m���x�56iѬd�Kh��$�9�P�N�~Hx\��섑��vݒ$u��V��R���X����k}�N�HK�v9Ѿ���8vG:�":���]���̴�J4n6�'*׍�\zF�R9!%�G\YGq9Q��Zt��:����v`]�Au5:�#�ԇ��G�F���ܨ��ǯ���k�M#�j_t�d��k�2n�C8Z�2��qr�`�l�e���Kq���<��ĴT��{O59�m\�����;�$f뭴9�=���Y${�O��F �����x6�6��F7/2�DK��ҀU�֭�*����O�0��[#����	��J��g[K����Rg�>+�����=�4/;�~��Zp���k��8���e�`B)��3�	��	�rW����hs~���s':�/o�2��}
�� hL[�},���|����aeZ�j��+��(�^�Zi�e.9��aT�[��vo=[U������_mv���mɫM1`Epأ��:�W�WL�l����ݴ'J�_�I�X��a!C�}V�{6��	a�;��e](���[_���#�x�ݫ�'⭧/�;��Ƌj�	n�_����F"��8+N0�����y�x�׽�(�����1R�
�~���r�?��� �δ=i�55��W�^��;b-_�gp�{�DWW�W[�bm.��E�s.O�|Y���$Z���r��d9i#$^�9�<^�T���7�?�{h;¤�����Ym�?��ċ,�:$�3���Xg�5���5�O�Z�2����dҔ3�ei��;��*
��h�*ȥũu��Z�:�UVOuѰ���r�>� �=a�bPH�-H��f����~��<!=��&�����p���ib���^?�(����l��z��t��7=d��|�(߼���?�	�C*^��\����������,k��c�	��[:,E�jW�2�kx�7[��U�� ��]�R�i�C�q8w�E�]��	s����C����݂���u(ea����� �pP���e��7_Wۏ��ŭ��ROYZ��uD�{I>ڣi�Ƨ�f���R~�a�4��i��D9�7c����Rj���B������'Y�
>�T
9�,I��f`/�|�V ����׻��q�e�c�n��VM_�e�m=����g��h����%�^�1�k�D��r�S�]Ys�3M�G2�������ZLe�9�[�eekd���~9��Ϙ�u��z��n_6RU���|,|��?�溏�4���WCy�g]un�A�Г�Nȿ����&1�H�|��,J�e��W	�g\�=�D4(�����DLZ��Qf�P��imZ�Pz	��'뼅d+W'&(絹D��4������r���@P�xY�@�Ɖ�<���7���)o*���2ў#ו�3�>(�Aζ�>
�ԏWn�[��i��.m�5r�A|I͢�� "�2�z� vt�|2���
z�z�fz9�sr�_
���<G��Q�g��!N�왆^L��6�%���r�
��暜�����2:���мY��u�j 綛BK.߾7�/�؛	�}���ftȵ��Ov�����i�!��\�<���(�/xaq`��q%>�7�i�{����N)9����>��RL��}A��͌V�E߭�
c3�{2���<;�h4�Z�㲍y��p�w�f�����Ld�"�������=���5���t/�#a�����Bۋ7 �R�g+��]�AI�����+/���) ���U`�X3l�1k|����Df㖃a�
�h�u'��%<��Ԭ#UbdjJ�X�vy���Yr׼�B	\�^b9޻<<��<D���W��k@+���H���Vɛ!�(�a�ᢜ��GB�\�O���)IF�z� ���S����a�˲�i2Rbb ��b���I��. ��fo�W�� ��_�{6��d3Ea�Cy�oM����@X1���"济���>a���/��1Y���6Z��{=g��q)�8�M'���^萳o��̈�y�e���v&�r�2������&܏�8?oz/*$7��7m�J�lbK��x�ӹ2 >,�my<1x��Ҥ;�։�=;����F7�j�8W]m\�S*�g����ͩԊb�P�W\��h6T�R�����?$�j}����;��T�N�|���^w�ʋĶ�� ���\�!���;<U5ju���*ty�)*/R��q1n�@��	˥�l�!���=��t�x�YƲV�$8c�ˁe��┗D��NZ�^[�wN���#���Z��Z��-����T��S��+\����QIf��&a�s)�[Epq`��8潝�k�5�E�ފKV�s�k��N��5�OT�����]���$���s�ƒ��|��4�L��ju�؞�r�>���>V�n7;,�[U�NK&2SdN�J�U���A3�U��)�2�4u��F�J������<����55V�I�L�� ��m�|4jg������嚴���|<�9�5#w}	�썫����4+/UgO�g�K_@;���
�%��e7v�a*J���ņ�gc\_�a>wzWhj��
b<0�u0����^V�B�Z�;��c���͓ŀ��һ�h�C�1��<�%�i���c�M��bm��pV;PaR��@�"�����Bc�ή��Fk�C_���1ϥQ
o���6@ɿ�/Wm�ݹ�+�h�'=T��gu�Z�[�#X�s��e�	��C]����4~̼�6���l�:H�L:cyVwe]���P6�P(xJ��,�L:<ͯ�N�N1ߞ�^=�=n]��~��[OT��@7��ܹ�k��b�����r}+�;������E�J(��P�޻{[��V��?!=(!c�z��T��?�ģx�H���uZ�o-�,��������G���zK�tIPj��H�B�}k�ZV��{�.z�����`"o�	-�m��*b���Px�_��&Ǉ��daJ{ɻ�ѝ��63���#��@F%�k�k��B�ͅj���ϊ �װ�X�Ϟ߂)і�n4�Z&�;�eI,'�`�o�����������Pݲ%�����X]{���Ez/�i2]�4YȔ�`q^����s��C�;݆ ��o����G/i��_����h�9I�	N�S��]��s��5��\Ȥ�u}}U�n�j�K�Ν;'�wMΞ=/gN�SM�Νmi�yO�9+�����D��N�xk1qnrZ/,�a_����,�n,���*:�\}_��?�3�ݿ��0�Z�IX��׾"������Y�({{�R���`�&�]�b}��`Y�`R����s!;ܩ�^4#�c@2k{tQc�y8��PF�K��Q�ꔮ��.g��}l�cgٳ��4������I*m_��:s|�,gKک�T ���W$겟�΀���.�\ۊ�4�9ujS3�'���s�qG��\�����+�x��L���Y�$�\����2T���yF��4aN�,�Mw��M
y�%]����툾9j���(�%�,�;wwdeuÝ=��\����[Q�"�ㅼ�����+�8"׋ O]9c�7����*�s<��H�A�L�\L�:Oƻ�R�y��-(��F~xx ��؝"��k�2fk���H��7�뚄Ɠ��ݎ6~�Gc=�n� 1�k[�q�*��O&lμg��{w�����=3`�*	n1����`B��eG�2u�2ޛ���1e㗮63����W������o���җ�RA�T�AІ:t���7����;�j�:���$���� ;f���!/�D�c]q�QvL��d�[�\�8k�Dw���N1E��ǅ�2o���äJv�l��i������O����
�2յ�J���Kk,�1��> ���$`�1V2��|�`���f�B�?8��:�2���a,�t�i�!�0w��$w�}��-���o��GR@H�SwO���n�;�\QK��5a�ם�TA(��]���B���\�XU�9���o���k	�8,ċg��H�Ν�r��$]䲶�ɒ<���ݾ7�2��/`��oo+%2鷳�U���y��G�?ڕ����#��te�º�y�Iz����&�������zmI ���ҥ���d?3�y����P&�T���Zb�kK�����G�������O?��<~墼xkJˊf�=�����kݵ��eh�R�P�0l�`ݢ�&�HŚ]MRb�	��tϻ�1��񎌏v0�,BR�x0��ͥ��K<=ӝy1��dSk��/C�����.�P��)�[-�9O�
5�eF�b�ּ���s��KZ��-f��k���zٔ�7�)�N���C)[;-[���99���*N
��2�g���P=��A���193ӺB��O,���n�H����˙Ñb���vD�zf]g�\5����@	�xk����Ң���?c�Y�{$�F7��C�("�\�ɘ�#�#<��O%<�ݕ����]mi\��xz�VY�0�b<�4����\8� 6O"n���k��>��ꮭ�p�P�p$zc�t`~i�WȲɝ�(�w��60~�~B��@Z��o�]�l:U������US���\�tng�N�����uUZ�P�� �o|�Z��iX�Q��ev<Rw�!��?���������SU����ʍ%u�C&���^=�8���c���0�H���;bf�B�m!O��]!ͧ�\�'5�㦝t����!�s��XE�fnOF���`oMqmr����i�(��2Tee�oY�c��}�JS�٢�ӾH�����
Z�l�R��$H��l"�~��y�-/�;#��@��ҙLY�� Ync���UX������L�y���I��<�J� ��M��j��ei?��g�kǲ��ȥ���D˫� Ɨ_~Uv��iH�Օ/]�O=��̦Z���Xa��K7w��D6�dt(wnސ8up���;Z�.�Ѿ|⑋�$6Z�	��W����wV�;����@>��0����Ԇ!�x��<)�|��t~M�x�M�~��dOp�?����㟽��Z���/�D��
��l���OR~x�;��^��;������9��%��$�W�����%~���Nz�R��6DL��B��p��br 3�X3�}(OQ5�^��JK��[	���$I/�h\B�[ф��Ka�B���5�k��>�#Y3N�&+�1�csE	z��%�we��� �	������l��ʹ�e�1�u̖������������$Q�e���8�K~�{�V�� r��Z&{jWBV7ຬT`l��-Q!�q?����r��)ia�B�����m%����BpvkS�$lϺ�}Anܹ�I��T�y��_Uk";8�W��@֝o��I�랆r��Z�/��G���תzC2MRd�9�	��!��'{P�\���%2,̙{F���թ�&���e�$��U)h�6�&t�������>�-ݭSz ����ݾ*�t��Z��~yM�
=�8��U����-��U(;w�������X���{�w�c쳶�ؼ��[�3�֑�Z.����r�"a9sH+�ɹX;ܫN�i�>��'�+��J=���_�'��5�99+��qa�d��i^=M�Ŗf;���cMŗI�>"{�"��>r��Ҽ�Cn�le�جY�����i�J_
��}���Pc��{(��x=ơ '����!�n`�N�qM����Q-o�4�Z7cĚ�w�����E�}��T�ja���luB9{���k7�>�M���cl�~�-�.�5ަ\<FO�*����_�Ek2�AHvCMRk�n ÕB"�*��ӣ�Z*�bߥJ��V�sŧC��qo�Noh���<��y��̩�t��[s=:4f�q�`X�T4`=��g?���yN>��O�w����v�C��6�59΃�8�Փе\J]��@O'��A��n�띂1�c#E�!��i)²�1��5,�b�ubY�Ų�	�(a�X2�f�3�M^�;���w4�Qz�I1�<�&��F�lȐ�i��ӽ���Wk<�<-��UY?uV�&gXO�$i��xv8=ц$ފx=�)ƛ
@��ϽUv����W��|q�������^�]cE�jZ��X�J��4Ù!�B��!C%	�/+XO��P���Nb��%�v����t�Ib���持L-~m
�l�U�肏��̑�0j�O?����G/���|�[ߒG�"O<��6b����Y�MW~�v�� �g$[_�](\��P.���1� {*�l5��\����x%O?�4Iѕ��޷N��\�{�c���W�8��Wz�|���kOS�����~Ҫ��t����au;��	�X�J��=��Ⓩ?!�=�����r��-���>�_��_�_��ߖˏ=!�g�P���9t�>$g~q�VOB�k�n�`Oz8�t���8zj�'�P~Ͽ�<S�MO�c�&4�~OR<C��[Dm٥��I�݁v��Nή��O����nן��rxr�Z3Wŝ�$M��_��y�?���/»u떏�������������w�����Ś�yN^�.>�H�,S��8�	���ϋz�
(�3�?���
��cVa;��i]NϞ-�=�T�?��>P�i�T��4�` �i
k�-H}.~h�1�@������a��}U��=Y�v��)_8Դ��d�����MY��	U�/��*n����eY�kB�_�@VV6��ҊUX�3%��Q�̂5���`!��R�
D/g�]K{t�����cA`<��CODē� �Y���Zk�Y����ī�ݦ�}\����fC)�s��E-{TSi؀�[?����X�q�l�1�A&x���[�Z�Eza�s����W_�O�����ӥK�Ԣ⑝���5'J9hܫ\�3w~���W}uyR`;���ߔ�;�`�Lru���	
<G������!��Z���.CO�P��T@��Al�7�`�/��P�]�-Iʑ���=�wM��#��mD�>��l�:';�GX#3MRs	~�
wZW�V>�%k:zT�<s-��Z�B���������W������&a6�l��ԟayz����D'�Wo��@?>
t�F f*m�|Ci�ky$?FK�ԅR9����Y��>ݮ���Q���\P1{�ɧ�s�����?�c9>>�?��?-$g&5�_�K�g���_R�Xߐ;Ñ�w�Yd
��
ȍA�f8��H���
o����j�6������y�����1�J�H3A��jd\66�d�;�7�]kē�^�@�0�Y�	>k�0�L��o�����s�_��"o����2�#ƺ#�����B�@�{��um�8�п�ͣ0����^]�uba��zװ]3�'ć�mU��{��e���֖~����yJԓ�A�9�p	�
���3r�AQa�)��,ue�nT��ot���8�Y���n�ū�3�����x}�%(X�Ѐ��L�P��V���WP�)�L^E@��b�m�̫6�~�f0�A�ZD�ͩ���5�y��u��*�/6 ���/���ٲ���v:��{nNݷs: h�@�H��ȑ4URyj��~q���R�jF��`���v�G�D�I�@#h�n�F�t��tr���Z��O_P6,@�\�Q�o:g����[+��Q忣��ȳm�H�{0����~P��,S,�EY��T��42c�OGT1FL �K����k�c���~�˲~7x�|<p�_�@2�!a��Te�^#D��]�M�L�@��-�˖f��f�NqL��@��
��� ��!�đ-�f�#g$��Q?�gt��̹��^p5=�@���#������U�L��|��i58#%��Ȏ��a`]˨(A�9�H3��(�c	j��a���$0s�X�0���B�]�z���P�y_��z�W�e�F	:re�H�1���$��=�j�L�8��x�̜�k��=�Wd 3jTjbDa��t�e�ʅ�2c2� ��W����0g1�JX䆻��л�\?@��]̪S�PG>�Yވ~������5���Mv�ң('�������$5hI�n�/v3$)� ��]@�kE��fؚ=�4Ӷ�=|���<ţsj`1��x�k���p1F�0(݃��ՑoJ��Ē�¬81ޖm�(�X)�J1�L��:!!.|"���Ț�M�`pN��ݘ��c1v�����x-b!CcL�sh��׉15<�>����Ը�J27;Og>56�q2t����k5f�p��RA>�v_�[˲݇? Fƕz'` ܁>b���	h�  h���>�giJܐd: �w겵]c��
�i��;h�d
t�̘�V�s� 4`�V&N���5p ��P����)�������7�d`d����l����ζ<v��|��):t$4{���M� ��b'�$ I"j�o]3%��!zo���eaaA�?��p�h�I�_p�Z��,ݹ)�ʎ��y�<V 2������܌�	p��v��*���cG-^c=��u�n�*�	���$	Q<��'�hIb�߶l#@�/�GN�a�=��5!�����h༝�J��(V I&nl��������wӚ��d:)�n}�w��F��X�7��ȿ�����~����G=p�_��#4��)v�#@B�F�jA�A(�������'�o�nX�|P���	�<��&3�)}1�t�赙�g@�Xd��6�$�S���r5v5�^][�i;\��L �^� \�H!@�̢����G�Xn�Zx_c�4FP!�1	P�)7M���r�K��e�5P���
=]�i�W�ɍ5�����B-�~h#�B�����`��}*�� ��`�l�Ga���n6�m��i�Gԣ[XV�`���
��<��-�l:=�.��p�yu���iu�Z
)p���ӨBd�g�Y��^f1v������*��5AR�E�QKz}��#;zT�-�Ƿ�d�2bY�ޑ�@�!h��>C��s �9n�	D��@>�u���T�sH�a�9�����b�8C3���vr��>�*a�I��COÚ#�=u�nh2m�bKy�g��K&gڤ b!([8p���w�ܚ�p���o��@�T�]c/|��7/����$57k�Buhm���n���
�N��|��(��W�{SQG�rxs�!#�j�$E�.x�Sb��͔B��='�G�^��j*���\��7n�>���f"��g�z�q���txhY����Z3bAu)4{��P��
���읛��q�3���2G��p/_�,7�]��}3t��^� Dq@FH��P}��T{'ub�.�	�\��r�;���"���?N:a=U��'�^"C2�k�18ꚼ�q�="�U�gߨ�9M5�Ҧ�5��B�R��+�2dPýk'�m��@d?�iA��8~�0Vvc�)^Ǧ ��2�|e��X	���?���VD	�t�������*��D�x�F�6���v^aLt��RV������;��=��K���^F� ���� �蚅��M�DA��VG�eR��:��Z��btEl`�� $1��v�O�cJK�2���D�˧�Ź��H��-�^�}.�1��ؑ9��υhq\%�c�3��h���>���|%.��&���9S��'��0j,h�\40���́�f�y5��PA�.�����އ4=�SY���}Ȇ:�Z�,�k��RٓJ30�w�ng�M�j�� �/��AG�n0�pT�;�D�ϯ]�H���>��ޣ���ԧ�����M�&<����:T&K��5���ጣI���Y��g�"�33)O>�W��������6|�W7������k�Oه���T���¸P�x���q]��@,��b(o|������Iv�&�qb�peuIv6���׳��L��PK �H��ǂ����d5��b�m�; ���쬈����b�N�(H���}�`.~�I�:1��8ݍ���o^co����JybZ��O��s�`[�~����wHT�H\R>}�m\�:�>�灛�u��k��_�!t(Y�AW�#�8�̎�g8_P:Cr��1��0�z{�ժ��A|Iv��}�g
��F+�%k j����=��s ��L�=t�:P+�=�!���u)�sG����F
h�k=1;+{���1��O���cc	S�} ��(�`��WDUE\�c�'fH�aJ&�������=vg���z�X���i�A��T��0��M�b��(fh�(�c��b�Sv��/���d�ؼ��<v��10����q�NX�p~14�ٿ�Fߝ1[��:Q��{����ц�h_����z�I�v�G�+(�iH��n�'!�b꩔�,�ߗ�������q]�!*v��N%�ހr���&ەf��VǘF*�l��b�h�HSNH~z�<�vfv��j=nn���f$�K4�V�XH���˔�B�p�m�")%��Ō18�3S+@83P6:&bOțh��'=8���K���Ǳ��10A��!]��A�zwP��FM��f�s�i�dimK�'E�2��:Ri�����@Ô_=�����N��l�ާp`�Fv��M5B��t1�c�e��p�%�LvV_@,ߏ�"�˄�Ǐ�)��7���U�x����d�UÜ	%_.I���)��y�jk;��V�)mK�i���D&+@��'����I5�ȑ�QYک�zeG3�2i^@�/�]��<�620�����8R��O���!+���D�	�<����Q'��Ե*�m2���7�a�z��&8��S(!w�{W�e����Ё�@\�6�k�����T�۷���TJ�����o2�gA2��h�J׊�R��u3�s��I1�}�;����A)ȹ_�"�/]��%���y�(5��R�\��5���qbU�W�F�8f]�Z�j@'��Ee"����J��E`;��[��ޣ��rYÞ��,Ld{�S��O{6���������i� ��S�{��P�> ��S����^^� j�g�?���y����z/R����2=9��oU>��x�D{L?L��F�	���>�%�gS�>'�[,��i�LjH���e�a�'�<q����z�`YN8;��� "�B�Y���ā�Qh*F�ӻ��:Ѥ'�s�8x�w��߃^�m�(���b���3�"{��cF�K��G�ʺͷ٢2:�NL�e&�8��DbC�,�{�;P�⊂�(hP�������/�������C�V=�s��F�p7]�0�pA;	�2��gɾ�Q9y�	f��}��\���F�)�'=�֨�-FRF:y"������:�!p$˦#�4W���E�+e|rBR���f��k-dx�k�d2CSFc_NY��~�?����� .��Yb&�q�|��ЇG#Nxd"}��C�ϲk{���f�+�)���m`�� ����I�e�p��P	3T�0���w�6K���Y��i:���q˔�\s^��1��f�Z��������O�4�`Ԃ��W<:�[*�N]R]"O�V��b[�=k���G�efn�#R8G��aH��nW*rO3�b8�F�ű*�7?#���P6��I�Փc�Z[Վ,֠\�d��gҕ�f��j͌�&dT�
���힡��'D���!H�F�SD���Iz|�y��YF��R�V�O.~,-�b�x��D��w�۬�<"9�ك����;�~���efj��z��.�tzq)ۢ0��ƎT[�XU�3��	.����my�ͷ����?��>���TQ���ɓ�o��3ې�:�Fg�D�e��"������o��m���҆ E�?��pj��M9��o��SS�-�w�y� /�ڴ��^��E
�h6Ց	
˗Fy=������Ir���Q_6�7����ʮ��Ǿ���$���R�葓�ѣGc������Ϭml˿��O����ڂ�t�"c����=��2Z z������(ܛ����}�BZ\�I���5��RF��ǿ�Mk@�*ZڜU��6D_#{�(¤	���o��#0���6��T�L�3���n���l�	?�> ���LHo�*�ڋ�iW2��?7��H�4��Lٮzc�{�j�:(�&�G61&�����1�o١�Zz�BR���4�m߶l(C�A-�'����}=���y�v�j�Z��͌�^�������T�x���8�/q �����Ĥ
Ԡ-�23��6�N�@FG��7�27Z���xD#{��~[�^���H0� �	�]��,2R���е�L
�Qp��D���6�0��:ʣ���G6�g�/pc!�{��d��޵���>�-w�_�� /����,���(��쓢ӷ��0�y��\ۚ!t�5��@�B/޲2,�64��}�)�6RAC&�i�̪��5�,͐��Ꮻc�@6?����W�Q޹�(����N�L�]RD�& ��S�Ե�`�d�C��h� �u���
n�nĎ4Y�0G+V[ ���Z]^"��������� ;_��$���cϕ%a ֐�A`C刮���xL���N}S��H��fG4��s�l	��"r��C�K��ߖ#�e}�ȹ� ��K��ʓ@r��!��çҝ����3ױa��L�9^@bXK ��桡W�2hw�f.]��68LV K19=%w��d�A�dyvd��<��~@оC6;�.D�|��z#�".|��dYyṧ����26=+���V ��j���XT��s�5";m��,y.���ruC>�s��.�k豷���yǧ�ĩ����/s�Օر!������m�~>��e4��"Z3 h��9�uC �)X��i`�A���}����u����벬�(`�NM�������Λ�X�+^Z�IЏ�,難o�8Bn�Ш� �2�)���p&;���5�uR�K��]����E�X]�{Kw5Z�X� z�1�h���T$��;�Ps�pUoƖ.�A�uC��� 
�j���<��C7#2������:@�k���y@�X�rlL9u]�=8xֆ��q���ߪ���~��}z���Z�e�T�Y��$LU�Zss��WpݾZ�y�X{=�����Y�;4��Ĝ� �TJ� D���a6;Ф=���pP(�z�{'O��U>�C��.8o�+��^��D�c�d�7s�%n�#Ƀ�#
zn|D�G�'27R�Q�Ǩi]��"D��vH'e��-.�0p%�c��������֎T4�Z(���d塇���� �e{m��W�Ɛ%�Jq�a>�7us6x��7 �"�O˂�3���$�'����M�y�����	�_�ߔ^e�Ղ��QIזd�����������,:���)����6��ݿ�E3��-S{��j�R����u���xr K�D�g(va��b�mH��]u��ʧ5��5���!Y�75� (bDJ��� qml�&��w����f�N�8S��n^�.]V�@G���`{��內��	7u}�;���T�1��X�$�k�
*6p!˕M���jX�@�F(��/I"�ax��$ ��LD_/�7����6���7�T�1�� ��N�i���#��� ���@����xd�dypP�i�Tȗ�fQ���OɊf�̸<�r�L�s!� :��m�o�um����1�ކ��9�~�A*�+f,.�v�I�	�*��=���絣ϵ�ϡ�� %�>lȂB� ��^c�Q��k�g�2u��^�lT�/��V@������]}&���~9̽��v��� ��k W��`>�oA�=��f�6EoP�#m3�U>��siTkb��"���hI��tA�;gp�ρ�O�+�b�4�u�m=�����z��\�r�0�8#~�g[����UeЂ=��{���`"�#��u��
�ܝ�H��F�rf|�f.�n[�H�>-]��[�Yp�t�i��,�S�$���F���nǉ��A4H��T�R)�����4\L��~����o����}�Ư�ί�6����@i����C�GH�fd@C�P��5`���ufALP��)��˥�Z����.��<��P�̸Ԅq_'��!ч��+���щ*P�04�;��dV��|IP0��ձcG��w~��4�w �Q#�	d�ƭl!/�Iڻ�kZ�&x�2
Q��ύ��.����w��Ր���"�f�lT��-�4��L^�~,�x2��dv� ����\)-E�f4SO��zN9����3'	ȃ#�r��P~�v��s`T������f�4J����@ S ���Q�P�:E������ۮ����Pb��K�T��$Y����7���%���q������k��	6��ߏ�~\���/3ӓT�c[�]��ջ����;�R~�AD=�xHk�j��W*�1=´+;��4A+��/�g�ἩI��M���to��l\�x�챜�n�1B7"��t8�3���}[G���=���8����Yg�Q=vXnܹc��zώ;&Ӻ.���X��������!M�Pq(�� �[��HV�7�7����D� '����ˆ��� oЦ7 D�~,iF�駟JD��,��-7�S�݁���Y۪�k8� 0��q�kD��@̨`S,lE9�>.�4(ܔ�������՛�_���A��h�c�	P���g�{VF��6��QG�;N[1�{vM����|���U=�"ZA$<2זTq$ ߤ<�̢����=��jK��Ɍ�?�"��w �Ny�D�^�@�k�4���G�D�}S�卣���ѩ�O���K[���ʎ�KV2O!�G�'��Yl��)�=��RR�A��g�P�d- \ɡǙvY�F2Yi��Hc��8Y��
��Ԟ��b��� �%*���+W���D}�fKyy������^�z~��][DOOO@DG�繹�i���@�:]�tqN�zkX��y仾�R�8S�=�Z鑔��J�ΫsWûU�fuG��iVZ
���'%�sd������x���9K��a�>v_Z��L��'O>rƔ5�YY�'�o���l��4�Q��Q$�ݲ�����	a���i�F�g&_Էl�5�k\� �}��d��V����$�`&��B.O�rE���V�Jj���2l�P��9=�ٙY�я~$�N�2Z��k��rO�+BMI���0��#kt6>1A�Nr�8��U$f�vr���>&�s����x�}�� � �=z�Ȓ혀��*1@/���WA��
UH���t�`F�Í�Up�x�<a����D�&9�P X5>V��|"j�c�yln�#O�O�t>�5�#[����g��
Y�͒{��&\Y�5��U=��2�65�򡻀2�������S�={��kۧb�G�]컞:�K��X�Ǡ�)P�C0�L�7���q�㣣2U.3()��܇@���-r�Q���x8����ٲZi�i_�x�,2w8e����o%�:��P��ȑc\;����g��y�U9��eFq� k�$�3�p�����q����Nz�vW�q�-a��D!�5���t&�w��H3[�ow��a1ӑ�1UL[���"��3[���%������8�B �>[��1��	�.�5J���Б}2�w%�%�ސ}S�Pa���M��'�������T�9��'҃.q�l���#$OY7���8��D=���^���ՙG��.9y�!����'����dcC?��g��N���������z�N�ȍzG��i�V���v��5f���#��ދ\I�PF֏�O�\�Mٹw[rj�\5��^FZ�Hf���H��o�Ug���7��<}�!���u��ɧ,9��=��e�#f,F���ؤ�h*�V<�4?�uH���'�"���ô�6����pd&�O�$5�I������1|�p�@Sm�r��2<�8��@H7�O��:qR^z�[t�nJ��k�;��H�:!3Hd<�j4���,�Y65��i/�Y1?kȃ�g�ئ+/2�꘤h@A$�|�"�J%cLt�1"Z�-2� -���9�{4@�:��9��/\��؜����%�����6j��^�h��8�TA��<����|)C���Q�6�����\.�w�������O>���#���ӧ�f��^{U�O��Ŭ;Y�� ;���Uo�8*��ьO��L�=���ɔ����QD(�V|��,9��)��^���		z]�u\ݽwW����:�c��3O2 �TK__`�Ғ7߿ �}.[Պaecp�NV��+7���n�f�YuҐԝ���?��.��������GׯJ�^c�C�Y�9c:f�;vrt���i��ə�=�A&�6�KM����J0$���>J�=z2R�K��!�?�-t?�P��=�o��_�����C͘����W��9���׍0���关�DAd���c���6l_�-����t�4kبud}�.˫k���`��<�0�� sa)�6���ű|f���{}+��~��y94=)�����ɲf�wn���d]�|�m�	�ia�;�������KO@>*j�����fü�fRj�;Ӏ!l��1�o^Z���TmFp�P��UiOLJ������d��=��[ӭ�K��r���C���ߢA��r����J�e:���X�]2΅��jl'����>�>bV�C��9v�!{h�D-f���G��l1/�����einX��
�=�#�ļv"�&��e�: ��!#�.����ظa��L3�u����y] '�:?�
�<9F��٦S,���*���"�zVߔ���GE�%����m�̦���8���U��w�6�h|��At�����]Y�'��V�`��!'Z!�&|��W8����\O���d�p*�nn�Ґ˦eϾR��w�����?}�|���5�l���:Z*u�A�R��o����,���4��2��G��瞓O?�$O<��<�����׍�* U�k�/_}U,��"�$�P�� ��ᑲ�8��o��P�J��tfԮi����/Ͼ�iU�e��mNm�8��V�~���{\���]Z�Ԁ���y@�3{���P~��yu���zM(WHm�� �8P}ސ!�Ԫ&��5���t*K�,RT�Ǒd�I�� �Ȑ�=a�=���1�/����FV1M�M�L���
�2d��%4�\�ۂ��5� 5�^ȧ���=���x�п��FN��.z��0��|�}Ȍ�d)/3#j����P�Kl�1�n"��hrɏ�����cjb\jM�r�,f?|�XB���Lx�Mm��JA��f,O<rJfgNK�A�`L���/�s��'~,��u�@���ŸX�(5;;۔���4�{�#+E����JS$Nw4�A�LqF���JK�x����Y��Sن�D:+E5�Ⱦ!汦���Tϖϯ^1 <3/��	y����񧟕C�������ȝ{k|M
D��3J�:|&	�E��7d��+�&�!�đ������9`RJ��xYr�;�Yu���I��%kK˲���ƺF�z��9pdpj Wsh�'�:�t`�-..���4{�@E���nvrJzV[��.�Kh�nv �e�mY1��f? �\��Df��0f�E�Z�I�j�Byl�r�Βv�-5u<ӓC]y��s���������^?wN>B���mѩ�`��|��\Ӥ4����kM�G�x t�~�T����ʟ��?�ɩy��k��k�10r�yߺ��7���4���uև�9>F�N�G'�W�`������Lk;����l�o�~W�٢^oZ��d}F9	��R�y����;3L:�9��]�J��!C�������'o�~���談�	dbzV�6+�W�K�́��ԣO�w�Cy�3r�T��3wS1�KFF4�,k�>�!܃B�(/��2�g?����mpd̘���ʒ^�=u즢�0�!QHh`N�6��I����4A�'�@"ޓ��|T;��@�`�>�Ӏ2�������%���;�������8��b�7*�9��B2�s�sƦAO����%ٿ1+�%���I����Td�RZȕʎDj($?"Uu~��^���m�	��c���b�G`�U)J��22�h&�ƿ��_IY��:$%u��d�G?���s�᧗��as���Жefj�%� �Zu�aܬ�ׄ�'��d����H�Gu9b��#/m�cz]�{@r|L�i\1Ǜ���G��Lv�mJF�¸fk������Y �4�����\�zGz�WԪ�����3i�8k���V��S ��Db�֡(��ħ�$z�~W�΀���S�;�����YHN��3s���Ƶkr��5����7�B2��:�/>/;F��9���}��7��@�Y�!A��Ȩ:T]Wu~~Q����jK�`W��G�z�����u|�& �4�LA0c�$/
h��o0���8.x���q������)���>q��i@�oY��=tP����Ҷ���f½���U� `���	���������c��6Dpp�sy~����������H�ؙG����s���v]�3�@������?��?�ɱQ���{�Z3^N0� `@uIF��oa.����e��]�+�r��)�� X,�2�G ���c��F��<<s0�������C@�g���Ɓ�g��m4�gf���>�k���%�զ~\�L�$ߍ~_��Ok@�_�2�x4��o� /<��L�G,C�6�3���ſ�`�Mu��)H���u4`lp��hېT��&�P����L��<{��'$R	��p?��-�d����F�'$��S�J���gXLk���_׭� d48	PX������T��K4.C��N"�n�%d������|���M���ʀ����E|9��_�~�{�?�\^��k�Տ�:%��׶Ը��|��F��1�r�}�}KSN�9��\�n���y���K��ӧ�3�/���� B@��<��R����렏�X�D�>�3��f��s���,��g��/_y�T#�A� ű�F�K�\���5+�b��/�+0�b�<K���6�uJB�5�o5Z��	�Hf�&���������Yk�&�`l��)Ns��xª'�]ʉGւ�� �g�rY[pő<��}�TT($�� ��=���ޣ��y9r�9rB�'ߓʶ:PI2��8�Ѩ��Y��{w�����A�>�P����hW�TA�/L�xjJ֝1i_���Vd>�9��$C��~&i� �����17�O!tsO��P��F�ԯ0𽾡5u]�gM�'30��I#�FYtQ����'��㳁(����Ac��Ē�XW���0�nq�m�g���{2l���GVAt݌��E���]`�=R{�7* �@\
�#BK	��L.-=\F�JrꑳR�t.�̀Wx��[o�VZ�:��8���L���B �1j
 �@.�_��ܾ}W<�G5=�pY̡P!�
���Y�o#�o��2�����c�k%.�ooU�#x���ek�"}�s5��H�۳s�r��A�V�e��-�л�F ޤ�F��>'\Q�w8���-�}���A��KN�����0�CJaDʘ=���%0����x���xp[��j(�J�2d�m�W
DkF3��Kd5t�_]�J�׈�U�I5��c�f���ت5像>�[2#�	3��t�ژeb)2��ɸS���I��'�>v
���O�H؈Xj �/�˹�>fO��Ò���,=˂���I���L���|H.�����f�(՟�pQꚉ�GF.g�qN�O���s/~��6�8��q�ߌ���NtT����a��B�Ҭ	�iqy[��ࢼ��yY�ܒt�,�f�n��m�Y[7�)t
^�}"�����I��� u��
�+��@�$@k���������� �-mjd�E��4��@�H�є��ߕ��Ui�k���Pd�xf8�,Fx�it5s�����?+˂f��ʜZ�QרĹ��n��@�)�P��β:�nt���M��a���h����S�F��=����`��#Z���8@�L0��-�h9��jfG��������f�������R!���Œ!D�뺱���r���)��h�� �AL�2�w�x��u��i}��<��St��k��@�W�ْ��I�Pg
�_�M�e��Je[�9s��Wq}���\ZY�t6+g{T& j�{� ��lI�c�C��E$����6	2b0��s�n�,�2CYX����E�G�(��5���F�\3���\��wޑ�~�`U@N	��@�;x��4�N�� (2̊������>��1Aƀ6���g�!���f���VBR����w����hG4�h����+��!�0&a Z5��Y/�H�_�����#�B/��Ь����@�NL����Fh�����|�Ź2:���鄦��!q�'\��b�Kc\]�v#��шS���Dԋ�-�S�agI��:*�Q��	��o�p������-[��<r��L�T�70�0D.G!�+�C�h�Y�����S&3Ao���y����y��/�Ȁ�X���R���cGV���<�����0c��dj�)�д4C���r{iC�|����Uu�;R��O3�H��2|s1���02��!�e� ��E�[��i�$ P��m*$��M���&Ȑ��� ��RF.�C��f����T��hӎ�cxY���P�2�#�`X�c%�
��VV�Y�XۻG����;>/��(pF8�M�����l��ҧ��.�A�� J����$Pێu_	J��r�h3���pu��a�U�ֿ�|Ƴst-�|e6d߳���d�����a������-:-��	��?��������J�T�|���W�^�����&%`O=��_SSD����%(�ϩ#]����[poff��w �A�<��61�}���"���W���׮����_�*&���3`�ԑu���r���v���>[4�u��k��������D�=7ְf��`���`(�(�.\��|�] �&g�Ѫ�Xd���4#c�g��XK�|	���\yd#/B��9����� 2�'Q���v��]���3OT����ޕ��q��Q5�d�Kd{�/ qH0!E��}+�<8���C�� �<�#k4DN��H6�ѱ66c�)}�gP��Z�x��4��Ѫ0)��|g�t9�)T:b��8jN���f	9��:�Q,���+A�v�n���k��R�ɝ{�����e���P`(�RF�P��董$�ѝ��u�z�~�
8���^��@�C�����o~��9��n�����~*{gg�j�%>$��@ �M;�(�!#�NP#��f�������p��k��Z]���N1ÊF�4���X�z�Q�BFe[F"Vb�k���]D+��
��)/��qS5@f�j	���k���I�%�)X�5�����}h��*r|�T&g�R�z�����-'V���F�AWiu[&��d�8+d�y��D�!�~�7�0�������t�.�/�����$�~%Z���$m��"*��U:=?%Y2 S��pl��N�v�O��	Y���A�ŀ�
�9HLS����cmM�g�������#�B���l:q3��d�A�`?G5cg{��qᓏ��w�˭;��U�0 ��K/��4���/�I����|M ��/_���.��hc-���Rm4住>���s��a�� �ʹB�)�l��Fx�Z�2���׻y�&�׏�Q`�Y�9�S�h$�>}�s�X�(����ҽ��ƶ~}��b�r�u����E�b�_�ap�����8�4[o�3��KG�'�qe�Y7 Rӳ����*��AI�K>l��O<EY۫7oi@�U��EVC�Mc'o�B��u�������x�п�ؑ���u��}`<G7�_���mII3��FA���ۂ�����?ן5*R�L�������.�Y/��4�ҿ����!��P�L�������j�9 ���B�T�aԏ�F�H_�;�UC�+�m5bk+KrgtDR1�F={,R�y�d�fۛ1\3���G��F��9Y[�DH,�e�%>��z��]Uö]���c�Ԑ����!�8�dc�Ŭȕu�m�fv:@oWC(�2� ��Yf�"�Й���'�od�l;��%�d0�p�9���B���A�A��z�;D>b͠�a,;�� ��l���6�ѯ��/�O[�Nv(2- �Y�ѡX@P�Ӄ�z�*��˲�]�L� =�#�s��<#$m��4�$-dnn��k��Z��)ǆ��2wĔIc�3z�x��l�3&�椼���p��;��G
�d�&�u������w[��!Ԁv��k���J�@�F��5Z�|�	g3)f鐍E�׃9xO������k����{�h� ��Xf��ֵ+�P�5K?�9*6�?�� ��?�����֛��/�ч��KU�!� �mZ^�N�ח������3G����O˂�6*kYݻ��|����9rD�w��	��pnXA�
'?9=#���o��Ɍ�y�ǕkWO"�Fe �E������?8v�(�ςE.5�H��=�8�Έ�{2���,������A0�֌6��N=	ؒl<	��v�8�ב�99|�(ER>�v���W��9+�AՈ���/�}W������ʎ�KA�{ ���@�̗ٔ�U�%�`4�e$�@y��"���R�o|��kY�^ssYں
YG^z�y2�ԥ.�L�{����o�n��ZC����t�6��ef���3�����`������uD�s�ܬ�̎����2U�K��nD��>#d��ȌV�Y�d�����A!�z��]y�Ïh��`�B�W=&������XY���2?5�6+���,2�(Τ��K��ЂF�w[���w��qkq�Ƌ�0�>/�23��>�����X֑�*���(F���Ѐ�R����RԌT'քK��-�&���l���j�$�@����iA�Z���ZE6�We��V3PքNx�}QSڞ�����G��+t�h�HLjT�絥�������
4�פ�j=�l��N=ϊN���^W�x���20�ѦL�;E�#F��v\���YVO�	����/����*[���L�NA�ĭ����{dsyU3ԊL�ek�˾5��
�C��g����Y���8U�%2 Ǒ��M#bJ�8 O
�!�][���{he �>�ҕ���L�_�)�>zF��{��5t�~��Ԁ��﻾]�_���u�{�L��Kp����� ׎�V�}D ��!�>s挜��z�Ј�X�a}�5y��Sr��q:]���ooo�þ!w����Çd������u�=y�w	�E�O�YY__#�n�P�����D����}*�7NtĮ7OAK���͕e�X]���6�)�J��	�����ɼ:�����n"xۃJ�P�zc�U+V�����u&`�oC%���?1������84+bGt�T�'5*}��L �SG�Wo��7�K6z^�Ҽ:�	�f{j� �qط����6�  j��#ɦ,����F$�����[�r���F�%����G�K�H���k���bF��v]�.���Oʣ'�K9�IZ_<�6����w#*�a�y�h5�jLR�y���@%�`"��Ϯ�ǚU�=����>5h#�*��Ԕ���#f��\�i7X�-�� '���(b�X�v$g��\��Ͽ/��x݌X���@,��qR9��H׎U�B���bc#1E�m�d�߃L���C:���\yL�hB��7��YS3��VWV5���VC��A�i2h�s��ܾqS��j���}
�)~��o���v�ݻ���wߕ��U���;@� �0��f�$U��+;.�(�q��:x8t����95"S-�"�Q㹹�f9og�Vܷ�ny�Z����yxd�D�#�30AP�D��{��`*
i�ְ��� .���L)O~��E4�眎���p?�tEv�9K:C@"� ����X��������;����>�b�0]H��㓍��mnȯ~��v咬�[������.]���nJ���[��4sޮ�o^}C�}�#"��ݠ��E��!C�]�N�9�Ν;��[6n�=�����i�z��T6��������-�	q��Z�t�l�O��W������Z /?"�˚��^Zյc�aPR��+�ۈ:ۓǎɋ�|�A�TQ~G�Ө7eemU�xK��N�`L� d�+t��3����Ou�}���Yz�0����~<-�#�Ɠ>z�埰&혤"`*����~�����жSqI^�*�D�c]��e[޿�7�[B�����8����x��ԼL�SU�8��k�R#��S�U��?p��I	"��	'����r�\ʔRS�3G孈j2�C��=Sey��Y��H�S��U;�����Qۆf�eL9� �fS
��<u����ˉ}<�0��Nr���f�Dփ=jh���*���H}M����<�&��@F�P�5���`I/�����T
���D�3xѯA�Ս���A��s*�����<zr/��#p��ͺff�Ǥ��t��`W?ϒ���7�gѐt�R�b�� ����|�d�A�Ͷ�Eʶ�CG���FO��%�@����ԺܺqM�ݾ+-{�Ō���g��oG�������3\N��ϯ\����\�eS\�����1�Rz_�0�3Ԍ��i��6:��S����Y�q������b�X�^gG0������a�ݲL�Ul{hA�hG�����Fa���w�Ya��zO�ٌg���/�P�âfz9�����}����]V��쬌OMR`��.6��{.�B *r�+H*8$$����ق�`� s��A��!��J˶:����t+�z��?6�}z�>�dDa���^���a��;��Ee�;��S���r��MY^\f��� �zl"���ԁon�����iH����U4�ugIH�C�i�	rY�/9)��R\�*O>~V���濖C{�dcm����Pg<���'N�xiL���Aya<U����(��\w+�weE�}0�a��e(�R��yQHJ�I�(q���"�3n�,��C<M��}�.'&ޱb��!��3�M��E�������ׯ�x�п�v�)�*c>�9��QH}{S5pM��1&��� �.�^�A0h5�w����4�����A���� t�}nnV����XG�QU*�<2�e�����1�mE}��_��|������(P�8-[�ؑ�o�?�b�F
�F����1���`=G�`C�F�.���j_7v��+kr�w����읛~�10�`Lښ�8�!x�b���!�jt,#sS���������\~{񊄚Jg݌���}i����M�pp�*v`�������-��P%<�i�T�N����q�4Sl�=G�\I�e5r���z���zE]3��k�SD�裏�܉�[U'l���fqr����3rg�\�}G�
�7#�(��#��@^yI� �>��<�G\�ɠu/������,Ɉ�ù���#BK	e���>3o�":H�sb�l:3�����Bf�A\.G����qNL�� ���"p�>xH��o�]aE)����4�r� v��,1�hG2g��u���>$���H��o�I1�'�0���~�"xr��#���@��;6�N;���;�cG��p���	鄁ntL Š���h�Sa�M�*Q��#[!�zm��PG2b�����o���E)�����,޺A��Jt�t]=��sr�����˲����=�م9^�������_0�)�+j��>���1��;�7O��n������� 焺
� P��l��K��������8�x��]�?�Cׅ�9�z���8L��� ��~�1�$ KZ���y�/�)���jZ�̫5W������ڲ���V�@48f��j�rP��X�f��M�r��X������3u�����F(�i&���/�T���:�pP���(� �h�3�p%��Q}��C�×�!�Ŝ�qn-���K�ɇ_T��&�zp0`�Bf������c)`]�Z�ܖt�D�Z�jzwF)F6Ձ���������N�s�)��M��Aɉʅ04-k�wdzb\�x���K2=]��G�O�W���,oV��N�e򴗺��%�bc��4��Č��%�6c^|%�Ѝf�$Rf��}[�����C����BV��v_�Æ:�K�0��2��DƬ�g����i��焬r[�K�z>���<%��J���S/7%�7&ծ+-Ԭ4�x
�p@Kez�ۑ�ŷ�\@��nC���=t�j�Ȑ72�+;"9�0�3�o�F� �1+�iVd�(#�[���h�����M��kF`�	����<�O׺#wW6)H0&E8�(�Kýo&�vg� �@��Ɩ��n�`��L3XU�� �8�g��D&<'�����YmI�^�F��iS@��1od�P�^!�6b5��Ν��v�q�'F�l�@y}�L�yu�y6`S,�=�~�s���K�w�:��o �ڕI]??8q�T9̔cd�JL���#nj�t?�M���ŠA~�~2��ɓ`.9���>)�s�}Fv�<�� ����g�� �������A���|�տ��šG++�n�Ӵq_x��F�s���m�u��%��Q��,5uW��~��A5��-�G��R���ц���c��T��Y��f]}��e���E��l�::�F=�f���3��zGzM�B�DybL��A�#�rY>2�&I$2���D8�C����z�Ǚ�^��<v��Wuӌ��e�DQ��ԓrxz�s�fW�;������r��mYZ[#E��nƂAA �t8��22$��v�~A����hv^.��^E�ߣ�ʬЈ���_]Y�ՍMf�@P���EV9_&'���+!0Nb�M�����!��o|�y9v "�'{X�+u���s	{��!<�ic٘�C�5Kv�U� Y��0�B+���!�٤g��4�rhTA�TZ��YmI#�4$jW�����cgKZ�(l��N	Bӽ���!5�@�74	d^; ���w��h04Q)M�3~@�nd���A~V�vNj�-5��e�&�V��i?�t���4���6��p��Y������'��C��kJ�2$�p]p��8��5�i ��=�M�g>�<K�P ����8�&	^H�n�W���^{��a����d(��2�<0"*p�AUD�'���v#4��+
�$��M�	�4��l�9�/�gٜ:�l���&ـ�0����24���`�bBh8-���p�6�Iʔ哹�X�� أ���%�1�D[����>�K����!�|��8���AT�:T%�1�ƄH�X�_�Nr�������R�U�o����1R�5&eu�G�v��DUmw�������v��3iÀ��(�K��0��#�pу4��8�Az�ygV6'[�?�S��>�v�q���Ugus{6����4�釶D�����d��ad���������e�*��N�����墤W�����y�� X�A�& (=8k(�eJ�-J*'!P�VZ��;5�>�3-0�E�]����Pw��F�ي�І�f��`��^�%:/���as����e	��05��4��vV���>&����pî\�&?��Ϙ����v���ETlu\!3�raR�ٔ�@�3�] �3���2�C�<B��<�  �QC���l�����7����:��p� 9ub:��jE���������[���Emu�d�[;�W�ɦ���/�D��S���o޾(�Ŋ��&�+54<�9W8
�B&6�(�	����IdRZ�����<h��q����Ј��9��+��>'�O4��o 4{cl�@1�)@U$0��8��L��']m`��nVD\��'�~x���GF4�9��,�֔�ƭ�w 4{������E`�FIWL Bc,��'�Y�c�<�?���ߴ���:R��P���H'1{��
��[F Y/�-��]P���]oh>e��R<��{蒏M���P1�x
�/�rf'%k�Q���I���	��!�/3A�x�D��d� B�=BF��,d�2�0��h����R>M�����P�l��*�!��s�D)�X�^`�6q_���lmv��r�37�!�8�4�T�K}PAv�j��H!/=,~�&[�+�T�	>���{�5������s��l�"��|scM:#:�D��3	7B��HZ+ɑIo�wK�L2����3��Y]ѕ�i`��$�q�l�VF�>�`p��8�A�f�9�UO����/�+��W���N�kJ�N��(���H�:HK 
�zZ��dˣ���F�z�H\�����F}G���f>�����y;�����wt����H�n�����Tx���p�����:���@�~lOC�6%L��sf��}�DY�~B��͍f��E�
���\�4c$�(XB M�b �,��dj�$�?��� �XY�_�vN��f�p��ۀf�t�2=� E�F��A6���8^�^��^������E�����������0��Kc��'�񳜯�kW/�M0��3��O>c�+�9���f���4�fNI��W�˛�}G�cߗb)'��-�~�E��-5"ٔ-�n0�5�X��ن�*.�s4��]��� ����O��C���3��i��`d��׫>��.��5�I��A�TW(f4c�������k�4{��꺬nnIO���;��_�=��� k�P�um�6}��҅�^<���xsu�p {�r�C�TP��H�j��b�kǹ?���Og�����cNn��ƪnF�ϋ���O���� u8@�/L�i�8�JGFV�gM��3k8 ?Gb%�̱#{���C$��7|�ȶ#;���v�]��������{0cr�q���G�zu0��k(%3crp�>�`A�gfH�J`d�n�V��z�s�5�@Ջg0ގ>�J�Noa�j#h�A��A�ȍo�`aW���=�Y����a���d������T'�nm��� 6�	#�c��8`��K�L�Z�������4:��B�)�j��%�I>'h������-�� ��b����`�0��㸚��qb�������k�����Ho��7�������c��v�j5��:�V�'P
�)]ȑ��S�����_��e��=BIHu�V��+k�\Ne���=1�ne�W�~�o4]�M���{��[�w59t��0����s멑�Q�٨O�F��#VT#qhjRF�MH�9��,G�"�;w���ֶF�"@Q�C�q�M��BH������:��fz�ǆn����b*݃k�����z�323
&+������w�K��b6V��1u֘m%[�fT�>�L��#���rgq����熄�kVԐ�,M�ͺ�����p � @���`6��UǜfvY��i�:�yu�����ǉÇ����D��衒qO߫��ʔ:�+�n�����?x���Ϟ��s������x��g�JFk�u��:��8803����̭Ӫ�`A������@h��\j��cڠ02��ٙ:QW�kU
�<ǜ��dtzZZ��E@�v����� ���G���w�����ҝ�||{K�mkГ�T�̙� b�,|u~�����fK�T��]�Nێ����ìP����~!3�3	�L�̶���F8`Җ��9��"��@9�ОY�������F���<&��D}J�fP�6t��|���c��k��ܜ]����6���J�C�i%��Y`��50�b	 +�xlm���왝���G�=${�g9�v?(��:H�󈎒K��z����B���������v���sU�ܸ.w��t?��AZ�!X@�&dd��{ou��L��_��h8���s��Ӌ$:r8T/�m7y�5]o���nߔ� �{�Y0*lxG�-����R�`�A����݀��R��o�۱��'��ng�̤�T1�^�2BQ����Q������嘠F�.���#�������<�V�E������[7���7�ZER0�햄���1ND^o���TC�r*_�@���2��?D_�X)ӟ�h�
a�2@љ�6'r��D6�;�/��ɵ>�z�U�bk�LW<�Yo��ah�\7�E��Ӭ�](`�������Rqc4�ld��h�l���K�P�z�K�lу��bUcr`�,��L����鵥!#�N�'y��5�t���Z\��:�q=���h�{�jC���p��:��Tµ-��\f_�k:[���N�&��D��S�>���� �y�����GdD�� '�g�����>vXZ������`�2}f�ˁ��K��L
uzn`��8⢎�����<F�,O�9.�:�V �7F��8��=*��:#��9"��<#W�\"��,��g��s�ސ���l7�~�s9{��L̔x��N��c�$[�!b��{��9�{���Gq�88q �Q:�I�iatT&f�J�\�P�k�����[�8��ȑf�_�Kz�(~F��ɞcg�-��F%|�����Z[�Tڤ��h���I75h]���{[rk�/�-=����z��)��m��}�]#�}��}1R.P5��6�x�2�ss�3�] ��-Ѯ�چU�����X��b9$A�;�(!{a�|�~ojvFF��%S s\��� �vN� ���]�ݷ�>j���q�	�#cp�@s��'��p� p��LR�b/�趃�ߍL_<"]+Z-!�y^�G!���ǟ�Ú��_�c^vV�@��O1�= *�6����I�L&��R�J���hQ�f&eaϴ��mʅO���
 ��>�'f.��u�y�~@��*�3B6�}�L`��>B/��ob.��2j?Zm�d�2� ��2���13A��`�%p�K(��c-t��4���o�����#y�C�a�2?�eh1�jO�S�!=�b�לw�Mv�C�~�VJZ���ʎ�͡G�g)Y�:U�u�ݺ�Hg񎤡ݍ�!6� ��F	˶5������Z@IIM�a��7�Vdd�^q1����؀���6_���@@���Z�d�X:���z� �N;����n�e[vӷ(��v"{�Uo/i�_�������)׺���k�b�i!҈���Q�fu���cV�ՑHD4�]�I�����-)��&�Ӭ��ܼ�l-#Y�Jmc��H3#�̱?�_5�7o-zH5���4J�A�҇4eP����9�m��o�R � C�;3-{'ǥ�O�Y���E�{��s5����2������5Lӌ�A����F{J9��T4�K���ӯ�k�8ל
\�Gv �\<��2��0��ܾ�98;���N��\ʴP���z�,��������5ˋuu�L�h�tHO{��*�8 ;:9s�3�3�c԰n�c�c%�%�V���G_�v1�����5;GI��0���|l���m�~C��&�R�l� p����03�i������A����#���0dm� #74�Z��b�1����f�w�ܹ�%�4윴����/���Y9N�*Q>ǀ#�2����nh���X�e`#F��d���Cv8�z��/���v��2L&ef��*W(U�dx�(�5�~W���9y�܃�\��s�v ��@���}��jM�/�޳ٲ�{v:���9��	%����F�0�]v��`O�惿��?�w���8���%QE�	��эF����ܓw������$-��O�`����s���}�����7�X���[n��p�F�ewfwXSʲ�P���x1�XX�<���i���7u��ry��	��3��>��1� �H{,����5�P��HF�'�@׎�I��,-,H�i#_4��L�z��gdE�C�g/^z[n����r 0B��pdmp@�23�Ā9b�
A��>�	��җ�$��wW�N[X�����7�6�
�Q�o}(�oIO�$�`��ooo�_��2��&A��i،s�`P��dN������(�c=���_}�z\��=F�/*lU�t��)Nt�*�hh����Դ�zm�칓�����|��?���e��;7��ϫ|��ꪄ�.�*����Г���BCf��
�C�Ό�����셺V!�A=���F]�´����~/�ȷ�v����O�Sգu�p�x�A'��A%=M�vt�ލ�����+�����mo��Ά���賳G���G��w�C�@�t��ʳ����<X�;Ʃ�f�srtqQV�eJ���ƚ4�aE����}[7��G��������W~(�����l�����J�d��Y��N
�d��g�=`�MWkrxyY���K��ٖ��|S��6X����{A�������I��Lj�]��`~>��t%���������Ĳ��A��Ԍp�k��"� w�g����(S̃�����V[v�z�B:@O>QGѥ�]�h_(˻�#��³�4ȼfIsjhA�[�/Q���,�Mc�.�[��p���U>�}̹�����ȳzK�)���P�|�lF�:ة֌�г��b5���uE�Me���][U�:����tƌ��H��&�p ��u-HWu��d��F�֔��9�֘�W@��f�X�,ycVJ�J�C}&@���#����q�; YQ�oM�A!���|�x��ia4�A��H9N�@:��9���w����e�s�c}�m��0�����s���{�0�	gR ��U+5��$Um���|����9&9����!��󲿷Cn��|��٧/��c��Q�J���zT�ߺIb���u�p|���@��ȞqD玱/��;q�؁�t�8�ٙ���S'u_���͑8L(���,�k0�J�P�RV0=v8�eA� h{S��f��B�i�rJ�#G�K#�����y�_�V�T�(�A�/�C�D%��_c耒�+�{��a'�z�Zd���7�駟�&��u�3�Q��~W"Y�Yh�Ie��1:bo?��`�j��B����F�^���Wt+��a����y�����Q�s�@��mً�`�/t�ڑƮa�M`��~����W��ڏT�o��V��B�E�|�]ȯ�ZY����v�`����8��8t=�Jv��޹���V7�d� ��#{�~�y�:ィ31	6u6 ��Oh��i���������N@�D9Fp���\#���Mf(Y�Fm�gXY���mjG���f
*q�ҟ���%�tU����Y���ȕ^T}'���zE�[�Ծ�y�i�%5�V�1_���Cs�?{���� 3e�,9 �\#��m�~N RwB�"�	HI��|����h\�̌��y�2&�Ha�I����7�ñ�'H��%���%߼�L�JijIV�% ���7ha��8K0����(����N�C,Â��D14�7 �!��lL�\��~]��R[m��膌z9��4Zh2��su��vJ���.4�z��e���-[j֫4�� ������9�A����f&d!��6F6�SH��C�z��˙���g��@����=hC�$*j��v5����5 �Z�U���:�i��:%tG�������ZmF2ך&9���:���{ˌ��z~nd���>����ĩ�������|�p8��q��Բ�Zʧ���z@xg��M3T�y��Y��P=����CB�*�`-���#A�D�ט�_���{�zsg��\ ���N��]���gXk#���AS\�A=��1$��_�G/�=&S����ݻ+|Knݺ%��ȑ��k��n꽶�@�#W����f�|��,j�Z_��9��ŤrϞ~�U�$�(�_�N΁J9�^�W��X�=�mN�RD&4�^��^~�]����̟8q����s�v�;�=���>"����c�C��o,���劔ヤ�U����Ǐ��_�`h���-\ь���;T����*�ыQ��&�k���'�ZR$][��gw�;�k?���h+B���YX�=�[g7�Ԡn�EA�����0H���r�C���R�3Z���F��8؏���uPY#4F�b}�#�aG��{�'E8B��(\!4 �Ue2"Ǿ���&)�"֗�y�wZ��At��Kj�>�h�?ϋ��)R�Y�<�`#Ȳ �(���g���j��
M%�0�|t}'��n�D�i����+�p<�}��҃{w���յCIƛ��4$�:�r\�B���׏�?����p��p��f}g<�>а�G�n��'���(���NBP��nǛQn���eE���{�J�Q=nj�%�Q��j⾤�����BiQ��zA�I*u=�L�Ӟ��`��T�f�A���ؘ�$%��G ���)9u�)Ow�4�׵��9�(_~�9f;@�2���H��6�Iaf\@�$��)q�g�sв��n�m}v�"�'8��f�(5�ԧ�!��"pԥ���$���'�����(��w�%s�^%�1�(055�bgu'jdg%�����?G�d�`��B�A����2"�}���f���sfX�V)�}�VG�v�t�$EqH>��H���fۑ��$�>�l�l�����:ӎ	�`6z�S���`�@\�7v�zz�
L1M���
�s��6D��h�1�(��3�M��}�P��Me6��b���*%�]�L\f�,H�cаFq�k�����q����X[L��%������c���ʐ +��679�pїh�pk`�;���E�p�I�
`6�d���妨M�Hg����ލ�7_|�9�6�i������n^���{�\�XC(#˄���*���(7�U#�q��[��nӰ�'M������ە�g�X��:��i2��]���ޑ����2�ptp�a��KYކ���'<�J��}Vy����_��T�{��%��O"��~�%��9_>;ұ�a��~������쉮heܵ e_���`���jb���
�[�`N<��9�Om���c0\�5���PN��eP5Ijc0�����A	.���sKe "�{�^�vDA6�ܺtiQM�%G��G�*/B�%��ߙ�@T��y��$��"N*<8a_�*��;P�&����H�:JոE�@�q���߶o���s�O��/y<���`��ݛw�쫡�iVZ�j�c_��=L�%X�Л���V����)!�G�#��,��(�"(@��h�N %8唭 Z�*�V�~�?��S�U�՛z�wRʚ��>tA�!W�`8ir�N�G,��Z�g�R��O�����f���3�Q�2b] @�:�C�B�k���(	�a#� �4�?b����Tv�7I��ȵ�� ��{��+���s�[`Q��dWǎ�Q�Kˀ3R��}f�@�B�N�.����5�[e,{g��4���m�i�D�Rq���`����t�9<���W�C�6s�`!p��*��0V6�l���G y�h������Y8�,��]ɫ���9�<�w�e��IY:tT6�7ܸO^�6ÉYa�c1�8cn�{m�*A1�f�=��e(.�Í�4@i`3θ���I�"@��$j�����=)-�0o�5 �Y�G0����ي���u���VH.��5��ٓB�s��˶^��b��~���{؟*@ � ��ؼ$W�Iw��}Y�s�]��� ��d&����>P�[���?�chٜ���(5��>4��:��� �(�l�G[���L��f�*T $�-��:�'�PE/gYڂMa�4�BǇ>uN��&������K_}Qi���3�o˭������Ʌ���9�|�h&ϑ,��LVW�-�f���?��)2��6)���ޑw�ݤX��Ɩ�?w��o=�3���������Hg�Z?��U��Z�*�_�6B�3 Y��T@�����*/��E������#���f�u�d� ����t�	�(]��iغ�8G�s>��|�����L^�w�jl�-OTL�a��8�ƴ;b��L���\�y6&�A)&n�����ۜc�O�U��A��a`�A0��ո|��m.����� �1𒟝D���
wn��c��Ώ��Q?bB
Ǎ��Ŝk~�p��:�
�z�=ҵ������T�}��K��C��]���`0S'�Ԍ4u17 �P�Wk5%hZ��F60�<|��iJ�r�hc�0�F�LiQytV��� ���{/.,��5=;c$,Eq�Z�����N>���ݭ�����A{t����o�m��O�{��/V5����BU��Y�Z�ÂJQ��H{����F����������v$TG��ۢ@��yi�>�p��:���sY�wJz��2�F���0:���m���`��L"�sB���26 ��Pm�1���,��3�2>$�6�SK"cj��	��"\'Ɛ���6+�����͎��dmu@iJ8sP�n�l���
I<�i����ôZ��}$T��s&W4���z@�;1�`�5+ޤq(ܿ�q������8 ]n2p����U ��t�6;����7��#��+�9���3�{>tL��������BU��Y��鿻[��g��u��/16���F|O�zCW��ha!�笜��1*A�ް<��vr�>ȡQ,	Y}���i]�
dk5hAv��k�"��zn�%l9(���N�<7:]~��`ǰ�!�a����~W65 �s�>(p����3��k�����,��E�!١u����gO�K_yQ�f8��W���;���,��M�D�������2u�P���  �y�~��!�Ǵ�k��ʌ�)vΝ;��Ӑ��>��Ğ�~�.i���������~�>t�
�\L���7[�<uR��,���M����K�jE�ӐDE�}�5���u�Ux������uy5B�B�lI���N㊵)q�����a5��l���L{���2�_��*���&b,yC��}��"�����X{�6+4f���'(�L��kd��~ًgG���re�f��[!�Y:�qe r�a�2��?��u��0幕|	NC!v<�$�b�3���
Y�B�Z��&����0=���V�Ň��82��2;;�|�t��th~^j������b����Y�!FO� L����㠎���0S�RIF���`=%V��^A�ȱc\�� ��k ���C�97�湶����//����]���B\mh�|V�����o�f��,F�t�/�H�eJ�}0�5b����C���%L�n[��� �k}�4��d׸f��5L��iW�MG˱��4��@G���5�aSҚ��Y�$������2'*�@)8wdDI�2M1��)uđs�9���*�pL���6>�4(��ݑ�~&{z�[�1�YH�����@1jjZf4 z��m�j�,��PY � p�����qe�Ǡ���.-Y��c[ޏ��rC�R���1����3�ܯ��
i�u��I]�1q
�xAd"d����5r�< �q2��3�\{"t���ͤ�N���g�O�q*8�Ԣ~�"Y�b��vQL<�F�+Ȱ&(��`�Jg߰ފǙx�SR�z��_�ٿ�=u��؏�qK��C@�2y�l���$�Y��,׷-\�c�5��$�� TK����db�eg�f�<EslR�b�|��ș��48���֦\�zE���rT�u����k�����c�I�N��FÄNP��yG��<����k���@�5:��&$L�dSC[a��@A���5}��D�!���]�y=zX��XQC�I��Nq��5�_۔D���׮Kx㦘���H�������|��f��6���S�z�x^����T�Ec��5؁}�1mNG����7bP!Aϙ�)�¾~΂�p��̰d3̛�����б��UÉ�
J�G�O��`��ֆ{擸�q��r��r��/eL�b��2���������m�~ȳ|�n����e�9�����ǳ�+�T��hbc{G��ėB�Y"�s�!*/,�`�����>��ǵ��A;�(:r=,��C��I���h�׾����j/ݻ�ݖ�T$��eW���d��\�ey�%
;�����,:�mfu��M��:r\j�D�e�Y�vw����Q>����nY�^�YZ��*�e�X<#:Qd(�n*���x �liB����g����Mi��Y䭟��S����{�C�I+6/����Ȃ"�s'va����P`�+\9\�aTc�,��(��Z<7}�N[����(@S�l��,��b-�:(/Q��ە3������	��OP��=�\*��{2K�ܜ��|aB��F���@�?bo��iB�4M-[��5�ː�1@���ў! �X��?+��6~��-�j�G�H�K �?ÔU��s�j��5�f��]f�6Rd$�3�7�U>c �"2�Y)ְ��{fm�8��G���$^�gr�0� ����٢�1�~zAV�5��[w�Ӂq�9ֶ��c�n��M��c��KC9�̌Ρ�sw�,�Binc��z��r�"�B�I|���i����W_���>q\�>������ۗޤ�+Z�D�Op�{�����2��R�>5��z3$��x�,}?_�B��K_�Gr�������4Ѐ3�����vMb-�<e[���S�N���4�W�/_���oɉ�%��]�����	LO��|7�;r��-sS-������Ox�]�%�ֿ���</A��F������,�.]b`�s�9��F����5�w��l<�+�n�zl�麏1���#�xEB#����ᰒ�o�L�ߊX����V����dF8Oi��Ag�r4�q��=ȹi���L��Ɂn"�հ����'�u�%�.�B�|�QrHޑ�� ��C�c�jM4��0����},�(E��t�8']�`�`˝(�07FO;�r_:��O�����I���$�+��cp�#�u�Ӈ��p�7�SH�)p`��S���(�֩��R��7#DV'3`��z�@k� ͒����uF���V茾�nt��,q�B���A1�O�@�ǖf�MͶ{Ֆ��~(��D��:�Xo��C+DtV㌠�k~(�o]'X�ޜq��t����f#����,�
p�xH(�1���֐�V
A� 2�3�s�#����s������W�{�}f���������$ڀsG6��G���� ��sg�0��ӌYCO�s3M���z��\F���d��h:퐭�<l��������Tǟ�=	�����cF,��?����d��B5�;j��
ZD�s�ݬm�IP��_#ʁ(��h\0r(|f�9�q<f!\Ϲ���?E����W��O����3Y��#�O˦뻻7R�-�0��0���;�q�W53d&h�d��y��*��u�� `����V�C���%M����:;:a���ڭZX�e��� �j�ک�Vv��AVf�>G�T;��_8$��(t*Z�e�x��U����2����!��A�! �v�J���L������&�^=-5J�U�T�kM9���=s��;0������~�Ր��e�x�qU3ȹ�L�,<v�
�o��s�d�?�[F�k�nYl�1�@��Q�������.�)ͤ���̨�}�K_$�Rgu��+�ё������^�^C��ڕ��z�I�j6���db|�5[�ʕk7�h�X	�� 1r����U0Hm��Vi�˛����g�&�N��1:������h��z/D�Հ��İ�O{P��W���~Wu_�R����@B�1=�GW�����������(*:A0�b�L�[���� V�a��O�Y��v��fFye�r'sI ��=�i�Ja�UӨ�����(*AV��VM��F)	��W�F�Iutq��:�F@nV��ԛ�(m�s�>��? �
�Bm�B�xn(~f�O�zo��u]'���u�н��.A��(t3��٣�z��A���{�����|�3�4 ��(����1u��@�fe�^u"e�D8[*�B�������;d)Vn�r
���s�&O�r�����"k�6\+�?�C��J��d�ϤD�SIG�pG�|����E�]Y��ԙ�2��捫�\Q9�ZUG^�f�4�t�ƈ@u�f1���H�Ap����<g����AN�b@��c][]%��S'H���Y�����{�[�q���o\�)۳34P@�~|�cn�9 Џ�q ��t��X��h���Z�B�>c�?�!��slgu���+�Ge�3�X�g�rx�c.���U�P�L�g�H��R@�M��s���\8w^jCֶ��G?�� � e�h)�6�qY�F��w�׍?�q���47���-�>�x,+J��f�� ���ٗ��>�!�����̌R�һ�É����t�pA� a�>�:��j��<���f��z_��Ʈ��7J���
J��q�����ht��d���i`�1�WJ�jH�1��YJ�"�R/��"�=O���tg�6r���P�+������!U�R�������gu���x�w�����C/|���P�Ԁ�x�ݷ9�`�Ԇfo6�%��;/ުȃ���V��?ޕT'[:�\i1�E;��a4��wok�~���3���>y���;�!��I4�2 ��s�^w~(�>������<{���j�t�������T���ٕ���iu���;�c�>dl�Y�"b�����"%O>��D��,����U���0���}�ߦ �?Z���Y�`K�R���Uvu�	�-�8�'��׋��������X�#��ڂ�O�W|�[��'���q#�?�c���x���/����������E[�f��$��	4"	0G� %��u���z��Տ>|�|B��á�ZIv ^X�wD�ҏ�����L�s��m�	%l���P�1��� K���������?xd��0�c�� �[��V2�!j�7���?��4Ԑ�<�o\dyyog��V�^������D*ͺ�-�LxVZS�כ��3�	;���Ao4*H*.gdِ�� }�&5"������=y��7���#2ۊ���3��o~S�]�JjN�s�5�g��YZ�c�A�O}���Mf��V��x�����Ц�K�Ws�X��`��i�;�s����Z6���5fT&�׹�fUǗ4�ɥ6ؕ��i>ۅ�i����NI8�� YlM�7��os������>ؐ�7?�a�e��D����HfWv�k%s�+�dm�������d���{qNxhY�K��l;$	O6�̒*����D�"R�VFK@�$+㜍4���2Ώ}K`П��\����QjΥp�cT�g�����	�����N&�x�������O��K�@O���M�Qw���I��k~ϗ��k�=�.�X,<R�z��3^7F�p�'��`O=$'����7�Yn~x��9���Qb�������)�z����ۨ�&erj�{�k+N�u��c��5�`�m,�I?pn5��O��wtn��s��m+�0R ȧ\�{�[	���>��g�ܹ��ݿ�����op
��o�[�'g.<�??'�޽"�4�g���J��2�� Ј6ҥ��^LT���-��Y�$�q8�sA�9�4�"����}B"��������1ɐ�Q��`T�4��?�����y�'�_Ώ~���'!�8:�KWo�H��̝S��Z�C'Z�(��k��*e��cɜI�G18�����d��� W�1���GT�Q�sAX���s:
i��S���&���4�T�R��n,/�3�z�?*zFz]7�a�R��<�VQF�bT
0(�j��r����YJeBu.p�hP���N�����a��K�}FV�}B�fU���/ȗ��e��+/3��&��Jλ�]��{��e׺?��l�����<����e__���h\}���+�r���A�M�_W���&�"���5!�X0��I�:��t�4#�k��̼4�g�Qf���M �H��W�����3O��X����`�
��R��L��(;O{�V���Z�I��Ɨ�c��*T�F��=�=7i�Q�9����B(m����Ι��֢����/��#�'h�W��Ni����z�`>����P��:{���{��qLy�G�Jyބ�p�� %�̏�w��6@N�3�$"b�<�@:��u���P5����Q4'n�ܐ���!#���6��<�N�j��="�91�?j���:<�Ad���mr��Ȟ���&Kʑ�L=�>����Hꉭ@8��z�>P�i ��03=�*�.fށa&�;"Ο���1 ���K%Ǻ��<ӵ�;�K���r����}�j�J�o�����˯��ֶ��pޑhY&�6&���14���J��t���=��^�q��tL�����x//�
�r���P/�F��	�͒5�OT��y�t������B�ǧ�/w<�.:�i�JT!�I[[���_�)E��y��F��q4Q�+d���9-;t1�9�BDڏ���A?��4�0��廙�,c��	hߞ:��l�X:��lh�VM��ڔtv�5�d��!9}�̬���|�Ѫ������+@����!ٺ�,�U�@2ɋ:h��C�;!�&������>uB��1����{����������W��ex��a(��$a�0��^K5�I�ըX��۶���������B��{j��#7n�IRk�T%����?�uS�V����{��sSri�-����=t�4���<���o��q�k`s��-y��׬h$�EC�z�U90(96Ofc�>���A�U�Y1�,�~���eR#A��Y8h"ą�p<�z#���Q��-BVR@@S��kȉ8�a��
��5md���L�of��<G� �A��(O��'��n����Z��a.#�Yr�����"g�c
��y��g�s����V��x=v����K`�{�����5't6�����
�F%��E9s���L(��pn���׎�r��66q���7��8E��{�_as���94/�{��և��N��0�:�V_��%3��N�:'�s������&�td<��@09�4u�x���No�@C\���;����U�?���Vl��0N�%>�A��F��g�a��� `2���u���}$�#0L4�A�2��BO�Q�&΃����ج$�(M��t��$Z����D���8��Gw����	 2-cj#��u�9��)�B1� �zo�8��Łh�ئ�:r�G��a�Ǩ!�h����Q�L#td�7ʰ��!U�*���� -��k�0��h5�饺:vJfW��v��Y��_�(okv^�(���U�C������͏"�a,
s֚9�,��eMo����;ߑ�VS��7�.5�@�.\�?��?f��7ߐ����$��;��`/5����]5t�qK�k�8���<��~|jwХ���	H{��T`��npT�-�����g��N=.�;�R�}��fLUY�]�c��y}�s_��_���9�΍��������af�p��q=?�<;��N�g`02�1�%�t��Y32b��>��3
������A�V	HP�o�c�sS�rԦ w�t����c�Q����h��׆�I���"�x�b��~�a����~�ꀸvA�WU��L.��S\_T�2���S�+�Kĵ21�3��>i�>=�&0���s�n/�]�� ��u7�M��3Osk�w�}��� 1
�d�!��f�r;���bP�	�SsU��,v)J������D��v�UG���M�ԏ��(Fږ�����5��ρe@Ђ@y���٨����)O�:����˗Y���?$_�����|��Fn�-��Ɖ�|T�� �G���5&2W(�ܾ�>�{���g����u>hb�E�{gPl#k����kVa����������Ď�'�B��mV�_�Kxe�m|ܘeV��K�ސ�2F�
���s�41J%/4A������D��<�z��oL5@�H�F� ��ƴf�����TkV�:6e�ʙ�%�F�d7�e�������Y}M"��;�������{r��}�QcUiV��Q��fM����#3j�|0����k4��"�ń�2Wȷ���r��qy��Y�v��_}I.�c���J�]y_��� ���N�M�a���r��k	��PW���(� �g���DT_9���Y\�!M	�t*�i��M���b������}�i��k��ưW�_~^>����Y��^��7���|W^��kj�)e���#xh�Z�0J�8O��e�v�HQ8�`��ǁ���T�j�]�'�0�*�X=���:O��X#�5:��e�s���T�Vf�6Ah� Nժu�f��
�r�cn�]����&��/(���$'�@9�o��1
C���8<�;	���>�7~�w�lVLxnG��#��.�G��	��M�Xᾳ����;T+��124:N0�y'TC��^+�Ľ#�Y�8���ck�M�;?#�b&ޡ{�+E��mu�ݵ�f��ѦѤ������9�&���=�Թ������� ��x����G�Yu?}萼�A��=G�z �0��Rm��G��α8_YvMׂ����P���%���Ev����.�hx߲����:AU�8ab�9��2�~�'�:C�(�雘�e�
d�?=>���9�qJ�p.ʟ ��F\�N���1�Mm,����E�ހ�E�R%�=CG��z0�36բ�|���TW�(�C��k`��D�-2���~[z�>�vZ��l��}_�85-��#'ɺ���ѧ���f����v{_�4�F�wv��	10��y�4Xt�H�����Gϧ��w������_���/��ET�dvnA~���=�ݍ-"�˺�"�$[�~4��Ч��r��+,��������R����q]�E�B^�կ��#�l�Z2 �
��3=3'��2�?~T�}�554�4j-�!k ��'��ݗ ���J^}��,��I,[��*f��j�,��0=p:Z�9��������x��x�Nv���%q
�i��[S����2KCV:�n�Q��zq�T	���� B��p��'}k^Rؒ`8u\GVV�ƇW(U��t�Ҟ��•V�fe"�+*�#��:#�܂���Cs'��x���('T
��8��@�����~�7_�?�BGE+EYe�B9�0(��"���E�*����al=4A �Y8�v�FQG0��d�F�o���9ZؐH�%�I���2r�����E�)CCK(�;�:���z���y]�΍��$%fE|��{jjrA�,f�{��8'��굛�}����ɣG���h��}���#��W�΃'1nW��ڀ���v� e�c,�پ��:��y΀��[���d��{����<����r$�F3N�$���X�G�Zyd���q�x,(w�����:ّ�������MF�Grp�����(�و�#b�#����9������٣(	<���̴nژ	� 0۱���Ew�fQ���lt�)$�r}���R�C�@�5ͯ)�R�iJF�1q!P�Я�8[��TC)���q�kbN7�������B����o�;���U>����jrb�&ёc�rh���<t>G�`��C8��^WsqY^~�-bz����=0^�!��tH^��oRd���b�Z � � &40�>~��4����%i���+�J��dc����ٿ�s��^a�������9N �D����{�i�G{���P�LGD��ȲF�-�� �s�$���9J��y3�S����AD"�Ξ�qt��{������3zM�N��Q���H-�Y&�}��U)b���"�FV��cZ��k~Z��)ه,��z�)��>�Q�$d;�k�[a���8B�ٶ�F����I�zs� r��<�k��F�<:����3�D��98�����(<�C�4��Xܤ�ˑe�^rp�C=��VEX`�j��z>�Ժ��(�"�לN|_��k�ޕ��l\ ��~����5�̸�c/��4H>�4�鲱_�X`8~����ST�2	��<`�c����a`�su}�v�^q$XS��]��3H��x8"ix,m�k�^���6�.��}r�˂Qư*I#���>ϘR��1j�lT����,�o���|1bJ�sـ��Q�N�l&�r�Q�%瀯V5�������̹��άmn����N�xhg$J� a��l�?����'C�	��3���0yhЏK0Z�}�3(��1UV'����@��v:�X�1	ô����]J�����?�B{�*a�& ���}R��W���\�wbr>4GӃ@T/}k��Эu0`�5��3�Gy�N!�Fy�N�����Ԉ�����?~U�W���|�������n�2�M���0��ۨ4p�:�#��x�)��'oaNO�:7�Q��9t��l�C���ο� ���{sڤ���Óo���4� ��{��w����\}�C��B���7��廙k�>64���F�mM�sT��_����]0(�����b��\���g⇪�ݝ��&����29s��LO5dgk�e@���
���Z��+���qr�<���I�bq���݂�Eh�)�'8�a0���w{ӹG;dK$"��Af�x�Ldx�zj<w2�~�����_R���</��張�R3n0k8[���E��F*` ����&Kב+��@ c�mۯ��I.�3�b���ʱ�363�yb���Xr���lN�J�Y�w[���C�|Ey	�sU�	T�Gy��)�u�IYQ"�Tp�r �g��F����ӨUda<ިBB
f<g�P�N"�P��]:��W/xo���e��U�>�q �j�����O�-��X���A�W�,����l_i����YK�5ˇ�Ȭ-m�{=]��3{���r[�&��N�#ᧀ��p<����\������]$�'�Z�<�����w�Ȋ� �z���G����V5S�}��ٿnF�M�#�|�0�iV��auK�n�+�ņ��2�3wc"׈�D�ѭ3E���`�p�Y[8��i�l}�|�Q6�w�m��^��ܺyE�x�'��ٳ2Ӭ1p �.+
7h���N�$��E�}��vG.����H=��z���U�5������k�&A�e�e�O!�Lq������qŲ*��ekm]�޾#��u�O?.��i�B�T�^�ݖǭ���ڂdN �D)ˣ[�q+���9�"��=���s<�՗,5�95��K�r���l��˽�7t}�m�+6�U�	���egw�8��4�]׸t��\i�g��}�k�q����G��$T ر�3��c�F��8�A�"���O,�B��6"}�o��YX��b`#f�y��������es�B�4���#7��cm�y� ���=��pvo�L�����3�t�%��a%�x�/�u�y�I��m|`1����� \_y�Q��2=���	ܻ��mf�B�r���<7|d�k
�	�(*����ѿȾ�@/s�5��pZ&4�*G8��6��Ɇl�p��T��{�G_�_W}A����L5��RB1���ٿ�63�ֹ�|Zr�������^@��B��Һ12�{�>:-���_���#}m��n�G�3,�<� :�]�W����d�ŲnLG̅�����;*[�Z����� ]D��1d���5� �a1b���i]C� U �0�������KvI{p�gzcגJ>긼g&i(t�d�J���ʮ:��֤c��5�GJ-v��Չ�o��@#w�hw�ž[൶C:Ɏ����R�
�-(��|�@ˋ-�������f�w$�[��S��G��E���;T��ސ��0C�O{=����B]|X,�|�U�� 
����]����ݻ���)�E��%��5:.G�$.k4u��e��e�Pq&�	J� ���[P�v�6����Lsk�༼$>�C�5�h�Q�	�h��~X}��7�Ӷ*�{W��
�������'��M��ysW4����#p 3��@\U�N��1�UCp8����{t�Yq�:~�����^<\U��4x��pf�Ϡ�K�T�ܾ/�]���|]�љO��= ����M��m=�`,��ɧw�G��>x��z$�J��>C\�'cB&?����6W��{�ݫ�����@u�D���
�$pT�e_^?��6�����ˡ������YӠ���Vq���a`(d*�����Sh�?����'�H��a����7��g'�sunv���(ɜ��)��e�7�@gށMiH=^Rt 
�ˍ범0vѿ���A�Ȫ�cL-a�DzoR��Zj�>��Sr����ǫ'U���F+���'�9L��b<��~���qA�~��{��{�3���pY��Q ������Y^�&t�9*c�f�&G[Kr���~��ڦz�P�����1(Ib��;��K�W?~Y��T{#y���r���`��z�q������l	 !��4�By#��0� K��
�Pڮ�}p��U��@ՙ|p�Y� J��V���\-l����Q�h�蓈��=H��_��\o�6���B}�r��Ǭ����y"n��pٯQK�"�!�S��-G["��!9��>�n�z��t~�S�2x��'p	���}��s�)6�g�r��/��k�
�l]	?5�[�e��9� 19�1-2Eƕ� Ka�Ө\-��\Xl�%����\L�S�@�,?�v��D��2`�	Ԭ�L�ρ �Ӂ�7��E��bwf�M�z����E�r�LT�|���F���1I�.�;�)��ad����}��(�p<A;9�6�y�y ����(�f5���e8&*����C�k쑍����á�P�������}YǤ�4xLn�_���z>|�q�,ʲ�����|��^���yX2h9Dl�4%�0�2��0��Q,G{���M9r���Qn� �
��>�ycC7c~8/����:�_{�E�ڋ�SV��)��&Fm��X��:���	��.�^�>�o�8�����Sg��ں<���sL DI���J-����!����C�mE,'BB�]����)�� �!�[�:����h1�j��_���!�X5��+Z��
��1�~{jҭ!hU��Uw���$��,�pMtSe���m��"�� �Q����3��F']ٞjt���N�����8��|/�܁E���k_.h�X��	J(a�S�iƄ���Ӱ�17�@d� ����G=� �vM�4�7[u�:��eҩ��h�<8B���;��1	A���~�e�c�&����É*��>����O�i��Q�!��jb�a/�3�7&�j�'�h���������C�G��}zXS<p�깫zd�,f2��� d8*��X�qe��p��̍:����a=B�D���@Χ�LkS� �Y�/~�!?��zn�jXm�I�u���Ȣ�ևQ�>p���ݩ�G���[������u�U��H��|z|���r��/J��Gu�_�I$1��NK�'Տ��s�����15d�Ÿ�M��I��ڒ������BQ�a�x+�%�����BK�'�#T������;��'�\�+�N���~Ag�E�\(D�ƙ�\$�2�� ��U�{bqAf��n!K�@��T��!�sM��Z��}�ey��:�ew�E�h=26(���a\�'�|� �]U�^w ��u��lo��c�H�d(.Av�GH/���'��(s�]B4|F*Ҕ�k`�����k��~P%���ΎLU��v$W|�/U�0��e1�����@�'�53
2NT(|F�u�U�BV!��t���:��Hh�\q�M�[�9���{H=X��Y�2��
�Ϭ�b����2*�c}r��;�~jF8�X����%�Hv:[�
.�.  ��IDATX]p�p\T4�O8>�g7�:T��HQ[����C�B���_�BC�O�8~�g�
)�n��"^k:p��w�zw��G0��|}�e�|z��y��V8圲Y
$��,u�(�BR���>!�p�B�QƇK�lq���;��L�a�w�����<�H9�FB�އj!\3���^Ϝ=�4SfUn��������"f��$Ǉ!H���8��Jn2�@���	��\�+WĂ�,�x�>y���>8��A0f����]Y[�(�xv�%U���b6�BZTol�����H��Y:-	ܘ��5[R"xʜ�Ѩ�'��b܇�e�b,P��U��9f�iUkqV�֋��FQ�Q�ђZ�)U����H�`,�3Q�~�H&��]�#<(�Ӷ�uq�����@��bFMg�9]��@��n�~�L��=%�ܪ>Z�<,7�S C'6���"�8#��W��A�\|ňX��s{�-����F��~�@ϣ�Yĝ�	��L�����r��Y9v��3?W�\K >��1-0 ����qp�&PB=攜?J���?����˟��w������u��t�ץ��	KԹ MP_�p�(je�p����.�p �<��'�"�I�"S"苡��Z���:�!2��3��2dh�o�yr�`вq��g�f{���NW�������n�+$r�u����C5�`��6G�c5�x�,�B�NY,�pQ�\2�J����'����5�\��(e�'��U��Ul���g�B�x��R6�,숑)b0�r2{��@a 8ҞB�͓���00^��$�@o�뚙�s���we�Q�Z2Aǰp$`ӳ�Ȝ���9۟K6�'�Ӳb��cRz��C����{3�QI`{��bϪbUu�QU���	�V@*���0;��G��QdYy�[ev��k�^7x��
�����w��p�_� ����ܑɳ����X<�w���Ǹ���>8_LtP��U�yF�`�Ba��ʀ�&�*�t��������}��,�Uq`�������(Xl�	��1�̌�k�;T�qc��%:���aD	�v0��&Y�f����iŵ �S]�9Njq�ht8�ُ�s�>q��T`<��k�>�-�O�f>�,���D�h`y)7mL�7��,_ifج�d�������{�� �
�8�PB��Wg	�#��tv�I�ݻ+�����P�ˆ��_oT�6���#j���:���w����89���y�&̷�W���3��wU3�W^yE^��Od��UdqeY6�v�13E@��~�=��M5F�ƃ#]d��tGD��}�K����&�s-�4hh6���qY�sCP�����L#@���Z&b>��F�klVAX�|a��w���=�&�'��5�R�{�<d�`Y? Ш0%0�:� "ɭ
c(a��7�4�TP�����'�C䣒	G�D1ǧ�� *o�R6�t�B%4�6(�
#�+^�&e�9��F��fQ9&"2"���5)�	��<G�XIf����,�k���B��I65�h;����:`fY��Q���4�_����P���r:θ�8�1�m�`�/;TV5����j���M�s�i����4� !@޿Zݑ̌�qq�$4�/Sj�^V���8�)��D���tt�+5k� �hI�b���ސ�ԝ�]�d��S�?|$��=��,b��1Ք���Y�j5����v{gO>�w�cat��������g�}�I��o�-.�9�Fײ���LY�t�<'��zL����3S���̖%zs���CZ�YmO�ޢ��P��L�s���;t����;����&h�=��،y&A8����-+�U�0�^C��ޟ����ְ~�]�����O�M��d?$(�%cuu8 �0]�0jA4��FG3f�`Ik�3A����j��`����ɑ�+]�Ȇh� z�0�}�cR+�?������ל�CN]�n�`�exoMT�e)q���z�PD�5Z�IC"�[B�R�p�4 :�s�z�m��@b��h��4d_#��5%{�[�T#������.W�<���e
�LMV�`(a��i����y&u��1��^���醼��s��0#k��jPs[6ܧ� J���f����l`�Xf"4+$�4��.hW{#5���K
�<�|�9�T�`6i��s�SHǒ�-#B����Ha5e[���8��������2�[0���b$�\@�l2p�֫]���w0�ZK��ȁ��r��ӥ�72Ǚ�9h�/=*Alq��	�b�l�o9��,=�I� ���9�#�_�����2St�d$�Q�������p쩣þ�v��������3g�{���g��4s������@_ہ�.�c��r�u�q�tM%.0���a��54L�{�e��U'p��V]F2� �B�gZ��������Ml�D�Q׀Aϕ���K��ǯ�I\	�~�Lzv���&!Ln�d���3����I&8_�Hz��]�Y=��D�
O��Z�kiTc�K�ò%�us
g�T�O�'|<��rR?[r���I\}m��#&Х��8&��|Y�ڜ�o�ܜ�3����b���Q�YA�I(P�p���Β%5D�h���NzZ��҂,���;0"�v�����Ո*$p���l\@�cͨ��Df�P7ALc��c���G��=F���J�T�|�F��wϞ5��:Qn|P�����C��C�w��DT$RA�N�"����&�ܗ��9뫩����.�!�|}�^h4��c�B��w���'�߃�kj֏ި8r�,3���!"�~[��{ي�������'��?�$ݘ�LxQ�֏R����.h�"�l�`%-���QS�{�6GM3�^�����#���Xh��{�l��t^�j<���ƶ��v������N�7닊�Ϣ���}oܸ!���!+'�թ/�$�8���1E�j�����<M����#��9w��EJ��?!�M���ن��-���p�y8r����t���,�����61&9�ť�$�8"����ԱU�\!Hr���<����ruS�Ë�r��Q7
f�\-�;'W&3	WWky�ph�S�Mڐ�����I<e��n4.�����a��{`y��ڇ[�w��g@2�W�s������`-t����������9y��K������N��'��ӧOS+�7ߔ��}�ƭ6�5$8��7vB?.��cj����e�P�~��S �#9Ϩ,���	ɂ@~T	2"���3����O��������1����"��e��QH	`3���ݹ��CK[d��D�r�(���eƏ8��2�ǈ�8�����=�8�����Ӡ/��F"�`���:�S�P�3r��Q9�?_�L{N�:ʘ�aDD��֭;��������F�=i����p��U
:�)�����Ȳ3�$��0JÅ���A���w�lb8�u�G�eƍt�l�z�)y�+̌[-����4Q1��f$��|�on�J��I�s0�ᚡ^;2+j�gf���mʌ��c�e��/�nߗ�n�]ͤ�5����:wu���RP'�S:&A�`X�ti��|�6x���^g���mo��˗�>)=��5 �z�Ӡ�{��{��IU�C,�`�V�Շ�ߧ� H5�T l�������.���������p+M�	����7��7���n��ep5�]1]��l[����@� ��Fmu�T��$�E� s��pXM?��Ѻ[Y�ęT5���8���͏>�3�CvY���&��>"�K�������]l����6��`f�GP̋�яld�Z�/���G����PE�1eq��Qr��/.ɡC����=T�/Y�GU!v=pW����յ�����|杘wd)�Y��I���<�}�%o��@�;���{;]Y��"Hp���ȥ���\E��ܛ'��cG˫/�,�ǿ�t����yY�o��o�7����ɓ'姯�v.�&` )���Ą_��h��{�_����������&V�?�I�5_1 h�p#{XC�޺$ih�ydJ�O����Cϳt��.���PA0ч*��^:t�ԹO��f���m���l�Y�QH�g5-�-��8͊i]ݏ�x�z��Fv8Id�~����t�-5F'4{:sxE>��Yu�ꜙ��k�Y�h]Q�xd����o�#o\z��.rr�f'�g�����B�%��>�L�8T��R���	��Đ�ab���H�33dwB�}���e�5[rW����:r��7���n�S�j �������������m3[D6����	Y<�߇��P�;/{Ìd4�k���yR�����A���ܺ��l޻-�jKV�DG^~<��:a42�[tA	G�w�������[��/��_�O���f�{R�ƙ.y�D �$'��$U��"�}I*���H�tkJzz�ȀM�$��!ӧ̪^;P��\�C��7��$aOƲ3���5Z
�����΂�/]�`_���W�fx�[����C�,���X|)F�v����Q��VJ�]��5�<?Wbg��b}{8V"��*p����}��r7��MO�ƁUV�PVo���j0���LL���
6Ad�Î��9�P��N����<!k�|P�BW@ꆐ/c̓��CC�|hT���[^/��{��1�6#���?2y+(�{,���3h`m�κ��ǲ��mR�n�bF�F�z����� �l����!����h��̔loo�Zh𞼩Y����os�B@���}Sd�����f�W�mOΞO��=��1��� ɿ�G5��&�D�����wN���i�GŐ�������p���8���c����u���r�G���z蘱D\V�Qs�+=٧��f���CIh�U)P���F�ˌ�pA�|���^I���IQ�i�a=MK҆�6�!�1��%�sǏ��e����>f�y��c��֬ѡ�=vD��H:�Lo||�J����h��u`�B���J��(%����P�p8�
	uܝ�~�:2����ƭ�Q���g>+/|�y#���_\>$UݘW��@�����!O�9a�M?�Ƈ�Y"KP
�� +\��5CQ��t� 8�˳S�<sF�������������)�[�pĔllnˋ/�(�;�$7�:)��U9�rB��[ߒ˗�[/.4�w���Co��}d�Q�lvT٪�����}6��i�����75EH��s�V��z���bF��
�k{�]�k�񼲾��	�4'�"~�9g_�;�1iZ$6V2�@(��}dr�4��U����ݡW�29]#>8��%3S��GCݕ`��%�n�Gl��\�e^��|����}� H������Yj&ը��*z�N�;��C 8а3�����M[��C���Yn=�4fy��=y�������ѣGYb��>�APL�=}�L௼���o���,Փ�L�e�ԗ�XN;�¿�t��1��}���l#�**��S8�6ڤ NN�zT�"r��6	TX�J�BA���ˆ��VŴ^��ϙ1�7�LL&�pP��Az�\�D� 	�x������u:mi��@��gP���Zi�5�}��Aj6�Q�*Iwy��|��ד^xaTߊ.]�P����jY\݂y�v6S[����y�}��~x,Ҁ���/�����y�?�|F�bG��q�ؗ�� s����Xz�l��� @���n�$�5�$(�;ĕ��݉>:_=� ���e�m��!W#w��;���,��h0�<�5��FE1䌥�#@?}�:�ó�ꠏ�I����b��TM�̆:{(-�E]#�M:�1E�@N9$��կ��ꟳ��[�!'��5���{�áFt�&�@(F�u����}@��A��,�F}J3?�{��aIԠ]�����|x�={�����G�#�?�= ��~F��!+9�,Y�F<'�l�y��\s\��kK���C�@��9_�k�n�>?;#�3-c��D�����ҳ б���@#v%��� -�, �v>"�bȁ�"����I��s�HcA&��r5���%*]X��hP�*Mд��^��GƦWM*4dWKӲg��d�0�4�U��G����I�"��X�@���P�@�����{ڞ"V�����G��.�$���~�F��������a,q��0�U�'���@d�:�$"2v,ņ��
����15 �V�}���$.��J���1���:%�`��� ˮ~���Wt���֞P��k���3�N��d�3�4-�z��E� ��|E�H�&P�6.+�a�
��ԋ�q�����~�J�z��_�;w��\�O�E8��**��y�sY[[g���W�"+KK���7	t�ڛ���_����L\��?8L��i�Ԕ�F�q�G��~655�@bI?�Wv���/ȗ��e9~��ͽ��!������v������akF2��s:!T��U�*y��B��v:�������?��	d�sz/�t���m]�y��AR�v��n����[iV��Zk�x�0��/0��k#�j*��7~�~筋��F����)��4����� I��0��b��,�I��� Mb`��2���kz��0,��5��84��gX�����P��V�s�FC�V�Q"X�?�\��@��;vG�x<%�Bc��C�3�0@2�S�v9Tj�MG[i/)\?�p#�	�(P	^�s� 
	����b���r��<��4��q�H]7Ld� S��&�ĪR�eՃN�@�d/����74b�ʔ��b�|W�t�r�(��/<!G����M�٣��(�cµW�R'���#g�9������1��MU�.�2��l��Fb��1l�GV�ȡEy��~����Ј/�N�Ow6]/�ƞ1ʅ�p��A:d�	#���(���9{��`tEH��nw$GϜ��5�����'�6v��\U��}V/',#�\�O�|d�8�y�����Sհ�Rh�K�\�3飯|E��4^m�5�e*�r�s��Rf�Qf :w�y@���IN9ϔ\�_�������|�5����1Tpp�(a?�Ҫ�c�~���3��/{�$�y]	���gV�������H�~HQ#����b4����bccgB��s#vcccc���*4C�4%2$͐�HI $H86L[ �}y�>������nr6(�1��bwWee>�}מ{�q��(�C~l1�TTK���0���d���c��! 㬳	|$������Xy����:���{e|b����T�8g c��uX4�hY[���A`�JI'	�V�� **�ʐ�4�E/��������YuB;�d�3�DB���q6੡~���k���<�
ٽk�\�r�t�AT˲��@��apט�;�X�V�
�����f����\#_ ������w���R]����YX�Q!i��3��i&[�`I�%������/���ڃI����!�B��}������������g�}~�/��J;�O��@U����i��фR��k�����;w�����ѣ��=�����6O�ͼ �'ח�&75 Gk��1�-�1�	W�'=u��iл'׍�e�ӞW��[?r��|L�'w��߷LN�\�N4�D�3���|���X׏��=����NC�N���Xb��M%Zp�D�\LW2 G�؄2Hݴ� Tr�bf1�o� Ih�ֳ�!T��Q8�����l�l��(�T��_�x���9r������Jz٦���:�\c'U��E�3ow"�ݰr#��	�V@�vZ]�����;���l����ߍ��V�����])��U�!Ի4;��P~�K�@l(����y�a�t�dѓ�憪X6O@K���n�Ary�B�� �s�r��U p0;5��v7���ںޏ��s���9�u�Z'�c�`�cZy�J$�:�����J�@8FǕJ��gT� G\?#A��i6><6�^7���\<n�C���e��x���jeXv��-K+�tVCCy����<��:����wG�wޑ��Y-n �e�� ����1ٵmB�|Uf����tm��KR� {�ɕ%T��ur��{�(�H�2���- -�Xٚ�+j��YXG�I _�e�'���j�:�n��7F=�Xk��ȁCT8Z���U����MHsU��� ��=��H�Ǎ�ƈ� �����}�6�{>r3�8b���K�>kZ\\��:s|���&�Yf��!�ѣ/�<4� ��*��	`@R�0��:VL���r1(J��f���]����F~`�j��0�Yp�L��"P�[w�Y0�\�y���)���^�KV���hG�C��nM����n��Ҋ��=������,��(V`8� ��gdǧ>"�֚l۾Kz�}��s���1Sl¡��GK�#\��S<�r�M��>�-���&��G۬�w7@�ZMuҸo�?��۴s�<������g��g�������.�,���c6�e D�b=�����/��W����Hע!�Q���~�wd��&1p-}ny�)��^�d#G@�͠gdh��`v���@6�/:ҜȴX�1Nz��0� (����+~�'&L2%N�2T)ʪ���~^��$��-��kPo����=�z�f��XY�ک+3��t��o�Y������ȉ#�IL�az=��H�[�8P��K, h�"�\d�pǔ ������2�B��[���%��[HXg���@�Q�eM��X��m}�?0��붺���Y(��A��) �p����J�Y-��]�^A)���s�|�/�"�~��Ԭz�:N��bGe�rO��`�h@�~?��q<�7��7������7o�O]��95�4�V�	��ؽGq���]����j�#��Al�^bF7���\9wNfnܔ��O��G���zG�'�c��F���bl���E�m�����EbT��?2��'-"w'�����%4��e\����Q���r\,��,~=����׿�y��ɑ����{�9v���=�?�����"��q���U�.��Y����xVJcS̆c�"��Z���$Ь-���"�����FJ�R�����[��E<�{<T� N��b�Ԁ��y [����Y�}��N�U��N���Z �ѻ�{����36;l��F*eV:�پ��$�^��DOʢk�*B�%��џ�q |!�DR�~��G	%���0-�߱��&P1�ݽA�ďj5���8�� �Y D�պ�v���1<�%k��崮�j�����l�2=r}.�|2�u�����8k�!�*��3|�h?� '�,�2�iֿy�㲲ִ��t2���b��������ԑ]�1+��~[��\�74��&������٭����f��������!�ؘ���}#�JZ�`2"ͶM=����qB��	��z��2��>�)�ڴ�S����'Ns���C���ĄbStX����ͳz�wmmM�c�<o �Gt������ATA�`$g�\�\��|u�c��,�C`��efc�ւK��ӹ��;4������{趎yX		�Q�!�W
n��a�`�;���XI��Ja1�W�a�ټ����v��p��%$p:t��ɨ�>�{q㊦8��lhU� �Q��U�I�+A_A0t��SF�%^r6�P&�� ~:�Dw��N��!l3逑�e�BW�����z�So�N vd��9��c2��F��ac�v06��TэRA5}�.��B�� ��T��3+W��bT��i�Ѳ,5��I��n�j��|�����p��6Vu��r�^����*&i���QL��R�]�疗�������nJ�lvlrZ6o�~�'�|��/�12�]�-w�37dyI��v@ _�Z��HE�ܼ*��r����`M4�oF!K�KkKjG��y�R!)Fݗ����\0 ���*�@5�g�òda��Z\	�2jǶ��-d��	�9��Ԧ	f�wi�q��	:�_�ܯ�G����+y��{e���j�rE�4 ��I�R�@L�%��YA�u|x���8jɸ��r�>L{Ҩ�i�s�ED��VZ�|
L�Y,6��G �*$�Gg�ڂ����j�(����z��+�������j,��P1��ĳD ��R��gD��K����_��,΃RwŰ�o��NC\4��2Z����O��u�މ��`�N�r���W��(�>%g`�HW&!z�9�t�t���^-j�q%T�K)I��{ƀlX?9��� d7XC����m�k��2s�::����<�_*#��3��}zG���Gd�����X{xhG����]��U��\�C�:a�:�)�m&��h�m�]\������hUvn݂;������`A�r�������ē̹r*�Y��U"��Q� Ϡ�g�+u]߫˫�����V��<���OL��Q�ʱ'�5H���hs��]�Q8�p`0��:j�7M��}����|F��m�p�jW�jC�/*S����u�z}��Ò_[7OK{}��F�,yL����x��M�}B��{簵��7$9�4��$!i��JMAK���ٵ�	P�V�`�"'݋%��g����MD����wA��g�~�����V�eJӦr���K�:<���+C9?Z�8�(���R��6�2��Ž�?/� K���W��Y}��
�� s�f��Lx%����8��Eq��\�w�Q'�e��.�0��9%��*[�7��3�lA"`|z�D���R��4$0��g�`���p��Whr^6G$p����Z��k_��8��~H}���&���4��"FmZm#rz��$�|.w�����������@����R��DZKݰ��>x����ڠ�l}aN��62�Y=��:�:C+5��X�ʅ&��y���5D�)��p���Q1g>��g�F��l`�u���-��Cv1��Dv	��}��[�Ť �X�P��
Y��4������m����zX._����R��N�I��&%}^�E5�j�+CѬ-[V���}��rD���g
򙱩Ii@�hr��A]�S#�Hl5'
#E�b��?V.�g�Bd�
�n�v�������h!�����.�y�-.̫ᮋ�%������7X��麒���� #/_��<��J��jWVVn1P|���#����gE�J_��M��,ʖ�(M����8�@v�	S>�&�Bף���z]e5�C\�	i�l:�9�X�^�$�����Q��cA�R�5��Ł%�Nu��!�pQߧ��J�(���u���ٹ{8ʹX73��ʺ���Y�$,�C��^���yy��I�����ő#w;A�@t��7���σ�b�W`������@�a�TV�W4�Ѡ�[Kl��!sGkB�t�<VkB�.����W��_���P9#Fr�ð_�LS�cL�(����}�˿�y�|�����ȼ�M�%��������=��\�[��ٯ��!ړ�����
H��^�������o#������=�I�y�nU�&R��X���l�P<�o Aj�I������h-\,�
W��������Bʏ oC��؀�A&59+���1aB]'��'���᎞{�I���8M|Ui�f�dOܖ�-]l�-���l}3�
@��ҎU�5�C/��\$xO�![���x���= ^�Dx��W�vzIG?�Zį�z��O�z��>Y�5������^^zu�"�A��pFn�V��¸�#�*X��E�rD�Xf_�=��͘'D�F�>�j���,ʂ#G9��P�X��|fJo�d�]ӻf�y'�YC�d
Q�.�x#�1Ƙ�:�{���D�f��[��եR�mG�q�3�pM�?���ՠ�j���52��eR���V�	�Q��}uR�tHGZ��z��#J�~�'�D(������q̌�d),�֕���#s����jܑ��A�
��f�*@A	�Rk�����gRIG)�6lxR�ݛ/081�L���p�qH�)y��6U4�)b� $DQ����g������w�H�@q��`��-"�A�z����l:�jп��S
*�m��tS�鄳@/<��.���wW��h�B�J�5]S�T����n��\ �GE�ݨ�:��m��=*{�H�t�>
�S3��u���>�O���a>(q����b��p��87�#��>Q�>>:N��><:"���0
����=<R���Ͼ�*�f����n�Y?*6�^45C<w��k"|��0ܦY/Ʊ�'�F�ILVա�:D��gLMofyn}n�\�F܂ʁ�b�=(�u8�2�[�@���k���Srϑ��/1>|��T�ZϞ;���Р,u6����  ?�7P��c�
d���`o�i��G�	��س�<���2�y3'!FJU�t�|��dfq��+���7��ِn��Z`r���ݎU�����"���(�?�<�W=CE�셋���!b[<�kl�$��X�0?�7&��~F9� �15t�Al��_$ ��h+����fKn^�$�:8���@%�d:������0�w���tvr|�?m-��Z�vC��	�����l���R����(a�Yp�p�Y;q��2�Ͳ��4,q��z�mu�-u�L���`A��G�l�f�8T�	�I�*g����@��I�ӽ�W�S*�"Ki�p#H�)��3����+ �h�5z�=��݉d��\V?$�8;��+�f.[xshb����^�i\�{�Ѓ`O��_}i����k[������F���'��0��q�.�ڶY ����P�]�A9ZtZ�I���}0d� x��+�|8y�Sc�BD���)[Y`���$'�d�ےU}�ȌكuJ7O���; QE��Ճ�#�;1�
�O&��ɚn ���C�/�yE�u��4�w��# ���LAN��6��!�2��NAf N��#c.+g�*k $��{F���Cb���L��q��
�*7{�޲ bx�(�z�E:�
�KG4{s�3��b[ ��co�!��'���0X�l�{�DP�*g��(tR����2s٢T��s����
�WKT�m��ʪ�]SbWx��Sc�rϓ�ɓ�?*{wn�3�~�����kD��g $��� ����P���C��\��K/q%z���씫��h��bc�Rǃ��,vfC	͗���~����82�,:8�y{�1˞�2KL�%<��"~�k��Y5	bӀ��9==){vo7�8u�#z�������:��~���
��vc�N�F�`��r��  0_�;ΥCf�U���`v;��B��cG�!�7:�P=
�����d��+��~��}Cѓ����~�A~��a�1�k@1\ˍ��U���!��

�>�@����郶�2S7�����c�6���s�ݜ^A�����$$�c\���c�f�ʑ���B`��:�"��
������ �oM����M7D�| � ����6�&�L�A'�;��ĕ�7���t��ڲ����sx����ɓ\B����ݩ9�Zc`$N�UG�Ϭ�@�gs%�}�Nd��B����>pt��wMn?9;;�����68���箁N��'P۔.-,�����|���ϟ�&�n���_���
p.���7�ާ�߳ׯY��r��
���WW�z�?���kl׏;�3��P'.Dќ�B���nԌFoЩn���3Dméیm�V\�^Ǥ/յ0!xa(,r�JY�%+K�,�&x�����(��F��]	����.��H%�T�j���~�Ȫ��A�:�P3�+TV�*ަ�z�eu~7�j��X!��.Vh\�4�ZWA?YSU
͚��R*QjX7��͞�,-�鳗�Q奡YGi�j�Y��j��&���
���B�5�e���$%��pyĺ8�/Y��?�p�?��l��7<6l�W5Cyf���%��f;�.]���}@�:x��?�`���4��{催jF���0Hn hVج�Q�J)��#��Č��@0S�v{���=mk�C��N�^�̢G�/K�F������>);�LQY��F�ѻ�˓�'���K���7fg�¥�jP��ȡòk�vW�<==Mc��/�;:v=���Y�s�X�^G΢y�+�Y��j��M�>���{���+�Ȑ���%�:đ�{=��^���POt�gI���$�[�[����z�D,�����7��=:���K_�VqZ�����Q�� K�g��J\���gr���d�����k����ޜ����8�Rh�sp�tC��a�S�D��h����wVNG%���u{��������7NH�Փ#�2�,�����2�Y%��n^�*���1޶��B� ���"�'����՜��i�4�߻O�w�,X ��q��|U������˯J���=d�	�!Y �
a���<�,���t� ��-h�S��ܷ{��o�ݜ�*����`��\(J[�,���Y�Ե9���2�Z��9�M񙺓G7�S7F֌B��O�vv��X�s�ޯK�zô& }�FT0�`|�{�2!N\,2Y�{"0٪�H����O.���oq8��3#�	naE��s�g��u�Jut�D��<��B�eY��8o{6�`S���!�{bF3��]��<�y\ȓ�� q,y����lR��i�^4��i=_�uBu�QO]Y
5�\�P�/K�z�T�
�BC�:V{�X\.��Ns���ϯ�<|���O֛�	l�Qu�C9~�M��)��TKe���R��͸g�6i�.q�d�Zb�;�%>55��IY��V��~�{/I���"��}èY�(CY�e�ӓ(H8��1�G����(WF4���1E�C�Q}�!�jhv~��;�O�����:8 �Nbd���NA���Ǐ�f�X�����ʒ~����x�u��0�tcn�����e��1�jp3���G�����'�଴��M&�#���Hq����o� �uU��~����Sy�ߓɑ����*��}��oݾ�����%��_����NM��}�)���?��_S�F����2��օa7 ��=D[���|���Y�q�ߪ�;XZ��˨8|�}x䝻�i���ߛ�4!O<��%ͬ� �B%�\�ӡW5���큮�,]?��U���F��Cx�{�e�vcF�zo��b���Bdzb�������+����^9�U�����7g��k���{
Q��ڼ?&V���*4���Pq�B/9_���?�I�Ϗ9@-
Q��R[J���E]'�9t���Oex\������qyI����Ѷ!��e�i25^|���y����{�%gTp�@��颼|��yy�����oJO�kp��`L����NM�%�D�@�R�%2s�,T5�$�&5�<�=|��]�?dUq۶���c���GǊ�F��C>84@[ ���`��� s���qC~��u�u� �a�d�u�/^��9A�T(I��+g��I�}��������.����_>�3�>|�ѥ��'�q���tڽ=�hUF�<�����g#s�&�rJX0��El��n�<�ƚ.�2	d�_�&�7���i:;D��c̨`YH!�a_N��y�|���g_��r�
A���@#����5h�
Ia���E��FE[�ݗ/G����Ʊz��ͩ��s�o_�y����2�����
PU�Ѹ�k����H����Nk��+V���)e�H�~W+,WG���N�F����w��;���Yi��P�:1��h��Ů�30��O�sܼ�p��pd�r�W�!!�Y�{����܂�޼)W�_d&D�}�yu���J�q����h�ڙS�����^F�0Wy�ԩ>(����e��U��j ��~�Ta	��Y5�h�#SFI��N�:��Ϟ���J�~�ƮOL�����2�ڹs�,޼J��RN�U��5�z�dێ�쭧�/�?�ň�a�tPnͰ��G0�kgsω)���fhD���r��a��t��{��͒eN��f����1���@�z��Z��L��1�=o�}5�gT�z����5 $D�F���g�%��&Q�֭�Y�]_�g�CU� �߻`-��4pC  �J�V ��������*z�~鳟g�<�5��n��:���fϺO�ڷ� 8ɿ���%�՚����,�#�F�U]o)�qϔ�29����^~��  >	��PBG`��m����,.-�u�h�D����l٪AC�"{v�auS
~����&�Bl�`H������v��G�^�3@�ib\�ٚ�z�<��eI�w;	����GL5���o�q[��7y�������}� ���2�	�3�+�UӋ��pO��9��4x�X�ޯ�>��gD?~T���e~g|��c ��}��c0 �>>�%(���{aH�h'�4?�=*����
ۙ�P&�͝�]=�Sr�m�w��t��K��u)�����Pn.�f��S(TL�8ut���E��K)AH�Q�H~e�6G�v��q��#�	؈:J.�����OL�O���x�����ſmo�E�뺐ko��4���ɚdb�\�m�|`�`@����r��=4kh�$�}�Z���"(�q��¹����Ͽ"Wf���Bƴ�� �������1'k�S�U9���Y���ҿcy�="i�DQDg_Z�������5u����<g�evnNN�<��G�%u�I��7��`��&]f�^rR�#�k�{d�7o�\��^�˗����~D9@�ȴf���a+���vD�"ќX �T�hl{(k@7^-��ðep��!��$���� $Fguy�ƭB���	��Ƽ�Lƍ�1�enU�`��2�'��D���`7�3��D�L~���HѠ�I��5��e�Y#�k�@G ri6�Y[�����n ��w�  �Rn�kv7,�ϝ�u���Vz�'��jAl��ݷw�l�ޢ���)�!�[�
�43.�I�E���1
��zbţH�e�F\���/�r�o�����[D0!G��i�k�i ���\[g/]W��A�]r`�nNA�87�%z>Ș�቉I��3�ն��5m�3�,Z��~I��^��Io������)9~�-�ݘ��!J�-��.��������
hw�ځ!b�j#Q$z�kZ���׏������F����:��>�����F&�A�����
�Q�3_5����B��A����'HIM!��'�A�Fbp��J$�!Ԍ@VG�+�S
��9���=u蕇�����/���+�כ���^�)f��٬��n<ƀX��2�zc���F	�X$�6^�԰Q, $d��͹i�t%��|��lid��������c����׽F݌��n�B����0��7Kq��꘷֠�} �fհ,�������C�����r��U�]�0��.k�95d�f���L����m���(���Z+P��+��Q61��w��.����U��q�ojF~��uVM������\RC���P� �,3Ք8� �yKB�oanQ^�l	��Q'�iv����6���ϨTJ��a@6�vs���Ŭ1��������3 ef���uB�{�9ٽuRvo���:7��"u���^�:#��}ZV̒��V�ߜ�#w�� ���r���>�yƕ,ayX�菠e�}D�OO��0Z�k�`��A�~MeY=v�A�'��~�A�w�8��^{�u�K�~��s���A�.�^��1C#�7��=@	������~ܠa���,^�K����p�n�o~n�Ncxt��m[Չ�Hmm�Y=��5k���p�)NW2��-55E��zO��d��[f�"E �8F�0� )@ֿ���0�@�1vњ��y��@�����C��[6k�Q�Gc#|˺N.҃����t,x�;(����SGϞ�b��@e����;�Tpۀ� E�;U�3�T9v�v8it�y��Y�û$6.�)�]T?����r�*m����I!	�c���q	`䡄�F����C�l�U�:���g@9��Vtt���v���H�2��,��d!�޹Qeh�Ʀ������;��w�x���v�9�R������ߍ��(��s����&� �L��3�,Ǚ"��CgH1��u�)cL&O`Z�9/��hC�Ε\6���P�k���]}7��s�`�@ ��K7~�����t@]�$�1>`dk��O����<�R��E�Hu�mu�m��t3D뢽 ے�42"��f�=J�N�=�q��%n\���=`/@�N%B8�K�����������������[2�9r�>a�V�٣G:��FX���9��|�:���A���zya���M�����zny5� &2��y���2�ҥf<�t�A��1�0O�� �n��e�����<sZ��]��L�V�clp��F��B���#w逳�����sT���+5�]�yϝ}��� ���F�=p~4�ޡ���-b�/����#]��	�H�2g|��1nd��o2���;@R,�n�� ��gc�ע:�y�X��������[�N:�W۵|6�K��ߨ��|�-���g�c&ȭ3�aPZ�{��\T�@|��kA�ڂ|&�f�s,���G�C'�N��}�:X0��9i4{�B_�.��aj&� ���ֹ�r��u�]���ֵ;���('$b��Jz���J]�t	m�UK�nO�=Oє+׮���
[�1����C���րEa�
����"�q�&H��"v�%n*njd�����6�`> ��S�f��k�C&7Q��5��a�vy�gb)�0��en	gx6n�V�1"������tmU�0��&�S�[��n�(����C���ܡ?�L�����
��͛�}'���{�3����=A4�,�J����8ǒv̞�v�z�=e��8g���,���k�P.����Y�ζ}G�g��(��詳��Zo��'F�
�.('��i�%H���߃66���742��S�B3�h{�)��XD���:�u�zY��N";�L`�'ވ{�
�s��]T�	@%p����tJ�lx|R�',�20Ʒ0�#V�hӥe5����	ئ�Z�����5�L�J�S�J4��xf,���9�J�(t0�ݓ/��X���ڽ[�t]����u�b5�N�z�ҳ���f4C�Fk���={�oQ*F� 2�s�E�w{��4�C��V/��F&y���ߝ�� �� ˛�!�٥G��L�#�}	�n�Ko0��7��!�i�yF��`w�{��|���L6
zcn����>mAy"f�Md�0�Ⱥ���Q���d
��w�u�\��� �,���tb��e��&�:�y��j���F�7[b\ ���B����l�C�y��)�r�����~��t��8����$&.���.������/��R�>�Lq�����p�K+�M�J���,��������B/"N3R� uyy�{cd�̪�{U�l�T{�+N��4sTI�����@Ϛ�\���}��L�qPb�>@,?���q��A�eemE�&F���曼%�V�?V�둬g���A��ۃH�~�F]��1�C��gW,x��b�F[qѡ+�#80Z�;%�w��{�W��������f�s��o���#�o��sA��aJM5{�~Qa�1�����0�+d-�v��_�d�K���8���o��Ol�w��n^�D��̄A��)�}��o����@���-��}�����!(�����jT��s�f]�6"jl88�MSjlF�IWj������yne��D"1ptpxW�
����'>!�G�~�oԞ#Ձ�s[Ď1�5��i����=r��E9q�����cg ĩ��عC>��ԈOW��e@R� �u�T�i��UPb����D608[�78n��$4� fM�W$�D�����-���tF��T�Fnue���Y����s�I�TK'� ��C��U��^k<�4�	��eh���p�a��d�d��,�(�:`��p��A68o0=���A���O�s҉s�D�9&aV��g�'΁����6���I��&�o�������=�+n��כ�Z�{�Y���o
 7������9���{�ʊf��_S֡���^��jI��18k�~�������bo���G'���Lph�Zu�!{�墁�8Ӯ���CK`�%8q�u8i0���u�]���k]WhW�� 9V��C���*��rP��=)����lf��}���� `j18��LB:M@(1�)o���9;7����X
�z �a�C���2�9C�c�όt7�P��DRI:@'-}�b��Z�=#<��4j��z�Q�?���\�x�/K��V����^��Dc��O����^��e���=}����o:���vwe���Z���|�H'�!�m$�Yc�"��z�a�����=��D�\�lo53s��^���b>W8W�K<��^�>�놺�@Z�~D#|5T����m���3`$��-�2�f5ȨF	��Ҧ&W.R��"��O�@���7ݠl�����dV�Ҟ#h :i�"M5���iO�n��۞ 2�h�V.�4r�JH��3��(S��u:r�o�����+?<&75Ӂ|#�	�K���,+[�얧���eL�5\hKI�h��^Y3%:����P�,����1�L�j\���'�$#Y��m%Z��D�< T;`@T)rD���Q8�L��zju���2`�]������)���u������'�tl�,��qx&4D����E� ��L<���Y�`s�d}��G�GLJV�ښ�~
��z�aV�����J�sh��կHd��>@��<�gԙ������rUj���7N�$�{��M����-�ᡢ��sϜ;'ud��\� �XG0���hC9	�`Ȧ����6��|��&~baa��javN^y�e��{�aٶe;Dd�p��Jx����?xA>��ϒ��l�i 3:6L�?��/[�/�����G7Q���m�w�3�ee�g�~�����}�㟸O��w�<��G�����{���2⌷�)�C����#�I��R�Fȃ�F{3���B������5F�����4��^�MV%^!o�A�A�?NZ����Z�_V���>ٳo�\���ՅEVOP�A`�	�W@�~a��.�"�s����k��P���s箵�����kwwZ���ApwE�4h��b�X�Ȫ��Aƴ���[������ޙ\)wLM��lv�f�X\�{�h��<�\E]3f��I'��:1c?ju��!�DI1'�����g&Cj� ��jf2T2҇����,n�iQk�#.���#��4"i�SUc��Yy�it��5a9V�d�^�nA�͕yW�;�=�~9�`�M;��ω�<F���lbF\�J���QU�
Y�lgU�{�W�����W�=�L.eߏB2���8`
�S(�}*��35=��]ZU�>��L:��t�= >���0p�!�IȟM�� K��G���\PC
����s���%#s�����3�WMC�ה��r�7Ͻ�q��A��o�ӣ�}6�ǌ�ԟD���{ �'�&��mC�)��C��X��h%q�կ^*��a���CƖ�6�r�%:'T2��Q����瞓��\�x>plk�:ecyh�@Oh��]T�戚X6���J(
�gp}�z�J��,+E���?"����D��F�^�d߮�6���cyaV��{����2i\C�Z�����xC����/�����?|T~��klp�"_��y�=t�fUG��{�	����� Z��9z�T4����2���ΐ�{�h�0π��������Ι�dyi���VT�̡�Pl�,�ہ�2`�d���-s�eM�2�1+MX������)���_s�_S �zѕ�|�� �w⃳�}x��c�������c���(f2���`�	��mR�̗�顿��Ϥ�8 ��K�Z;u��\&���ݜc�^4�M�_�2P/q]D���,�EY*$�����_�����G���rp�l�g_;!'�zKr��.��t�I`2o�c|
Yz^��֩i��C���S�Pzj(Q�Ix&�nuU��5#��F���Y%AcT��б�����8����Ͽ�����6���i��,?ic9�7�lb�2ipA��*G5�(s�䪻unyM�x무�!D�q��c�C��J�uuiM~�_����#c2�����~� ��\��^�# SpD6�]�נ-g����$����A�d>K���4Ç�K���e��+5B
l���ɱ	Y[���ù��5^��WN(�jU�h�	AyP�yy��r&�+���{�Q�����Uڠ��`�dn���6xp`poY w�3�P������a��H�<���C$9���:
��Y����%P�&Pl��&M5�� n~iY2劌n�"�~���$��񱒒ϑU�o��R��<�>��Bi�س�m��}+����ϓ������ګ�p4�c��l޺I��e��7�"o�;��AF�{�e�V��G>&Ց!�������޵�A,�'�9�����'� ��x���pߠY:��jk+,-��?��2\�˿�7_���Y"����*y�)�t����˽���ٳ��O��g����r�����o���IΖ_�r��� k|���<ih#f����Q�s\׀�pʤ������F�躂m(dK{k�B[�(b���r͠�R|^�@�5���V�j� �� t=���%�=�F��|��` UKhd�j�1z��I�R�1D ^������g��9ztY�X��N��rz
�+���I<�3���ind<�t�������K���H^3��I���&��F�mS|C	���{���(}ayYN�?'�φ�v4I���SB")4bh���B~��ʺ67=4Ta�P������u5C��l�����,^��Q1��46���!1�jӃ�B_�Uc7tt���4��Ll�]6�CA�:59%���rsNFA���'=N�q���g�e��u�-���EY���~[��j�Fo`���q���҉���b3ڕ�0��g���`b|�z^�,�)�cZ]n�X
��)A:Ru�� `-�$�VJ���僙�G�))x�^�˟�e�A���*u #�p�� �2��h�}��1= �����I�tc���!��nA�euFH�2Ku1���]�%(��}T��9R\G3h8�}AV��3:PT�v���^5�ѱ.R��sI+zm��y���"��.�v��߸q]~��O�^���̑�e��M,+�9s�#� HBMn��W��ӟ��P�ݑy8�_�����=<<��9����E���C����� o�e��׳}��ܸ�(?������2�ܷk����C��y��5f�����o}�k$�0~�~�J�]�������Uq����$���[�&�҈�w��H�m�:�z�p�3�]����y��~Bn޸F�"�OP;�� �_t+�s7���/�E0*�V�L���Y�Z��	��5>������u��Q� �=8~����g��KGS3�z��6F���ݮ�iK7gB���I��Ш�@�A���{�T6�}��4��9]䔎,�&4� ��6����_˱�	����PH�"F����V����f	����0�@��A�9��#JY���H!ň�1zv��@�kf��F��좼z�{���73��F�����cz��H�udt.����ܪ��`w$N|g���H���o�/�"�k�ZpT@�<��^kQӛ�;�0�}��;r����ܹ��i|l�4�˩��AB��H8M �80�M����^�G�&�DN����m���#�h���6؋�ڏ���r���0�M�"a��kF7�[@k���&@��:N�"A+�怅ӛ�Rh&�?_[]��,�_�w��6�?ձ���&��|�26�U��� � �WãU�'b�I�ʐ,.��Y�.��~Mf�_�@huVT���@��A�!����;�_����"I!]�7@�����3-Sɇ���|��!�������,��Ȥ�߮���H��V��	�9�i��y��Y��`@����Qi �.`���B������m�S�I��C'Lȩ)d���f���3��4�5�w0�Y@e@ZdӰ��R���wȪ���I��9&DPA�9� �>��n;��7X�P�Z`^V.��`���;�����\i��Uo�8��2AѬ�na~�z���'Ū�E�u�V�������a�������ߏ;7�'<��0 N��љ�qZǁCS(E����A���QC��Gf���`��<М������gx@�����9s��ٵ�1����4�a$&����=,x�y��{�5c���Q%S=���TϊY��,�!�Q���h�yt'F�Ԉ���I�83//�2�9������_�'�&Y���$ /�1��3��Z5N|G��r��L��s�v8�s����i�DӘѠ����5s< ��?������������}��׮��)�����A�P����j��|��Jd��wԃ�G���w���`	���9w_�'�v�����a�=3'�G>��B�7T:F���V�*=[�'�����;婧��d��ڪ,j���g�#��r�*z^ם�2i�Ȅ�''�����ݹc��7zr��)�?�C�WXQAK�֨�i!Csߎ�i�:9)��$��\-x�@���dA���R��-�"ǖd ��0���3�kE1�j�I�|��=��G�c}��a���L�!�5p��D��u��k�{߃�/��gm=�y�����(gN��z��F4軦�	�����u�u�=k�8��!+y��c�����B�1����_������1��s���z��x�P�k"((�7��m�ֳߕ�37�N���S}r����p��>F}��I>˷�|y�sNe�������ܬ4ke����@��˗� }2��2��!��	S{X�;ǻz�q�?��@_���؜hd�B�dy�$P+���)�(SS��03�ߥ����xK�m������%tD��*�O����4S8�f�5%9r�.��_�y٥�or��YK��lX@Ve�[�#�cQ>�pŘ4���͗���qn��hs��9�L,+�U�J�N8�'^d&�ר�R��*��	2��`R���8��!��*��@��3h�N��0��lrF��ﶚR���Y(���^�u4(��n�CG��c���1ҹs猻@�� '&i��O��سW��efn�._��|�;6h�_~$C�1H��/O:���� �9���Y��ٹn|@161*G��)����@��@iU�D�,n޺U��U�� 8�����\'X e2�;��0���5N0  @���#��'z��N����
�aj���8��
��$��0 �EF\�	�`�@8�s��q��y2�%�-*�(���g�;7���繴&����+#�¼��qA�>95%; �+�����ΫE#/^CO���"�	k��\�|V��� {A�/(�7����;2�0/+�`~(�KW.�}z��/.[{	�&�,�"�{̍��3YQ��X��Y�-�jK©%�s���C�����[����@	{
�����|�S�b������j����E�]��0彀��V�d��V�G ��8�y�������&�f\9lu�J�'�zD�uu��ۜ։9�L�k����N��n��?��q��-�5�#B��.r΂� Ҡd�*X�����Jք\f$�X�LJ]:1�v���~�t�s��&���"nx�j��I5C�)P�+��ۧN����Q�����,�,��vȗ�v��1yJ���^�8�>'����⢼r�5��A�
��D��1�2N�8-_�����1�A�Y�8^��mw:�@Y��5�j�m��:��yzJ����Y���ߡ����P�5F��=�V���#�{����$���䑇�j�~̎�S4z@�nҌ��_�:9s�O?�Af��r���[��,ö2��17���}�����,���Y�����cj��~�<;���>&G����+W9�g�ʐ����۳���׮]c�NY4�Sc�t�����{x�`/��!i�><s�'2�N�+�(_|��lQ`� ���i�Y�b�Dz:��PG�Rw��R�k8�EY'���wŪq4��N/�����o\9�`j�u����5S�ӿ�ŗ��_%�������V'�A��9mW1�H��CD��1�O�Ξ���/	x����e,�*m��4;�- �������u��|�Hw\*Hj�ZbP��k ��� �D����;%^{�\����7��k�˿�Y��Q�ܔ��n]���#o������r�����2�ǔC��An>��'�)��=�dm���3p_1�}���`�hp��u��IB٨!��i�%���;��$�juJr�xW�;�'<J���22�+m�A���l#J/�\�c�k�9e:�˯:C_j"�%k}dO��L��*�9�`�I�����L`$2t݈>���g	�Tq�,�9.G|�կ~Ք�rF�Yk�C�|���������P�#��@G�{vq�8�Ӯ�j�
jku"g�*ef2���@�l��5!jA��4��	���;x���&,	�Ǆ�DD@�	��zHFG�\}�q���l�
��v���k�q���ٌ:k5�7�\�#����߼��ڕ�e�D�s�=�q�M�D�"�x�}���n�;C��Fi��}�h8i`�{:t��{ָ�``p����s���&�dj��:`�mS˞������,Q��y�����Q�������lX�Y1���zK�����-�Kn������vA�k k�@?`74�o��E���l޾����W.^"���9w�#o�.1��ۃ��٘aЃ>(��������g�^�2i4q��#r��!���"��������*g������4���J��N�;p�Q��4��꒾�E*YaЎ9��w����/ʙS�eX������,����%޻�z,�~�C��#"����I�{Y��H�U+
���M�f<� C!�W�\��-`�� 4$�{���%nSRt̃I���q_��PY�s�f��9u��~��v�WOK�+Kޙ�Y/�k���ϟ�(�4�3C�*��٘g7�Jgr�.w�OxdK�$S(�kS#U��%���Q8uz�����l��&E7�J�e �@�O�gjb��b�ǲ�>#,�dT�#a_,eeV ѫ���������ₜ~�-�g��a�� * g!���jnw����6,�p�$�Q#S��4�	ho1�����h�d5]�W�وJ�y������xht�0!"����M�%u����E�k[�4��D2���*�,#�46(��Ɖ�R_�g/+�>|vUƞ\��⽶��%��}?$�ܐʚɶ�*h��w�f��>{���ݠA������}���~Сߎ.t�fd��Nz~���7ҝr��]19ZD�#��P��`eA{�<��;<2*3�sԺ�\�@�����K��}F�����=��^7�A�� �[A�p�p�4�ff���YL�z��)�s���@v��'�\�UP����'��?<�����������^�u�����6�������?��_'�@W1&���kP����IW2�d��fÉ�C44+ַ��܅�.��T�*	d����/Y~�Y>�ɏ�3��pľ��o���gx����z�|�WŲ�bYr�ܜ�б��*�-p�Bɥ���9�$qІ,{����c�6�y5��:+b�:|�L躽z�&�%�3in#��G���b~�Q�����5J퀁��_���^[��l��o�}b��OqLc���0f��0L-HS���*�� Ӓ;ǻz�q�?����^��5���z��۴�f��Ee:��/q��x=�W��ID�gT��N|?�>�M�HR�Ӯ��gO��o�y��X ���/�8@ ���G�(�M��$ɖKd]�{c�7b�@�]Qӿ�H��c�~��^G�;+�L��u�1߮�]d* �U&&�0l� ��qN#geu� �q֖�gm"�1�D��!}�qA�9ʞ�]P�����^�!�{vn�Y͖�|�S�g70.�0Mw���{�����3�ȑ����>���i����� j��)t�@b�Tv�<&�F��,����N��-��>�2��n���o>C��ߗF�����|E�Oo�׊����!��A�g��s��9+Cx>�~S�����{5�\�o=��,,/�u`�s܉㧤��������9p�X�3����O���������|2�U5��������p�QAB�sߑ+n�>|�F.u�>��ﰕu����T�V��~��5�v��tm]�x�����y_���y�;�bϾ�X�<~�=����_~� �s��<�I�\�?Z5���ޛ�}��R���#�Y(eI���˯����/��\<w���5 .5������EH�<>V"�HJ�<0���z ��^�q�^���U�u{����y��{� ���(��3�Q x^���A�`*�E����>�Ժ��?G��}<�R'���MyVـHU/�A��̪��>��[���e������C�	������R2G��dG�xAl�.��C�D�n��<�|�a���8�,n\�ɹ�nd�1q�}�挱{�8V���=|�@��_βǂ �эƠ"�IR��k|rDZ��V+T[ۿ{3#T0��e�4G@@�k�56:A��Z�A��@�P�ڳg��(�ӡ놾r�AX��E_��5�:�;	L�,:d����z�4\/`p=E �H�ˈf��>� �{�獲.z���L�3 �gp��U�r����55;��WY�?x�`_�j�������Gz����{��c�v{��>��ǭ}t�㞛��� bt���XJ���"���_�����S+k@U�댾�9`E�8<`��l3Ḧ́	��xр��wueMN��ڶu�����|������ҁuW�VA�c@�6U�PeIm0w�I�7�0� ���/}�OeP��iէ~?�Z>�����S2� ��AO����{}`]���8���r�E�'r���ݶE��d��Y�Ԭ�ę�"�D�Q5뢕�'ޔkg�hF�c��P�`~C[leaV����p�{�2���\8T�b`���=�Ԉ24�[Ce��O��O�>��Jڡ�'���+�:Z��}��S�o|���K��#��q21�� �h5�d��7H��뾚�R</�2J�:�������7D�r}ؓĩ�e#�&�:������vg2R�!5#����.wn�Ox�6�)T�����Nj�l,�2JT4.��f��A,ċ����~*J��#���[ѭn�͏qQ�ȕ�B���"�pw��>At0�������a�*V8���IV��`�����?�if� ���7d��ݲ}�N��~��#M����Y���U���C#�j�F���:�	u�Ȑ��$s��eद��{�n��adh�<���~����҆��5u��U�U�w�l�&Kg
���E�Qb�g�Ԭ��
8�c���7ԡg���)�s����,�`����P)
������s�p<v2�m��N�r;˛?n���v"_��}�>�o��J��E`�=q�X0u`�C��Sk�cm�lT��,�QH��R��	�Qk���]+���Ժ��o�;���G)$�
icc������������F|=�l� ��� t���{� f�ggo��W����3�<���#R-��UD�BO��BR ���,����ٲ�?|�u���ߕ���ř+�X���	��T��#������wI���:�/TY"��Z�Fʔ�q���ܑ�5�5p4��ί��3o�w���4۱��*Y��c ��D�QC���ڒ\9�� ���_�b�* fҊ^�9Hb��@���C8���뽟�}6^�*igmtIV�(ṢjB_a������`�$��|d�T���e#�ȁ&�(Hg��8@uI�k릩��/�8��'����9~��C�	����a��}_1a���:t�f��׭^(1�%�bΫ�AN��:��,]O���f�a��l/���|Έ�g��-�ǎb���B5�����> [6Miƕ���ܼ]&�7�Z��{���Y_�'yP����pӮ:E �ӘAH�	I`���fM
�ш쇆ʔ��`��COr#?������R���I9z��|���޻K�m�V��Ȏ�ۙA���PΟ{�}_��#�QB���L�5`�U56Фo���:]D�,B-����@?��엖�4p�3K�6$P�J�z��J�n�����oj���+r�$R��l�?�p�����`p0��� `�s��Z,��W�c�6_(�9�^��Ib<��flݖ�e@d���x����RRַA �De	�s���8!֐fo���|�ߔk�.9�HQ�|�Iy�G��_��x�c�d�K�E�s���\\WGO��t�Q�Y_]d0�B$u@G����_hp:!�r�Ae�����ZHXF���zM�JV�!>E��t��WF䇯S��&W/�����7���u9�g������UO�P�oB8��϶��D���h���_B�O�eD�JC��������r��E2���$y�F�65�����O�_vl�JfC��$?�i3��WN��?�җ�x�.�;�,���xem]���dSw��_[~T�/�oݺU���YM����{H"��{
c��R�5�2���$��	Y�C��k�#�B�l�C�̎驱Ɲ�ڗk��0�s�٠�#�.�QWm�	�\;�8��0�僜�3�ٓL���M�0
�����f3����H�mC�^6��q.ҟҢ�^�t���C�3�&��
H��;�8��iW��2=͙܄a�Cڹ\X1}9�x];�T�L7�F��&5�l6��kTg�lC���P�aiq����J\�C�	��b��r]�	�e���)�8#s�X	ؤ�
��9���:"]<�����a�%rk��:#/�[K���`�����D
t�Y��1q��1=���ݱKFFJ�yrL�6m���M�2�6�����,G�>�ѧl!''߸ WΞ�;h�cc�6q�����U#�]�q��#c�;tP���3��c/�$�c9�i��}˔f\C9�<>�ϯ��O����D���b!�Y�)�Ŭ�!t�3	S�됉�0���uZ�]�|�}\4��r�L=��$�(c�IuJ�3d����ac�0���7|=X6�#@��x��`?��3�ۏ>P)��]�'|���.8�2s�8FF3�X
A���IX��m���jG�������8E���)&�i�ֱ��������% �۶y�ͪ��oA�{@N�} 9�?4��@��P�L/!�1�PN`� Ԧ��ȃ����?��l���۲���:�ߡ��)�D����D����6�*�j"��e�^�B�k0z�PS�^�A�(�q[���o=�:¥�҅*B:|w40�2�JZI����0���ޣ�oR�9{�dS���%J�B�t�@���>��������1��
�h8�@��K3�Ə�`AF7C�\�f�%���������W`���� �+B��������+G�%���X^3==%[6Oʪf�+�Ȭ���-d��`JL��b3�l�T����dr������^BTteUu/b��D�������r�0�6!��E*�4��ǳb�΄ag��S�n7�S�\	�+��A��GL��6�)�?�~f�M��]�ˇ���?�y`f�Sf��XO������Gc	��Y�7[�iL�F�E3�C��_G/��L!���c���=?|A�����A\��a�~�{(;���#"�-[��!��F��(�1ջmY�HpY����:�$��ax��lb�9��ga?�&������%3�C��gܽ*q_�jW')�h(%���H�@9�)�p"f]��}j�N�<:�ѥPm]��UWG�鏮�Dm�l�����a���"�˲}|Dvo�&�Ɛfsv��l2����y�����pEraJ4r}uI
��c�Y���&2Ρ[�������1�}��]��a\3z�ih�$ht#v&PO_�*Cu9d��~i�2hT�]Ӓ&S�V���`�fĩ}m��>X:���>X�����pxP���3���y'�R���g�F�X
d6A���
O��A�����_6�q����Q�hW��P�6���t&���j-f}�4��`׎�S�8���"�O�<���0^�<������?�uC����i�e�U%��t�w�r+3k�%Qh@C	$�4AZe�,d������?�?v8��F��2 ԭ �T)��\YY�Y9o��x&ﵾ��w3�'8ێ�����2o�w�s�����k�	C�|��%��4>x��+��� ���� �K���^���Dl�JBP��j�z-�pZ���{��K�ȵ�����ӫo����v�#g_?+���~_z�A�͙���v��Q���F��A�5Y'G'VB�`5�z]���w�>�ģ��s<��F�ͤ�����i�s��p�RR(|�����)���5�?�<��|����6}K��K�벭�LCw=�I!�%����=S?[]m�)5�F�8ڮT��g�ȝ�`�?�U����/��Y�A �S��p�p(��0�:g�0u�JL�D7�!/]d�y�;���'��E����l�(;�38�mO�U�a|zz��-�Of@'�I&�vu�X���v}�U��N�I~2]�K�>%�S��qS����8x���l�3��O�*�C��&��Ȥ��$���.|Le�5��l���8KRNF=����!�&�2��-�_�2(��JnU<�խ�ac�f��t�ӟs�4����=s�z@�����t�(u���ܑ\F���rC��6	? ơgy}u�Ca>�>��ޔ��ei�!�� ��:�s\��l��>�!�{�0BZV�~C�N\J�XP'��LDŌvp(�\���}r& 2F�	"�2��~.E���꒩Se=D~p��qp��-.P����8����s�CWO��
��y�e�Ծ��xu�'l��F�zޯ�M{�p�!4��>�:^>�j��dJ�E�k���f����)��G[%z�����<x��P�Z9șmԻ1�7���!#X���}�硔�A�"rH��A"w@��9�gN�.k+jg������^���k����h^��%r�demC�ַYχ�QDMÇ�>��c�K�����V����>��<����2�H��L(3��`t�0��=
r�k�t�h�� �p����9
�r��%����C:��LA��b�
ty���p�΁Щ��He�*6�H��_�}�Q�9���8i6}����7Z��tXXX�������G�7���q����~T��o�i=O00i.
�3뽮��TA��kC�X�)�N߽�Hd�Ƶ�%�Uk�2�x߽��^IƎy����	�S��vÎJ��d�t�qi��Y���}�ւ��	+����S6Axk`S�Ic5�2���X������;��U�k�	�@��֭�@)�[��1�n�����`W��k�7q@8q��5�k��6��6܇3��1�H�dMb!j�`����ܥ-j��A����lu��_~�9w�7���KRo�$��Lc��JJ߻	#>��Vb3xr:�oY�=̼puzȤ"�T�-G���:'Ya�D��w �^A!G��C�D`���F*d��|���O��7Μc-��}��iT��z���gK�;my��S�o}�CaVo^�(D�톌4ڞW��'@[�}3�@.�KV��Z4���"ǹ���e7Zap�|�����a�� :0�C��{���g�~��ޓ�"��m�y8C 4@˿�3U�2�u��q�A��&l:�Z�jOVQy�y9�������Ɉz�yU=������J#�Q��羛�w�3�|Z|�4����ͻ6B��|���ӵ�Î~d� ���(T������K��):P��ۿ)���s.횹� �A����#��C��ʲ̶;|��5��SO=%/�����i��F��ޡ��/|��}��|�k_������V�)t(B�/����G��O����/~Q.�}�D��~�{���ID��(%���^(@����3�J�[�֮S��I����Htkk����-�q�v�6���l�Ȧ�V�9 �!E�^�:�GO�/J'�8�����j><4$�ӏ	v����%�k �?�����S��~��N�D�3�a03�lom0#��(�WҒ�x�ǝ��@��"��`W�e�J׽�3Y*����=<����] pt}<�6�+�&FND��.$��%��-�f|�M�I��d�$�rf_/�#":87x�K0�i�GeA�+/�MFe����8ܯ�dC�yy�����3Ap��W�:3��q�rI��.�|I��d��f���o=H7�!v����k`l�A�O77��}��2�&�b#HX�e��ԍz��t�+�hM�!U�zX:C-U��(H����/�:M�c�r��V1����H�95l��v�J5,}�ċ�8���ԈH` P��5j�b��x쳟��r���I�z��+���}G>��O��\���S�h�i$~��;�;�H5*�s`^�=*��K.\D��s̉G]��2DϺ;v����:#��� wT�L�-�TO13]#��yH�f��Cr��>���dI�̙��=[����R��K����A�1���d��,��	N��!���<R�uv2�N��n�{"Q�68����du�U5��8T�"�����>*��Co$�^t{*�vq�����\K_K#60�}�gIB'�
��}{�x�y=x�$jt s�uz��yY]^f�[�����?��T�^}�W3��G�����4�6��_W����s]|�G���ٶ���i@ق���`���wA���#���S�=._�����_Y�|�-?�ģ����O��cG��҆��_>�����^6f<K?p�˸F���\��*'O終��H�p�x-G.�t���rXY)PS�O܇��)ut P3�����hU�S�j��3p��`֣~����W҆yW�u�e�o��L���f�A�:���s,����<��;�s%��������m�R��AB��'�c����;�
�i��V����zZTԃa��{S�O��KI�7X� ?�����:P���^!kɌY��ΐ2���1+	�B9�u8*�x5T��fy[�?C��1u�����3M�7��Qǁ��(��Y8v��1��JRκ\[�s�(����
������Tyۍqӡqrn��A�s�v�
W�n�tJ]�e`�%/��$S���0�=յ���x�7����0E���9�;�Sb�#���A�zcֆ�@1���$5x���#j��F#�;��)D=�t���͒�4v˄)�r�ƭZ�W���>��±�A���~�����#��F��n�!?����:���TN��c[ŽH5NG;eT�M��X^|�E���@����Fj����ZX���T��>�Suh�f;r��Y\�,��C�����zx����0B:3�{���u�pD���P����|�?(������C�Q���K�'�y֌A��;�qFT��=z�:t��pH������{<��r��"���UN�:��|�m��UM��f����O*�����+g��d�}�������!
��-�dBO>"�aZ�Z�w��G�Ş��cG���0G�>tP֗�ʖ~o��g��u������0V6�}�gq���A4x��?w�'���|�+_a�L��.�����xu�Ѓ?�
��К��C�Oc�x_�OM�����<����?���Vf[����n�u_�sn�M�Y#5�h#E���Zd&�v�]�{O�á4D#��~;�Ya���l���V�x��<��F��^�\d��'�sXɩ�8�%chrl���>��N�>��ݒQ��>�z^�f T�/}��T���G��G�Q�Y�+��P>�_�7��/�{�ͫ����l,��� )��mo�3�{�s`�{8��}p!�UG�!�A�_O�"\�ti<� ������{�$�VQ1�����X_��7���F�a��(aia��^��q�ك� �u�ג��a^|9��5��j��k�d��=��Q��R�vPVa����5�M(�{��)��[��l�TQ|`=^��!5�ϸm�&ൡ0R��dY�ѳ�g�#�~+�p�2~R�Ha�V�Q���7�dR5p%��!��rw���
�A'���n֚���������7���)3�D�@��T�=���}�uE�&�|J��i�E�$<zJ@!���jN�8���&��"�W��j�q��^<X��;I9	�⨩�t�}�5��D8� �X�҄y1�O2�GL��1�C�C��^zLP�7��#*=t�lo�0���H�ߒ
Qn�jxn�f����$ǥ��c[2QҐ�a��!etC��@�bKҼ���C6ey#��Mk����nn�X7����M���9�� �����Z���g��٣���P3^$��s߷8�Q�
=�`��ĳ�'��]S#rk���^�ꐬ��Wϙ�R�47Yϼ=�^�O?�4ے@DC�T�V�7���Sr��Q�LU�j��Z�/�#��E�����W_�3o��1��N>R�A0&����sG����^h��ӧ_ui�8Q��gS��;JU$������AHÇ"֧c)�r"�p?��w�;�|T6������+/q���.4b9��<��wɵ�5��Q'�XN���p ��Ɂ�{�Ƹ�Fl�~�k�fܗA�:�(������{]����7�E��G�Y���d��\�|�j{r���SG��߿pZ��)���5)�$-Z��J$��=p�$��` �@�k+��N�U8��GY���GA�[5�����-N9ĸ4�뉵e�ALD��rggKΞ=+_�ҿg��#�~��0���ݒ�ޓ\?j���}�ϙ�}�Z��A@�fC�K����>���w����UD������hT��jy��{�����~�,�χ��a��쇭��kC^H���^)��ӷ�[y�Ջ<��(�]�Y����3���63<���e�͕w�����m�����V�ӓ*�h�+���-�o$��ߟ��e�^��ĉ�(	�-�#�;C��%�-0z0\0�a��1��i.�8E��0x8���FTq@r���7hY��~�1�;��+�H�_�铱y�=߇ �JƏ�Z�8Ti�#�����qG�|H���-�j/TC�i`?���P_C4��3^���s�!�����=�p�b�F�ߙ�u���e�;�B��~u|M��РW���i��^��5���Pf�[��oI\F�҈}V��k��9�>�~�Z�E��ܷo�3P�� �]iF��胬C��F�VúK"�q����&�C�����{�q���	���Jr�����mطwQ��ߐ5��!��/�8�ԔLi(�m�ݤ�G�66�w�e�F��5�>s�{ʉ�ψς60dk��@�� ����:3z���@�"���b|)��;}Yػo��k�c`�A�G�X�0�xMe��AaN�ዯ�,_��5��f���G�O<�qy�>��L�CZw��]2��J?~���۳����~`l	�̰+yĵ�Y���	��j�ȸoP���ؤ#	�����$�s��5��j�/�������$��3��{���Q��F�'x�����Jv���z#9�g����|����o_x~|�+�
Z�龱�I�k�Fl�þD�����k�<0б��7��n�	��oi�8��t2R�С>��$Ѫ�ױ���F=���+_0E��֔~����F��3a5�+3s��<q����J�pW`�N�c�8�J�g�P���#��ɯ�L&g�c\�.xD�$Ρe�pd��5N�,�/I���h �G&-���mn�[��M�L}-YT���a���i�F���P��ʅs�E4��z8r�Ӑ.u�����i5'T��ӓ�����+����S����A١PÏ��6z�us��FtE�G ��$MEl��롎����Z�>F��ܥ��
Y��'�MW.e���]gܕ7Ν�\D�Ha����B��3� ���"����KׯQ��$�&�͍-��]G���Ы��N�܂������8����[��yW'd^�׫�*b�~�r*�{��s���C��,����Nvص�@��L����Q�N{�d�c-����s�!'����z�� c�5��?Ĕ�	��=L�&����N�0� Y����lv�r��%I�ޯ��Иu�p2fi|@$������^�L��7�q��v��yy�嗤A��T�j<�cUc��=��N�Lk]]�gt����€_�(sqN(ҽ�N�i:=y��$��X[�Κ�Jl8�,�9u���GI���~�-Y?����?H�R�밥��Xc�`sk}|���6���4emQ��}���aG:1����!ǻ�Þ�!����$p�� ��2�.G�Z�8_�-��ܕ�Y�T�/z��,օ˸�n F��Ra�i��L�q��1�3��DWu*H?u���>�KD�|8��1�8��)t�֦kQnfq�$3�wf��`0h�P�
�vl�D/�(&�6M���>�Qo��޸�R`HA�zT���*�ᡅo��u��K�O�}��Y������E�D%�F��to0j6k���F^����2�l1L%s�Z�" :����6�9��G(�U�����]=��t��u������}ț3�l;B�^�a61�~�W��R�v�œF��4�to0t�%=x�hʇ�R8љ����)�o��y��㒡��шi��0[�h��P�F�ͦ���eva�m=0pb0D�baȌEED�"e��i���*r��oO��qw���-Fx��������~{�}2 ��x������k��w���e��F���l++K�`��������aFY����/q]����߽r��NݺC�裏��0�n� �ŇNvqq�Y\���}�+�寻~�;*2�9q�&PCk\�d��vd8p�8g��Þ�ٳg��p��w:�P"�@�@��ߐtK�0�@7VǱ�(}��аT:v�ˊ$��O���\��kZ#��U�n��c���C?2kz�о	u�7ϝ%����;c���{�=�{��VԵABľ��[�/��q^��#r���c���������k'hC���4�H��5R^�{{]�'HS�u9��<�?�kvFL����u��ž+Í`�=�]9 %�N�F�9>�H4��@q��,�`MI��?(kb��0�~��� ,@�@-P7J����E9����P&�(t���,ߐ�z�3��z�ظ��kU��5��-''����wqD��a0ĥ��N!���;e�%�{k�!>�Q�h�I)A$����u�b����X�ؤq����{���88^y��]Eo����o~�Q�oj$���_|��?s���tC�������y��ב�GY3쫱�p����g�i��ɼ�{B���=�ً2�J������K[��o}�;�G�ǌ^��IK#��o^��ո^�s�P����6{ҟ�������?�ȉ'd}uM���g���kd�c�4[3�c�q��/�Փb2�{2r�d��c�:�$a�v����=P������.�s�2�h�˫�n�5��!|Ҩ{��W_?�,	�dkvN|�����_�Y�p���-�5��(�D&��OPC�7��͋�<<�u�SÁ��b������%K�jP���QC�xԝ��s��d��wت�Q������H�=�{�[ߐ����z7K6
��wL_��*��A�����j�j�a�������K2#[䤒��B�?�u� t_�:u=�����l�h8@|G�ߑF��kk���*}��{�G��NV�nU��/�㑭j`v�g��F6�{��s����J�Y��0��욦��4�����������dt:�zF�0�N�m��h#�}��]:~T𮰊�����R�hܲ�Q�`�����2��&=�^���GԘe���gYDm��]�]��;D��=�2/r���Bi�pa�^0R�1�4������lkVz�AIԨB��(Z�n�\�kחeUE�A�đ�\�Dx�zA���0����`����{�uh���k����3����Q�� ��s\k�;d}uI�0�Ψ�#�������>��9�@�>�w�~W� ��x���"�m���������)[z�]�~����j��=,	6��t�slv7�s̛3��V��IQ��E�}��A��:%����W����1�"���tո@��̑����ḾrA��/g�3\V��;D|[�����C��t+�?)C;a�q�59������/�8���Ϊ��L�O�*��T���<x!l��I��sQ�2�=Ij}���H
���ա�^9"^���_�+W�;e8��"��5``��UN#?��W._�����F�!O��{Y�Y�{� �d�S��=�Iy����?��_�.��:s�>�i����y��S�T�DC:�1�G>���O���`���'�v����CH��C�0��:���՛j�չ�E(	�� @�[8��O�9f���w�s�K�$Ȇ�N��.�fe��5��Q9���L�FK#xL���U�����!�Rj��4*���~G���fZ܃��`�a�'bO��N"ǫ�Y@�F��:��}�S����H���:ǎ�Öέ�5
���b}#�`0ZђI�h�h[�7r4:BG��8g��8�A�@��̱��Z���N �sA��d�w��E�]�$�]��;D��"j��� -k��Hg�>�5b5� �%��9�k~��1y��#�ة#��W���`:�����{��&�^����hĎZ#Z=�ȩ0A�+��2�υҞ<~�91���'G����T�B(�ax��$-������#�~�U���z ���ғ�A��fcc�ξ��ߒ%|��B�;�X�#W�F�="&���pS��;%��[�k}�i��v��K_�Ӷ4+z�l����믱�٪˦��gސ���K{f��KKK�A����	<|�"���o�ީץ'��qS�mO���g/I����=�:뛮7�:=�wz����	�#��m^Ǎ�E�$r�� ȉg�;�6B��}_�ԅN�u�Jʴ2�<|�z�<��<َV��Cq�f���P����U5y��$K��� {0�&�q���R#�HEJ���Ww�z�4��g��zW���x���=���6���Ȳ�pF�H����l9`��BlF�[cC2����Ad�k���E�uk��ѽ �G� J�R=�1q���?%��`��	����$��Q~A�����NG�����.HT�O*�V;8P&t��~'�3 q4�wd�qA� ���#2���u��ޛ+���Gn��˪��	V9��::+p���FD^D9?3̈���߭��
)D�s�����Q'#?�Td�"�*�) ����!u�ɗ�n�իW��}�{EǑ]�<��P��.��\�:��>�2�x/�>��sY��I3��nG�mJ�������ZR�<��3�w�b�T�b;wĔ6�k�J)5�^�9$��<r`Q�5+�7���� ���׬I��1�;ۑ�3��{j�-��t4�F+WH���+�yQ�I�����Fڨ�Av���~�=s�	!W�᠇��ֶ|��`mmH���mﮭ�VH���x�}��pz����w�یv�T`j��?&�4�1afNC�"�s�='/����������)y_ʍR6ַH�9��=�j�&E{Q��p�~��'�Sv���w�S��թF+��z�`[�2����8U�j^#�g�� 8/q�C��P?#,�tA2u�7��Q���aM�C����U�)�Q9���P������vv�����h��O��H��wȦ�'�MͶ�ة�Aw �1�^(O�Q*)�� 6���RgP0lM���A�n:�����p�￠�����&�dEv�e6���2"4�}���O^{󒮧�mVp2]�g�H�z}gt��t��uC��5ɫČ�j�#]3�Ĕ�m����|�;1��.[��F���ְ�����Kv}�a�s��Ύ�q#=��I��#��5Or��5}��e�`d,J#�ֈ�-7���t8ޯ���˫���w��Gz-�92M�:��'	��	K/z���Ϝ�Ca
�ͨ;гh��ٺ�}ymU^x�=_f�aPs��wr���x����� v�QG�z��Qϡ�R�����p�V�*2����ڳ�
��8s���{wG�<΂�Tɒ��N&
�%�k�n*�pW`��A�L=��s������}A<���:)O�<&jೕ�ԍx)fT�I�	�0E�N]8vP�m֋���k�������0�7X�Yz��0�a�cV#*(iޕa�iZ���u�-b�
R�dAO;f)��Mo�=p�Ao�d]L5�7�V��иohT�6Dh���G6��@����yh"rb�0�z�crՑ����pߞ�L��tf)��	lr8T���{F�z���V��ǟ�Y�lj��H�M
V-�gB����`��K�+D2F�j�ȉb�\ ���:$#����H!��:b�-�a�~�mw��8��x�U�Z�;�up��ǽ�zt9Xd4�E�zo׫~�Vt��6�꿷��;)����EDYw*X�����a�ú:��� L�]�bX���![�ϭ��l�:�j�4P>��+R�h����̴� ?�?ec��AD�%�ub>mh�זdk��#˃:o���>�\d�/����l�r\��s&��!^W�U�﻽��n
���U#��;sFZ�n�=�߽�Q�~�2�3��Y����`AͮQ��HO��U�V"���<d��@nC��'tڑ�@���9��"��y���*tB�ƕ�
�<�=�s<P&��Z�h�nӏ�s ����:�_��7/\���_��wa^R��phqw�r�u	�'�gE��=�_\`K.�3�W�Nq���?���[�؇�=��+z]z��D9b�K�FMc�8�À3��>wvI����
N2qLO�=�`��}��ay��c2h��QGM��l�a����a8t�QO��{��%������E}�kNPEC[W�e98��L ғdO�,���P�E�|��9�_���Y�8��g�k�[�GT�9�	/��3,b��a�PWg����K���~G�߸�zgw�/��u��Y
F�8u����~D���1�`�Wu�s$��ϐ�D[�vh�!+���Z�c�X�ыN�JvA��eh(��MG�����y�!S�y6d$8?ߡ���>��d�i��t���"%6�Qa�6ĊY�;n���E��J����\'��I�]��O2�+�ާ�v?��S�7ts�>8
�Q��U���w!
:�x,c�]߷��]o��T0�[D�y�K�c�5*��H>��C\'����F�� �w]���}������j'O���WoJA"]{ssNZ�pm�N4������]�*�k�c2V(]]�tU-����U�bV� �ԡ�P�~s ��}A��A�N�~p@�KH�B[�>7��Q�h`̏ѐ��A�� �]ѽ�	j(̈́3T�Þ�z�z����y�49�h)Cڝ2��"�j��k��օ����"(���'�:+�f\��*z���w^|�Yt�D�+ѱ� �V��/�Ѷ��o��2�U���^L�"(+�r?�]>�H��V����>/�i�Ӓer����%����^d^���e�A�Cd��ǉ������%h��C���=�'��-�ΙWe��&��e���Yzӳ�b��}�0#���uY�ؔH7����>.g�_��`�3U��:s.	��Hq7z���%�_G?/�0)�����g;q��s�0�+Z��=t�='@+�Z"��%��\oo�Hz�q�!��ڊ�jy�k_�uZ�9�z	9`�^�tQ~򧟑������/�6W���-+PYC�T7���0gІ�%�w�5�A-�N���z_#���S}D��Z���7І��V"��-�"���o�#C/ЪTs�R��H�툽�ҹj�:�:���?��A��H,@:���ގ�]E/0dN.s�0|;L��� �Uq�"U5���wfR'yGc�9�C����[�Z 
�z�u�#r"p]�5��\T����=m7k\#�J��������[Ő��udj��g�,����^�ɹ���-�7\ȉ��H���\��Nb�b@<�r\�� �j��4�k�=�E:���\�|I>���F�����Ѝ�����3�P9E�6At�CYv�
�^t�P���r����L�?��F��^�h���N����#r��uY[Ybv��a,}$�)��k,��su0�&��u{9���t�v��������A06���\'�Z\n��S(p%38:��a�Ɩ8��� �1���1qkl���0Q� �RҞ+A@(L�4ģbw͎:������b$�PT�N���׮�Ɂ4r�8�����$D��n��"�c
3�e�N���n�����G��JjT�$__V�&/<�H#� ��{�*��D���>�<��G��/�_[�a �ZN�)\��z�,z��5��7�7ds�s�Z��d�z��us6����9�E�n|�G �n�����٬;��8�p ো�n�u�XD���=�a�}��-[0P��(���E��H�}�V��59j��4
���jW��djl�q��mA$��W/˪�.Qp�a��wZ��[[��smGJ�/vx�"��zІ������]�ѱ�	x��󲡑Z
�r�5y�<�n�i��3������>���W�G�/���V�;�+5��>_D��o�3���Mt�z���k]�O>�8�X�C�B�:,`>�[�硍V1(��SN�� ��?H��)�/�*�{s~�F�=5�[�����T؆�1!DC,��w�A�q�����q�[Ҥ9���;Ͽ&AIؘ&�C�u�b�ۇ?�A��?�3y��e�S�{��Hs�#�8���mb�V�de}M�<��n����r]����3��4,:0�9��j�c�u������1��N���1����oʂ:����Hרm�}Е3J�őe�С�E�nܯ���L��wT6���UR�3��#�r�_�Ǟb�=Dw��a�"U��s��9y�F�|^��u��qq��k
�(M�c%��B?���a˜����!���a�h��4��+a�T�W�"��3�w����iR�B�ؚ8�q�&ڏ�����7�1ZM��}�A�y�� I�!@9��9Ҟ�deYV���a^�< g�a�c�M�9�~�36t��WyՏŭ}�3����Ƌ�j�А�{�R�N7��@�#'�
�Ԧ��ƈ�?`-���56,����_��~��g��ߞ~M�!����I��ξ��5��Fl���.��]f�;�Qw��Hw#�ό��<_���;���=�)Q��r��]K�^[m9s�M���!��k�CJN�:P�N�w>��~�}r`aQ���O�=����R6����!������)%�֟�SGj���e��!�F숇h����5\����%-����>�JF��������%���V���魃\*��� K�^�A�@�ҟ��^�Q&��x����?$���'�Ƈn�y���Ɏt=����0�����J�92 �{e�&���*]���-f	��dpp����j����+�Pc�AE��b8�&�a<j�icC����勗��O >wp�>����Y����K���<x�qy����ڥ7(����������F�%�!�ip4@��N�����6+;=��@"�"�Y�+U��I�.��t�&�w�P��qm�tͺ}
��T�������3F� ���-�kJ�e�9�ا�YS��"F{��9c9޷�E�����ɘ�:d��_*���s
Í��yud�r�)Ҁ�]��Y��ުI�y09ʳ�����~~C��!�B�G:͂��"g�]�2"˗F���0�~�`2*��.����V5��ںyPGG�r�Y��=bF��^it:�a�
��YW�,�p`�|���H!�p��;Sk���`�8���ƌ�t!���Fn�@�mJ�挼q��l���8K�/�t`I����)dq��x+��ǌHB�9����"3 Ͽ�:u<ݐ�(I�ÿ�ԿA� ���i������WjDA<c*��]FĐ�:,Z�P�w��� ��	?z�/�k�b���M���)��{"���k:�᠏���"x�;d{F
5r�s����W?/�j\9"����\�S�-�?�{�o^�*{��k��_h��%}�U��epKD��H� �6�Uy���2��8����C�t�o�-�d�O������]J/���V"�����נ��L���;%�����ӈ�3����O��������C'�ˉ#�d����_����n�HA�����)(}�G�������d�J"��ۖ�K���N�=��9��_d�%l��^���ih5`�����s�����	��?��<r�	����C��񁯍o�Y����-�(��h�z�+�����Ak=�a<�ǡ�Т���?x��os�!�q�T\t]�9;EQj�� כ�T=��+�]r>��;��̂ĺ'6u��MZ����~u�߸�½ 2j�$<�O�k��.�� r��Fz¡
_7Gʜ��DO��w���H" Jd;��mr!J��]&���3�Y:���#sa�[W��B����T��:����]5���#Q��)e���s?0�,�87�|����]��;Dؠ\�36����8�6"#:�@;���7טΛQ���i[��꡺t�<��,�~�FksԥU��)d�AO9�<Wc�f�h]#J�D$�#�4ݔz\'ZK%����Jz��m�j/
���t$֯���'1�a/����!)�̑������>Hf���CϮFTHy��H��*�FD$������/�ka� )<���jC=Q�~�j7:d�����Ѐ�VD-�hꭺ���!t hg�b��^���ɟ���ސ����c����Uչ�E����!��y�	��'������,SҨ��>�콼S�&�������M��?}ӵ�X�K��Aq�U�iu��?���w�sD��>J��N�";�1�SdA��ݔ��O�<�a)�������yM^�{O��g�y����'z-A�D_伣Ǐ�aΑ���t�7e��Ȧ~���˜~7�Q�G�����ҫ���*�W�7b�{1� s4��˫����-y��I�T�������ɾ�^Fyj����d��l�������hp� Π��h� qL_Y�P�?��]}߭������[Aӏ~�=z�4�ݻG�f����)Јy�����'g�?��G�[������ݑE]�I�-˗�K<ۖd͇t,�}����s~���o.�z��E�~�:u.�XS���\�C;X�7��H�C���A�Lf��A��z5]�]e�,���^Uз��%��9'�˳Ξ�wE
��h������S�ck�&��y8﷜�O��	��#Ix~���Ĳ����#�n�:��$@��%-D�h�dV1�yI���Xb� �/c]��ٻ2a̰3�w���e�*��y(;�o��(�C63j̇��\t�b�zזo��B[�!	l�x�5
�f��Lp���$;#N4���t�3F|~�J���#�"�yD��\k78�aM�,F���P��V�nT�9t�Y�Y8J7*�Ќ>'Z�
��S��g�x�ԟ�	�*}��$oUƫ.1z���Y5.=&<��3,�a��}� Y�%�-t1"�p<��V��	*v(� ���ܑ�;�p0���#�Z��pLm�	fa�0���;���T>����3)2Dò+��{�Nd���X��u_5HY#]{��)9��s���%�IF����c]���QC���~�M��r���шx��5�:���xN6ז$��9��P*�nI9B�vS��^~G��F�1��}MN�����M5�_���~>�Z��J���8�(�N9t��8������- ��V���r>Q��[�\�������\�|�S����g��'�̿����^a{!#Zj�ǼL�S�;/�BÄ!(H���
3�r��8r.g�iQ�ߩ'e����k������x.��R��F~J������="�h��� �.�lГ�M�J�Gl���z��x�{��O���:�.���J�^8�hh���D|��a,b5��;���������Dk���r7C N��Y�q����,&j"Ǘ�p�i�$n�a=��.��,w=�� �+B�_��&	9+�kH�Ȝ6{]�̓���&��Ʈ5#�"�i�җ�ސ2�qsV�6z����ڲJ?m���^���xӺ�t^�(t� �����1`��懭R�{�P�C�����K:� hEA��t�ņ����.��H�ii��#�xcVI>�ΝDd�Y\�6{Yϴ7~�[��|84�<Eξx�6�H��j�o�d�"�s�_�=�F;��~+$v�42<zbkܪ�7k��!sPi�$���h�Bt�N'������}$���(uS�HZrƁ_���e�t@���u�
�t����X��/�1(�����P��ď�t���b�N�,�/��n��f��6���ՠ�demE6:�����D�>�`��o�m3]��`}e��aH)�<r�r��%�gѾ	#؀�HP��B�a�ݝ>u2
2�"����$Y�������B���B��dWD$g.^���7���y����ǩ�w�����РC���$/�������r��Sp�0n��{�������Ò�o_���둼y�<�5Ў���a�1�~u��{XnO���R�j�������S�o�3'{�vh%K|� s���р�Kٰ~.�?W�b\��@���o�2ލ�Yk����U�h�ϼ
�Dۜx�]�c���:1��w���Q��
�����{#
':6�_"�USw��p��P�A�� $OA]XDW8Ȯ������1�-��i�|�)czp��3�Ӓ���\"�)�7�ܐ��c�^���>/�仼�5X�09�%r56����������/8b�	̈́��*~C���YHu�Y�D8D74���ٯ��4�DJWdS���Oq���o��k����S�Н������A���7��*h NԼ+��ȷ	!r�v�����|�9yף�K�ݗ��:������`��+���8`a� i���#�����5�o`�H>�}r�*�ل���JŚ<���G��.D�a1��~��:)}���������^M�z�*'�!�;��ޘa����ʊ���iٿ� ��q�@���"�i[EK��]5�+r��5f�
O�;~�<z�$y,�}�yy��F�x}�������܌�<q�|��ǶXc�q��'!:R[���_ҩj�!�K�BVyZ�[�F��#���I����B�����l?k�+o�!����&K���{���ި=����_�:-����a��f�� ��P[F�����/I����Bvz)ʽ�
�&J�^�����'�S9v� 籧z͒��;�\��Xa�����X�x#xW�v�����V/�c������߈�J|�v@ ��9��ve�%q=�Ϡ���rc�sߒZ��A�5z��>��4�X�&tg�w�YO��sDn�����I�}_z�U���)Y=�A��0�~�����I)���yY@mb��/^�'�I#n�pԕP7��'��^����"��hpym]g(�l�޼,Ͻ|Z��4�D��
=v���&f^<C;�	5� r�rH��ob"@��؊ҷ�UQt�;���Y��&txd�N/�2�i����셯S��ܡ2��ǌ�}L�xWT��O�����L�m��a>����p�'�v�~�WC���O�������K��a/yK���NWR���s����Y�}R�����H����='���3�Ѓ����&��/���;�Ņ�[È�kutF	�B��=ʈQ%FoctFM���(��D�aQ��}��ι{/��~�j������W(j6l{�y�ъ�摭yb��'o���9�^�Fj>/�N����?۹����;e�)X��7���|�"6i������I�����֠{{�q&o�2�Z�9`�.�f��
�B�+�U��F{:�Ű�L�-2H~Eu���O*�TM�ͤ�u�q$�C�ۢ�̠u&˟�͠(�������'�[4Ny���mX��o6P<Z�$)xݰ8[Ҧ��%i_�5�
=��f��>��J�p���쉚{Π�N�nkK���j7��_�u��s����X�)1=��aC(^"�8�$��ot�u^��5�`�=64}��2P�R4�����~�հ؞0�O���2I�P���Hz�T��H�$S�lwB�!��6�_�0!��������]�۬��{��L9�̭��?^�{�nN�����v2-���C�E'������_K����6	�'ᝁ�������W���T�U)o�-g�ɀ�R͡:�B���{v^�Q,�KY��w���,�W�P�w��<ϒ�+GaW�uh�e�3�[Jzf�q���rM%�	Z�{�N?#��!Q�G�egE����v���̪�E�娢] ��/7]=�'�W�k6���z"z5���H��������q���X�l�� _���}�;*b+&�Nj.�pb�w:����������r���p񴧩��LA'���*�h��j�0���p�"�����}pP4�M �z*�y��%������m���S��,')\�9��@�e�l�=;���#:�k������w�^�-��;���[����R�o���G	���p�?�=�,{��T�А��왵H��Y���cWFRul��j�y��%%^�SEyL6AW	�o������m-rx�E���%�X@���y����o\D��L�-ZFҤ}�Y��y�?����d��;��(�P�u���l�����LV^���	BM.�C���6��o
*��1/b�D��Jߋǂ[���e�AU����M&"�O�_�qeE��_��X�]=Ȼx)ͽ
3#���[��"Dݤ<̎���΃��'X��ؑ�2h����n���x�u��0����h��s�(i��]��<�@Blh�,��N��p�� o�q\M�6م�l=��kai�PbY�?��"e`AR�.x�hW��L�;�+��NrN�� ����ʲ�	Z���rb������@�L�#��i����5~��$tP{��r��h|e�&�ōW*������v\��z!�Y�ͧ?ݯ�=~������?��S�m-�zGDnM��`C�x��X�񁯏�u��,��u��-�T���<z���L����2{y^ `?hB��Ey�sm��+KJN�=����*�LUH�a�PmX<1=��.~�($�^���I�Co>>��TX<����y�I0t� b
] &�O��o2��iZ�Q�����3;����˰�(���C<�1�i��w�
%�}耺���X#l���Qo#�O@7U�4��u���R+E�	,��rSFQl:���Wz;�j���j��N���7ݹCu��3'��'Uk�a�X]�$e�I+4�H����f����`)I�-��n�}ZEB�N���oG��=o�����nk��KBR�pY'��#���Cgo�j*�?�)3�x�.ʙ#�r�Xf����(z�P1��cw�����R0V��E]��~Hٯ��g\T+.�s��� d�⻜�)v���r��9���ώH)���I�k?؊���g�.�3�9�\��>�g��۝����V�y�>����}p�]˹��,�nC��Cg��`�\Ӆ�Ĩvؚav!�ɯOJ2�/7^���׹w~/�Z�� �Z-�Pڗ)OE7��z䶜Q�� �2���O���z�Y�K�~��G�&[��b$���_���:2�����G�N\�P�f�y�&]41��Gԫ�M�WZ�R���\����Gѱ�a��2����gp��/��$�Juҗ4BU)tz���e}rg�F镱�>�~��V_ܪ� ��؆MP��;E���V|�0�׍WQ����`9\k�Sجe�.�9�~~V8��,WM��d�o����t���l�dI�_'D��xҸ	�64V��d$��>�7�U��l�+�O��>��<9y�*��E8zq��b�+qR��I�x$3l��r��jF���qJjX���c�$�r}Ԛx��b���3c�u`M�	��� X$`�+�����6����{��`�b��	[](X�܈�n2��<�ý�@ �MF�B�����IB��Sݬ
E,b��g}���� �9>�g6��L�ڡW��ϙ2�`#�.o_n��:xQ֭*��(e$Ga蘫�oG�ڤ��$�`-�	�>k��+����*?ߖ�������f��T�d
�y/�.˼�����4j�A����;
���y�dϵw0Z8��y��������#w��AOݿ�h�e�$�@���؀��������?�5=�+٧TA>,��%����oW���i�O=�o����2(���e����]EF12=��7�����X9u �f!sA����r2G��J���r���*����:��A��w}L�ez�2�(if��,9ƭn��� �&,9?�b]�� h�UIOH�8$5�Xz;�d�wC��8
R��t��Y���d�CL��&E#��f*�%ɳ�U����VndЦ�i��8/T�̷8������]ƒK,#z��F����$�������.?�2�f5!̲�7P{�|�*O@NQ�(�.��O]�W�o_�ȇŁ<�d}R�'��Jx�r���w9�\7o��i������y�.�}��լ�
g��9�(�3j�+����Kgpn�������{�`���B��+��e%^��M�J�47O����iR�^r���z����$fH��<������8�S�#�g��=�/�5�d)[1|��,I�*k��<Ѐ�g_g�)��2��8*� 	��p��J���</��>q�-�5_�%��~�e�U8����t��Ҏ-OY��f�9�u��� �S��3�c��?� �	� 	>+(�.�U�����uÿIV�6uQ�ͱ�j;F���iTTg�F���O0�X�9�)�N	��2�K����d�,� R�|�5��/C�n�,�΍� k(�,+�S&2R�D�.��+��aُ�6tۚt�'HB�D�S/�e���p�����t3������g�o^��J����r	'�J�䱎w Y�������L���@V�@͵x��%�j9TAGH�i�a���}HD/�(��)��Y�����/��H~%,jQ,�w*1��8p�=��%v�<���XZ�60�S9lt�C�
�Mxw���f*�s�eK1o�L�3�r{e�`��h�1��|�Oɠ�р��2�#��yZ-P ��QDI~�W�'�UY����~��PM�\�OH������� TYAߪI(	�c���6
՝c4kW�����'�L9�b���k����Ko�xȚ}o�p����Q�|�Ñ!�{�{D� ��k���f�A�Ǝ��Be���%~w<��6�)|զ�Z1�n'���GҴ�_���+x��)�ј�Xg��0�)��b �FzP'G�:s��x�%����l5�͘!�/a.@�O��<�!2E4A�r��H'p��vw��p@�3�#c²d8�C�b_�];�s�f��(��CAA�?�o%|e�dq��:�x <���s۹���K�	��a�RzY����j���.$+T�V4�h��{�3x�XDXi��A��>i��p���{h_� �'j-1 �e�{b#�O�������A$���\W�S��ؕ$c���b%U���{(0u�c���W�^d�A>�VK"L�Z$��u���o���=2�vk��JM��M�A,A��� S<�T�-���:vfya���n�i�j3R��Q\O�7{G g~ӊ5�ߎ��汶���B�]h&nC�j(씼H "j��'6�*�/}ؒ�y�����9`�|��Kyn���*�h��Wӷu�,ej:��U�w7��	2�,�Dg��-x,0w?d,)Z��(۠Cj�J��b"��fԵ�n�+�vWah��YN�����(F)+���5�����������f7k��Țz(g��<B��l�q<Q�d̶d\-���T֦,/�|�QT�z��n���iU���Fcz��œ �WX[!���2C_�Fp^�~���ڣ���b��TD��i �
��׀-�*����s��^ow��P�=+RBԖ�� ���Ȫ�kB4,���/`I��|Q�d�����%ex�_��B��G����T3��q]�����<-H*��ٳ`�т�<}?�"�+]G};���US�S��Gx�T�X
0�7�f��4<��W^`��qL7M���T��-VO�l嘫��g�6fغ�5$B�4���Qa�o\p�4��r#j��ぅ���95�0�=j��ϱ>$��m�r,6�@u4����J��$ }��m��9���\�Gq����\�,���bޙ&�~1�-->��
׺;�s�����b���S%�6s��l�O�!$����m��]3̭�<��ԥ����3G�#��AP��3���U&��,Qm���X������T��iM�~�^c���?��B ��U=������wA�E^�{�:n�d���uP�{֢�0dg,w"�~�O�[�ww�|P���������Ո�P	C"A�(j������=.-�,�К�3~,�$w�(�W�@��2~��5&�s�͒�ò�M¨
��g��������A_��Ϋz
K����"�p�󭖏S͖�13��V/ɠ�7y
7cŀC���56��=����#�Y��U/%��M��#��}p!�m��[;�k�L�9�@7�8g�Q(q0؞�m��<V��7n7�RZ8��vp�'����f9�х�nfh�>+�V[ܧ|�į���0��O�$Q�:�9������g��Ѝt3��3�ۢ&"�?�VO�&���+7�V)��S�"��X?S�v���M�E�Z�e	�=��M`^��|}�u��p{-/
Ϊ���cJzu^%/���{���<.����s��ͫ&�㣔39���B�����(�6�z�g'K����I�L���$&����]�=ͪΐC^x��U�XA�o�s'O������5k
�@���}���۠���ҧd� �N?��@�8}`������Zx��8ZR�tBO�� ��$����G��v)V@�1P0���i^ؠ+�����ږO�xw��6��͛B7*:���7!�<�����
�n�D�+n��:�Z���7t(����wsZߏ�YD�(j{��n��o�Ne�.�I��L��b����Bw�H@��YX���b�Ԓ�](��7�����6XHP��/&* ATh{�^n`g�BFKn!a��N"�S��x�_?���_�]�he�XԯX�t,�F�W����� �,[���0���]OI�O�p�h�S��|Yi��+
���;c�;��Js����M�v����J�_���oPO�i��2(]��h����͸�]��o�/D��6� �Gc�Ld�ݢD#���	{��Z�+����؈>��/�/�/�/�/��
���+����$v���� *Y<2b�
<��{]a��l�v�DY}��o�p<��Jn�=��i��U�ؼ�PK   ���X���-PC I /   images/af9fcf8f-e29a-4021-9780-388d342ee2b4.png�{�{^��ur�vr�il۶m۶�ضm6�ۍ�46�����ϋs�s�7��f�5{f"�%`q`A@@�$E�A@@@@  А������}�8Jj��� �{@SiqA@���D�T=s.z����R��/�_�:�zP�bI��A�?���������X��)��ݱ�rQ��������� )"�o�>V=�V����þ��\^��t�_|\z\��=i-�G�&IG��H���9���9�1
�u�F��������{�6{ay��R��t������EB�?�v�S��F�Ŭrg�q��{g�����a����k����ϕ���g��Z�Z�ْ�ܕĦ�A���Y�����m�Ň�7�h^�Ex�]������盧x ��|a8A'�_��)(�g��~y������yl'�ɄM�p���6�+"
���п*ʓ!M䐽g�����}�uh�z;=;20��VX�p�|91�z�3�ZR����Ŧ�#�����,=�y���i��8��8ĩ&�LY�J�`��1���h4П�����^{���t}����w.ԩ�=�u}��.�I.v���}�����H���O�N�s_��o�&D�6�@�tp�:� 9s����P��MD�������w�U1:V�C��&ڗ|,���}���.�D��e��������E�e5��܆M��:t��>�}}��=�\a/�+`����I�۲�|iT�yM_Y���D%`W��
T_�0]� �ެ�ĦC����R�w�+hl�����m��>�!9����$�e�0�/x���w�<'�ʷ�_���\J�,ml�1Yz�/��$dd���"!�?	��!����gѤLR�Y(�A����Κ��������	vm��߼��\�߶���d�E�sm<0���V�}.�ۭ��W�r�`���kI`�����U�@Ԥ��e���>9�D?5��2��� L�����Ͽ ����0G��fl��Cm�>�����l]�1�>��'�N$Y�?7/����}�3-n�5��ͧ���-��L +�t0�I�dz���#��}�l�iL��m`eP��{i����]�3��@=A�W9�xy?���dlיcp9�k�}���|��?[���͞Ӕ�����$i��c�;�3�L&��nj=�������~�L��S@�~����1���M��9��Y�gB���z������F��am��<�'c������߯��� an�O�P���sB���y���>W�B}:ᢨR����!D�N����µw������������Y�;�0����׺��k��-Ɖ<�A��-�t��К��2�ӤܝZ�/�6�l�^��e��ӞG�[n6e��]��~4è�vN��K�e��C�]����M�~�8��O���q�	-���a�)�\o�)t�n�?��"�{aBx �c�<�b���Ӡt�f?����>��&3Uڍj.ֿi̸�?��X�����_�S���|O���i�] �_6o83�o�iL`�mU7������g��	:�Z ��� �Y�1V�$}Ȯ���b�a����[��������~x�eg�r`���B��v�1��8	����h���Q��W����L��2�������`w{
I���C8
�<�<�r\�|e���}���>T���?P��v4�Q��1P{�&��5�|>_��=A�c|0�.������)~~�ߟ��7c��Þ�^^j��	b�J�/��Ir/K��/j��w���\i��
���2�Ŗ�T�(v������U�!	!
�a�N4C/eL���<:�!���7��y����劊�D�4����r���.'���
)�Ε�`�xc�B������鐎��`k�bڿ���`��1�BN�0hL��?���d��r���K�r%N��*�Ð����z�_� /�����O���^�~F��`�EKR�f� �k^��f���=�{,�oG�|�i����$���ߤa��5�@�e���G�"��*��$�O�%�9-��N��� |�	t��W��19���=[�������G���S���|��������_x�os��3Q�C�S�?�?�}�P` �]f�$0#�d��R_�N��֛�*&S��##��Vh������C
*sB��V�gЁI�.x������K{#w�\�4�]��ܕ�����wH%}��QL5���T���h�r�Vj�����=k�����G�A�J(p7��΄��Y�:i�o�A�}�v�N }n����������?D� ��!���#_l���W�b�{�&����Ls�}<�2��>m��g��e�Փ
�.���\a,'O����O��������*F�̆�dA�C�Ct��˱�18s=�s��ý���3N�t��H���B���3̆M�D�3�`�!��ԑ$2���b�tum���[��}Nu�� �K��8�¬��$�h�sj�լ�~B[#~ެ��μ߷֖��K:���y�}5miw�o����Y���J��c�ˊ��j7�y�ޮ�E����dw�͕í�f>�χ��e_���V��|�V�S�t������g'"��x6�K�O�t�C���s�?l5�3UR���*%Dp4&��*�N�-���N�����s�E�����1>b���V�m��C t}���f�����߷i��Y^L�˅��{�ik���
��.�����|+�*�ZF��ؒ�AlH���kf�{�|�m�A
�}fo���={c¼n5�z����A�p��i�Av�Be߰!p��l�̦�|�"s���$���M�M*D�����\�!�s��Lr?�/����$/��C>dw��¢N|�HK)��c��P+T]֧s�;d���<����ӹ*�'���ĭ�/���zߍÚ���Mx�.j��,89��'�h�m>*^���Y4�z��i�����+�k���_V�
�J�#-�uT��J2L����=v�k6�[n���%���Kx@�>X�/��%�X/WA�P�u���|}z��j�̛�S�Nc�[ƚk�(�^7��������\P,Ĩ�v�UO��a�h��J�4]簿ջc�������J�j���*b}_�-}z�~��w���SWd��Ҹ�"��'�֤l4%�n?���Cس��Lc0�Th�$�����֩�kԫI�N��-���:��q߹BD,,�U�w�����oO|U~���G>z��d�7/䱇��o�>a����sbg���F���nc[��1�%�/~�|x��8ݲs9����l�
t�~���9c�B�'�f�B0�@�M��W����^��N�+�V8�a��5\_���w��&'�k*6�_SICU��1j�$��:�2!η(�<aS1j�n>��DZfe�˲S?qQ�&L̎J���9�:
]Nye�Z��Z:�O��[6���즋���~��CV�p�[��j19�.5��^9X��u���ǉ�6�b=s�U�_���Xj�0�O�'���C/ d,�"�k6^#�p������2W�$��2\�vX/�r;Wk��ɧ�-�n�>i=����R)J��>=_�Q����7�P<+�1q�J�-�s���D�Cv-ӎUb���W�B���L�6�l=����=�"�TZ��Z� ��F@]|�	uk'����hZ�
�k�R��j��w>�:t�S�R�=���SϺ�x�(vx�2ş���8$� ���V�� ^�,q!�Vu���~��Jm���:�/���ئ��������jD�0Ҥ���+�e�X��EĄI�3i�hx�y&�S�r��~�o���{�N6))��V`���6����D��|���o�Z$��XR�g��)>��8�*�/���/ua������z���@�fq�4�������������WL��)���ۭZ�L�O/��XL��Ɇ%�5��&k���U'�պ�}f��&�}}�]o۟�z�a��;�qd��EfHqA8��;��l':�\�v���P1�]�Y��OaH=U��{&�ԭ�_T$�E����˰n��h�m�W��M�R��g��l��g��i��&v� ��)�g�7�MF0 a��Ţ���@Z�f�����߻#<�@���Dؽ�`�j�U�\��R���f8�*v��%$����F��+�~ns�L|���������"�%�0�hJP�� ���]�r�:��ߔ%��V.e�������tg��ʓ�["6��2���Yy7Nf�N��?v9
PЂ,��p�� C���d՝3W<�6��Hm?y̾����NU<j|�+D)�c}}����,�"*�F�!ro�D��1���Ź|����",@	I���<�n�H5��:�VF+]�y$��]1 ���`��~���Kg������uO��,�M#�P�2~hi�3��99B�|�[�g�l;��P��5v����u�����7M@ԼHxA-K� ����>�L��{}�H]�d#�3,���;#+CԹ�%��Bֆ�F�K�g�����l���,��WPB�֌>�TO��wh�1�6l�]�.J�[ث9�N���.�9ʐ|e�DF!��i�8{�x�00��:�v�����̉@l�x��O��� 	1!�B�~��^[8C?J���(!F&R���f�~Y�ج!vӇ�"By|D������/X�`=p#������ur��Q�n��Wè��QÁ���c�h�- ~/r�'���?^r�ku�ݿ��5�0Y�9�M/�����8��|��e4��A���!Y.t!��b��fވg^�,n����q����J��Cٕ�{(�m")@�ɼ�|G�c2��>��!�&�OVvoN�J��1���+�`�P='m�<�
g�<_s�J�4`�e7L&��}@�b���r_�jNB�/�5v�����b�dd�2񭌅��c1��^��D����X�i|��8�`��C�����0�%2��<Խ&&��ݾ�avpc;	�q����Ċڻ�8�Y���ɖK6G��1lrA�xpIs�??88�R|�7�	hDw3�G[�5�{\
5Hg�G5
��������S��ə��QG��`?��|	4ޏ�<W�F���垾*�o��eW�5��S���<Fz��<�H�eX:eo&9�t��x-�3�����0l�>�ɨt����H�_�[�_z��o���|�9v0��$�K��?کa�ԯ�E�|^��?6B</�<���(p9.��6m�6���+�@��4����R��p!2���s;up=�tM�ȁ���v�a���}�b)u����C��Xh��<`|a���)�T�a ��b��b�۷�{<�����A5�/D�ab9�׏rCHs֜�YYnTC�&â�9r��"Jv���lɢ�aH�<��ϯ�G��޾���h����6o(fG�˿U�Y9%�����u)��j�k��|b�ޔ>��X*n�7A�k3�	�y[q怯=8x %�p���n&M��K��ѻ:AE~�<��e^�jί�����6� ����M��A��+��a�!Fk�[OC$����_AD5�\�1�F�+ �����m;]�~��U�Y�=�y"�����V�k���Re��P�jIK} c�1�+�O���L��K(��R?,+��+Y	��$-|����l�!��e���}��0�?�&K��0jNT����d�� �[ѰP@>wg��#�m�b�$�c2|���^���K��r%$_.��b��Qo�Q��mN�.ɷi�j�\ELX�מy~t��}Xm���v�=e����L� ��<Ot\}M�Y"��k,6�R�o��ǡXN�����H���Xt��\�]����͕k�R5qty��|l�AR�(̷��7��9��Eu�E�H�j�W�� ��:���M��pB��t�!?�/|:�������s�B��X�Z7�����}�op�c�T�=��Jt+�x�g��U~�$�1�Ti����o�/��yVJ%�4��f|��g9�`���C&׷��L���v�l�o�r��C�TGv��Y`��iR����i0��!}㊠(J&N�`L)Z��^������[�_\���5�	)4x��XM�&b'�����LM�.#%#�	~����OS�r���*���SZ��,�7М���R�����a�|L��ؑ��;���ө]�>1�����H����uZ�P��Af4	����r���g�x�Zjr-"��4���k�Nb0h=M~�qQ�	��ZF�q��'�����a�Ga�ôzޮ݇N_���^����Q�ǜLQ]�aMGN�!6����������{�q9�y�W�NV�a�H� ?K�
@:`��A���'x�,�2/��]P)6������ߝ�D����n#�)Dr���0�ΨC��lnH�Qq_�A�p��$C�����4\��۔����O�j3 ���D����2����*Mb���j�	ws��1{�9��^ ��ڕ�*,���9z"9�F������~K�'���ڥ��{� ���jr�����s����'�H�`F⃏Z�۶� ��ߵ������?�%��j��2@���I�������@���V��MVU�BFqD
wcX�OA��~!�a�*�~?���i����\�`Y�J�";G�/@��Z}����[�P��mub>cj�iD�-�+5����tb.(���TQ�V�
��:��l<��V���.G�͟���Qb7ā���E~7��i>�6Le������9*0�,(<.���Ov��?�����ڲ��U������!�)V��)�jK<H3פF���p���� 2H�m
	>H��8�6oPmnշ����%/�����M�x\����Q�����(}�����+�'��@�&��?wLUZ�V��JI4^S��� qF/Z[V�HA4:��IUi�h�.d����l[S�$z�N[63/��Yg���c+ڣV3�����y�a�"񠵪�X���0�$���M}�h�7b6<@3_�z�T:{������@Y$�[�`-�������[�X���ݓ���-0����sKl���Q�wk,���M��V�)�?��;�(N�=$�X)��,�MS"?�eDa�0�A�"O3Pb"83*�����N���y��"X�G���
1vH��P/֤rVf����z��`I`!� �v���ldd{ݗ�qʩ}�6�J�N�����S���VS��N8�>��+~3J�5��{�8`-��4迾Y�r鑜_�n�t��_:�V��DNf�ʎ�R��M�g*q��[X�z��l�d�M�Ik�B};�_�fq&�p�|4�mۭ�#�~xF���aI0"	â_����|a3����J�;U2�_�1���&���aC_�a^���8᪛!�͢o�Ma\;6��T(�2���-6�ϵ�b��a�lbj�!��h��H���ղt���D�%MM��:ub��^}V=�r.O{r-v�3|.ǋ)�NQ߸p`^�����gV�'��F4*��g,XO$nv9y�r��'��3�MڢMY퉟�6��!�av��e$�@m�q�T�<������T߮\�o\��G�H�ѫ���iX�Ҁ��}[(w-<e�=F����z�˄IL�%�[�5u�3E��SBSA��9!F Z�����%�B�T���v;P�D�1rY��&�ł^/s�m�Wx��S��l�WBv��{ԃ�^
L�BF��oz.`ʌ��B7�ay��T�UO'���e¾����Z���4����2�#?G��հ*�ao�,�<�t��T�J-�x�ܮsB0�g*��:-�Oe�z�CO�7X��*.��ʉ�4	���P���7p������z��T�k�]w��Vi�T�&��V�]oy��dT������ZU�H*�nX)7�DD��Z��:Nh�c;���?�H9z(��&J��DR�J�49U֭"��Z&���J���K����Pp��l�`p��s��r�@��a�[m�P%���F1KL��xK���*�$�O�/�5�GUW}p��Z�cm�_�v"��P�'ŧf$/��NP*�4��~{%�:�w�{^���vm$�P���6�w��S�n��ٱT���Kw�e����,Qy{�Xl��/H��Q�L�(��s��r��oZ@[X߭��_�>�kad��J�
�'�a�7��
��!�0�����|�(��0����5�d���}%��Z"1,��K0�3/b]�DX��ɂOXT^(��6���oƙ#$+}el�Tk|n-Q�'F��Ȅ�%�cZ7�,Wg�,\���5Wy�m�Xs��(�0Z�sl���'�b��8�_C#=h��7���y2ST#"]&�����L��}ݶh.S���J^�d���	�h)��23p�$��i뵂<���64;������A&aC�p��з
�������U��N/�bY�E:8HVHT����O�In����h��R��dh��J"�f�T�s��8�k��Pg�t¦�>�� R&{���l�0��j��S!B�Ҍ.�M��eE$2`����Л�Qb�9%r&�F�'O	1��Z2����g{{�{�q�/���F��ÖN�s�4 �?�7ݓ��rn�n�9�ݎӺ�<�L�?�j�(ߔ���H/jEw���%�s���_�`��b�4*��SH4J1��G�z�K��Uv�N�U(�0fJM�70�I� ?�!�����ݜq�ɪ.�vj�I;X�LTde���a�=	��,�?OFb��i����tGj�B٬-��7~��4��S�����`[ �yFK`�("���=UQ������tP'A2�24�*��p�D*Q��5ũ�	yN��Ă�%�at>���!�����w,�o8̨��=Ƙ�Ē��I��P��	�q����M�~��-�Zx^i�]�kI�F�,\)L�#�=T#��(����b��Lc��Y��k^� �鋈��.1�f���+8�<��*+[���/�`�+-"$�p4����R��;ҝ� l����|�:шу#�P�J�x�h�̎�W;��7%�@b`�9�~v��X���3��w�X���t	8���`1���,���0q��U�,�o�+�����~M�,�����&8���K`��P�kG{�m�CZ�ܗ�?����W�о^HemIJ�w�V+�D�����qť��$O�*���߉]�G���������<*ƥ�u�g�׶JY��,�)	� ʤ��f��=�,��À`�ݠ1ußj�TO��l�^*c�[(��B�f"XyD���h�n�f� T���-�n9��<�Wu�0�5�a7n.3��M��\1���Q;�)z,��	��|�@gxC�D�^�Z5���+/Ns�� �	7c���ϱn�WM�q�t�_��n��2��Ϝ��'L�UM�U5ř߾t�����ċ-�o�|�"�C�X��z���B���6��$����Ꞻ�K��)��eF�j�T�XXf%���Z�5u��>5�HR�f��Z0���Ƒ�
Y'ZY.�Ɵ�0F�7�xN^4q��˾���S3�Y��TBm&�k��'�R�㠓)�`��4���瓦����2��+2��m1���ަ��c��h)�7Z+VM��aW��xK7k����)_e���|0��g��m#��F��c]����̸b�А���s^�X��~����	gb�j͵g��뜡K'ϓw�7/B#�~�����!&�$6B�]yD�w`Q:W&��E�%����]#oF\A/]���RbS;>M��W�����hA����B�I���1�Ej"�Nf�Fޑ>��cSo��{9L�;i5�@�ɲ:�Tm�
eO�����Np�̖Y�G�OB1U*��[�V/jF7ح�!mz��ɈN�o������2=���U�&�|*��p=WR�룡Cg�q�>������uA�SY���6K)O�8�L�P��hГ��BUP�I��s"l15o�Q��f�9�׼����8�I��~UD�$���
�e$5**��Ö��$�I6q?��a��f)�bk������۳�V�}q�}p��S��nLL�;SY�2������)#3�՘��D ����L�j�VjG���勽�ŁJ��@�\(h<�\Mwl���"�'�/%[d��P��k(�`��@����><o	�M�J5R�(X�����hL�Hu��x1��07й���"���������W1���!ZL}���7=B<��wQ�t��E�F�<���U��Xxg��1�k0���j&�d1��$�o�$e�<IeZ�N�l�巐&_n%�mܵ��i�>謉��_�>�؛�bѭ��Ō�q F�a7�3�)�pMeF����o��t��r�Ӡ��ݽ���A2���0v�]�G?e;�NSѩ��D�"��\�2>	�X>7o�#{�0�U~>V*~���i$��, X�u�)��%��T�"�K��,�S+c�e~z�_Q���{�(꼦wZƱ�;�DK:�?��\G�4j%e�I��a��z+N{��p�أ������:��PMM���`t2#��N�)�ƭ���]X7X�0�{�c��L����zO���/v�`��K� �?�,��!�^$��_�},�B^qA�$�d�w2u,�51Ϸ�V��P:��XR�R�"�͘Q�EH�P �"!j��T�����>UB�!_�xc��?7�ԩ+;=��p�f9I-�m�t�+����廃kiz1 >,��"��[�Ͻˑ�R�����/�����"���q��Z��9�z|��/���x�?��'�}�d�=�AC��D�k�B?� 41JX�Ԝ��鰰�����R���y�׬9��J��2e0����V��GX���Ë�y�Fe�҈g�9�7v��j@�U�E���mۛ�B9�D�E*V�:frE���2-Y#6�ϧW5'&e���*���/������g���@I�ȵ�9,�F�j��E���AD�>�[��B�lϨ*�/�Ɓ�rm�um��;�[j>ڇ��Y�Pם'���0hrg���Qh��v]�:�����k�X����L��B�v�`�JWp�^
�qD�Z:�z_�8���ۓ��E-��[��V+l����KQJ?�#��L�>"H���F�����l�I7�?��_�#Xid����1I�H�YIo�7�\�J�0��iK�-��n�z�6��8D5!F�qD�h#�X�{6Ϫ4�2��~�ep����)i�!)�6���@s�:4���9����,���g��[� �д�q������o�"E�?f	"��R��R)����n���0D���烒JmUB��b:�<1(��0	��m��|X+fj�E��㻡��?T��$�3��{^�{1`p~~�x�U�Df�g�m��Q��DiKT��[o�CL󪶈��bT6`�S-� $�Y���5�{�U���٬�*�O9��ai�Hz#ǎK�T.���_ԗ"�\P�/����n|����X'X���#��Y�������fH�9e�b����]wC&:e)��,�i����1���G� �=����0Ψ��T�����2�K0��d��,r�Fp��6JѰZ+)�:=fש���n�ЯR�&�OΆ.��@����t������_A���q�D���9=�-�����	��F��cɍQ�Y~gR��,n6�&X��-L��2�5�]��!�4aic3�H�R-}�T�ٗ|��׌��a� |tN�=p!B'����)uk��W�hp��� �]Yms����t�߫�Aj*�X�g��W ���2[���ÉC�}4^��9�̐
�2]��v�<��+uk�!�4j{�92�1��e�d^ǎ��+=h����hR���Ӆo�����v�Aȍ�ag�9e��eq��E@dէ�7E�c̺:e���+QP�h��`S��_C�ĳ�� [O���
D�B%-���Jz�Cz�Fx�Ġla �L��Q4*1�}w�{|�6*�+suײ=L�����&�6�����-U�I�5k�"��'`y�2)x˿X�.��\�uAcmLҖ?Y�D.[�N����r�����-�1�p:�����f<8��>%`hw����n�x΀��x��,�-�@��z�B�Y{�'�>�A!4�b�"�M[�-+$!�3r���ُ��V�����mY.�-v��\�O���2?�Met�}���<�f�Z͌5~p��
����%�U\�):�ϊ� ���t���|Mլ�EV�8���z�� �מ�C�X����JKB �|n��2�uy8a���\�|%�w@�������nm��ܴ$K���Ot��'*~�3�1RE��+���۫���ᢹq0{��>�Á8�ąǩQ�[|����y���^�J��Ix"��ߤ��M��_�Nf���O��\�W�C��ل=��.�p�.��ɤ�^
|1Z�ғz4���4�&Kk1����
k�$�0w��e���5�IG�4��[[P_g?^bW�F��XT��8�/v�S_VJ;|�/��-m�����1m/�
��13�vGŞv����	q��7�֙��=�(�5��uo.)�dSS��,m���،�kӍ���i�>b/~Ӣ�,_Ϩȇ�0�1�Mfx\��\���pK�?��J���z��c�̟��p쭌%��Nփ[v�<�`Ӑ����2"5��]�f����i7���f��n��D\�"��ΆO�R	U�f�E�.q`��'}(Z�l�@�/��� 
q�Ά�.v��e)�M������lz�O%�N���
�>�F�U!�]u1pޜ��VUD\��yn_�ϧ�7F�A(����]���}�����y���@�?h�n0&��n��1�q{���Րn��t��u���+�C'�EEq��QG���=A:�n�L��I�<;Qa��/ń��� B?Q��"| pFR��8�d�sDQ��&g��6)���lh֍O��sV����
��z8�=�J�	��HF���鿼��F��;��_��.�`������9��� ��ɴ��@��s��?ʄV��Mx5o������O̱�L��%��+��=�����\�����J6�t��������q�.�d��2w�����X\�>s��|PEV�%	���H��ߘ�����Bx|]Sh:/�3�����������h"�ɍ�s��lV��=惆��K��==r�,�*�5�Rے)��%��������m_<pqa�_9��l�F�ݠ��������{�ǰ|��� 7�]2��ٿ�����6A����2_CGL<�0��{>��U����R�Jagn����?�O� �__U�����l={�R��1ZQ��@�Kũ��W�ՐD��,J6�D/Y���qG1�k��33I�� J#|�BjA�4���*�\����_P�A�H�@;c�8Y8n���/ �B�l ���wc"��y�l�o�c\��v���.����w����P���#Hwh�ø������Nyu�y������U�L|?*��ڨxIt<Ő�l�@_�����S�x�/( �q��-R�ؓ����*����l������R�0DS�F8���N>�|5Z��\',���INp�����V��R�x�8��h�k�IX�����o�t���zWEHdI�^��!i�s�\�V��T�X����+��(��eÝf���B� $ɁV�)�V'ɟ�}3/���A�J�t}�]�;�j`�m�q�%=���!IŢ$ٷ if�ڜH�nᅗ�-Kfc4k����BD�<փN+��֮I.^�7����uh���w�p��[��c�:	0"���y �|R�g����^>���wZ���w{�:ƨ��)-q�|/p/ŴQ2%B�G�ɪa���q6qĬ�R���P0�0I\�1�|�i`�����R�Ҍ��^r��3<~g������#\�f!nׇ��������Ȟ��*{�ap�댎�7��
��Ğ<�۳ܤ7��z��ϔ(�M2�4�mO��4�{���L�7nN��W��1_�@�e�z��;����ˇ��;��˴��!X��g���F��%T��za2NG��@RR��s3*�m	&y��l<.��M���Vl�P)�:Ο���R�ݱRDs*�/*�4�g��o,*Q���o��L�?I�b���t�lث�%���E�=e�X��|��,���L���qI&;��=Ar�m���r,s�QT��i:D����,׾,�V%y:�C� L�|*i����)yYU���a��#S=e���L�+�dy&�T?5s\�)A��Y�T)�d#�i�7�&�'� �!mm�?�c��^��ؐ���~WUH}DY*8FqO�e�T�l�wFsYe����±a�>�{ ��C��Z�IH톺X"2�
��$|��h����	X�z��d��8�g�}@H�*4���;A�z�&��.��;4C[{��Y�i�:�x�J�U����ݨ	`�%�(��O�,|T�B0�����C4	���4�7�V��8�ۊqC��Z� �D���)��UH�K����t��q�Չ��$�s���N��(�0CWyK���S���;ma�*�_�up^?�,`0c�R
���`��0�7�Ų�m����I�Ȟ..?>�$^qw���0� q����*��8�ʅm&�Ou��?i?e��&�0qp��@�s��^Af��IM��z�F1k��5oV������=��ݔ�>�q�S���O�Z��Q���39N���dU�Z%Aғ���<hc��ٷ����lOK��ZL'�I�l��;B˾n��wq���
�7�D�7Z:Kj���פ<c�"�|�<�Unj�f��1ßc4S�k,��o�d%=e�x�E�?,W��G����)± �A��b�Tҿ4��O#���#L�D~�
�ܚn�Y:LK;&��E#p�I�{�����7��L�Ӈ�3��;����bk�z-� � �ځ����v�n�*i��̣���6
���,�(t�N9i;1��7�k69t��Yz�����a�د����CJ[���;~�ֿԘ�1C��;�d�c���V��Em�,�v�-M!utq,��aOV�g݇���5�n֏�zcg��Y���v�b��'o�Y6���'��Ǘ�E��i�^჎�+�Ƭ��5� ���b$��&u��GT[E�̐��%-�x�M8�儐�~o��_w����������Ysl/b=P�W���k�jB���쏃28���Of���E'�D���Њ���+�*��ykc#���ˣ���!n=x|np2n$v��%62=�AAL|ٴQ\e��+&x��R�6)r!~�$�OI+�I@�eHG��T�7�r���}�8$�B>��K'JI�2�;��t��~�Ţz<˨h��:�d�t]	�_=�8�*qu��+���#1:Ri�^+�p6U,I[&@�M��TT�]+�?4pV\��H�� �ݺћ!P(��ģ#��I�6KȢm�
n�SV���'y�׏B�R2Y�םŚ_���u�͞��],#�@~�8X&�V|�D����	"�Ƚ>��HD�D5�=��Bp)�m�x�eyIU�p8z�!��|���G�P5�s;�����n�X�FAEz<���M��tqP�`5V:"3�{�S:�4_��$ݒ��&�a��m�]�a�\����i�f\V��J���h���΀sM8?�/[���4?C��*�mr`��U��$�I�P��"��*�?�WO�K����dU�ծC�:�t�~@���.��{�ۖ���&:Ҷ*���߸\�~4tF��Ly؍0ԕ@�I�.����9�� ���9�%r�뀁QEHGG������On8h�b+�����Xx���<�u)9ͥDW�r�!&�����-�خu�J�&�`��JS5@)�o+�"y�����A�A�нd1�b��=p����6ڹwd������>�����E��wwWWV�C*2�mW��`b�MJ'J�63�
l�b�.�B�a=�v#�؁���m��j���~�,�,�F��Mo�@ᜰ7�$LE#zS��2:K��n�����k	��@���lk�-�����_#D�C��b�h_�`�9Ѭ�O� n$�ݠ"�hY��95�kUo���(��MoQ;cӨx��pU1��GS������?"�KTL�y����y*��?�m*�����_JҖh-��|"#�'B�d��a�ʍn��[$LّϷ6Ш��b�cs�3��e�ӵ�~�kM�ۓ�i��@�"�XZ����E^��/���g���޾�4�<�B�6mN��Os,���G����d�@'ep��9_H�F���M���'B�NxE��2��r��Q�w|%�<�2M-F��ʩ�9��~�Oڿ�Ԓ� ck@�/=T����b�d6^�J��xLb��m@����l.�r�~Z�>4�i�3X_
_�yT�b�q����Z�2w�(�dhRFGK+�G��9�!�Vr&��nʅW6��=N��U+�`"���e�F���x�-���-+G/�s�9_��9X}��1m�<^�'�R����#KJ�(f*��&�TGZ��{�Hu�c�1�r]LOz��(C�����K����51��'�K��;�E��M�wm�9���M3"6a��k����_�c������OL� ��=�B��y"Q�u�Lʕ#NSl��9l��W���#<�J/0��}:)yfa|6R��r�"��$�����gL�V��~��:�~S�O)��J���ǞFqM?�w�!���i�� $ua�%H7	C���aRsU
��~Fq =�^(�EM��H��$�r��r��"8�l�؋�C:0����3>�iL�Ms^�б�i9n����Q?�|��8n�}%xBg3pZ,ĮT�Q]年[�

�d�+Ș�@�\��h�ʌ\����uN%�Uv����ݺ9���ndf��g|�f�lDk��N��>�DIdߕ�5��O0jzV�c����V�.�q�-�'N<O����)�<�man\���E���0����>d&�l��3�l|#D�vUby��E,"���Z������?r�N�,��(���>-��FZxHg~~��q΅��#�·3�B?+U;+���]B_�-�����z6I3�^c�ta�*��T.#��ٜ�\C�Ym�r�s�����\�qcGI0
���pt�y7������:���{���"�)����k?�C����J��ۡ#7�}k߫̿��kn��)���	�Nˠ�{����ww!�߅/|�#�폷�)���X16�W亪컛6m���ӱj�
�S���۱_k+Ҵh���h)����#��.��%��R��KcC�̣R���ͅ�Y�)AV��$��0�����i<���7n�/,\���t#f͚��:�Dys�^M��b]R�SU�]Tcژi�gL���x<�ހ+�)\�ӟ�;E+EGЁz�Yt~��6KZ�2i q� �'H��Ŝf�	�@��/��a�q��N����F��7��A�Z�mAO�,f�1���򯜇C�:?���翅G���P&Q�VzĪҜ?��(��]�6�q�2-��J\>�<��Y,��}Z�K��%L?Ո��6f�������|������w?�^|�����>B:�4S�k�F��[���g�z���(�!�1u����\�����uba�\y�}���V���cp�_<�dT^ڀ�O;3��������*<u���Dk-��[_�
.��7qW����ǜ�'p�Mr9��k�6�dN��5�6?���Ċ�Z(����~V��a�(�R��"�T��?�?����Y���b���$�țG�z�P6}n@�@U�#��8Rq��8`�0����q��ඕ�q�`ݚ.Rd�j�4��%�o9 t��,��܆'�H�I�b4�3�=�8���M���~�z�<T�E�HL��H�D?c)��< �;�h\���ⲳ?��Wm�M��c���Q�O]�RC�؅��]��z�|JL�#Z[���ނcF��{��w����tƂG��fE߫k
	d\t�|�_N�����O|�n�q�b��촘
��iJ�uĩ[D̢�6�^`��/�J#�HB�Q'��֎��>'�oŚ��q��`����{�)1�rD�k�*r�{?�6�}ŏ�I����}�{��u������'�0UZ��)[������[�9J5jt�P��;�A0PeIQ����E_©�>� |��7ix��7�.-�I$��&{�<ŤB7��<� a�H#THq���)�����:}��8�������$H�����#x�ߏ�g"o����f���������E1�Q�݌|6+~9�R���Z���JU��9�@|�]���}�w>���w�/�>�m���%������|a�Kj����o���"�P-W$7���k�z����q;�ٳf��/�+������˾��t�V������}�g�X�=�0�������U���/~���p��^&��z%�N���mS�l-d�s�<���7�;?����V̾����.P�Y�Q�V!^U=���Q�O�A1��M���D�e���/��k�;��E_Ŝy��Oɾ].�rp	L$�7���~���& �C�(= C	a�O
�V�Wk8>���p���������:���}�ۤ�G�y2��ڡV\z+_������ڢ��r�$�>B�\B__.\(!�S�NŴ��I0�r��/.쬊e��N���j--��*fO��e�=���Lb�ϛ��B���["�Y0j$:���k=K��WÆ���E��8���b�D��]Qg�`��i."��:,� 1����7����M��'q� ø)��p 	3)K�h�ȶBW��f\�tk��޼Q���"�}e5�x�)��*&�?s���Ȭ���]|�l2�<L��`��[b�}%aܝ#F���G����1�r��?>g�F��*�R��ظ�p�}�쩢VyQ�
�w�8�����]�&N?���A��I@13�LV�7��%��Id�dgS���ڗ��F��ډ��VH."�)9m=b4��JJ��5k^���#5H���A�w
��w#�L��Z�� m9���C�I�.�K�������Q� B�lK;���O�tH�s~��C��R�*
�S)���+��}��%��w%�n ��о,̙:�|F����:�3w:�H%���B)-E����J��F�U����s����Am�؋�S��K�~ �� �����o�k�I�.����:f[r*}Y�L�9U�13m�A�Q�\¬Z�d�*�*�h>��\<6G�M�H��!���E�#�2�.~^X8'׿�����qсר�ã��w�"�T)�2�rP�ᡇ!�ܯԤ�-ͅ�$O0�D���'�7Ks^��#V-�ca�z����NdI~�G̍�_vʒ`�1sk���['�;�kD�І��*����w.��p�"v��~񟥈����n�j�II9���G��"�͑®3���B��C�f+VږJ)���\6����f�t�����y����"���}��l+E \# ���@)'��k�|���A;���\C4�*��8y	.�L�^�<]Ƴ���z�?g\J��G�K�j?�g�t�:��J�n9��%� M�C��K��~d�rr<�髈�B���*��Z;Z������Vf�&� �@�A[L�Q��l.@���S,	svL�2poE�4C�!έc���4�H"o����W��6-��8����=����+�#�Z���N{����U'���(#^�r� C���y�PJ��(��T��H�0�#�`�}E1�t+���K�N��[�C�Qr�w��v>�@b��!>�]�<1��V$M#��(�5��3�/�������\�}O�I-���p`G9" LIn`�TF�J#��לt���%fi���C� #;~6$�_ͧzj�t>3���8�ؐ�NV����dM�R��{��l��=r�7B��dSh=��Hu|�ȋ!�SYz�[ 1C��P�yM&����\A����_�0�'j��ܭL�%NηU:�[�w5_��$�țB�*l�$4�L�,�%fG�㊲�Tʤ�,Q�.}Ԓϣ\��"t�=��il'4�R]��JZ� V�UԦ�%6�,��Pێ�l:O,�_Ք$��ږ��������X͗�v,#>$R�ub��
�+�o�lJ@������l>M���A�)�犁�T��@!�l===�,�B�^��QH�����8�ԣ�`�hg���V5��R\MG�Ų%u�F\�\�y�����o�k��:��&�u�\�z�u?�K�=.�ƾLK�Y\�黧��u �%�����|�?�B2Sg0u�Z����V�z��<�(l��\zrd��=4~^ xRǈ� &��I��-{Y���omI��i�b��T!+@bVU��W֯�K�Vaw�q]�-�;�/�s��dܸqn�DX��/V�R�����uݫ�`И)bf�^��P īV�Y��JI�Ш�rmm&N��<f�X�ZQ��Gk&O ��ջy#Z�[$������"�#���8��\{Zjb2��|9���f=?jDt�*����KG5��9m��
vGM��mc'�X�
�yE	2
�ܙ��iI	o��R�O����!��vx�֮]�M]��Z`H��P�bq�M�}3s�O����n���)�D��0L5F�g;�J��Jv�r���$�țW�z�D��S��Q�K6���*HbԪeQ��zz��K+p�����/A2�cR�kn�Q�^T�͡��(%&�żb�K��_��n���� R-R�:0��jdŦ�4G�VK��8"��e�q�ޏo��j5Z��r�d��������|"�G����_X�7��z�pͯ1{�,�� ��.Z�9��r����j7�=bX����{�̒%8�m��?�c'N�l��ʊ�*���vZj��>��9�v�i~tP��}�,y�y�w����e����a��F��S$�h���@�\V)u_*�0ph�-Z�i�&���_���&J�0w��kD�D�j�_ݟ�U�?�`,�#����˱�g%Z��%���{p�7/A��h:�Z�h�PŎf%�H"���esh��݆.�J�)?�R�.׏4K5���J⩸��P��xbC7Vn(��@^]�0�k�bk<� ބ�k����c�!�p�7���qԴ�1m�0��������#WZ�����2�|� Z�6<�|���]����:4��XIjdlo�ۛ@��' ��6��;�w,���8�}��o�j�)�X�G����_D�)pCI�c?�a��[,b�p�#Ob����~�7��FlǪ+X�ن��R{s˘�϶�-1s�t?����3���q�1Gᜋ�����9���1u�8η�J��uL�+�q�/g����G���	��[�����b��e ��q�Q*0�n���J�W&PS�A��
��������0���'>.�s�e8�?���S��)��+��I$����j�ki�5�Tyzq�+�z�F�>�e/��Y�~���E���e���;�:��+��d{LP:���~to+n,k*��̯�ۼ���1�&�qĬ��'���6Hr	MaVʿ�!����D 8i�\�������p��F��B���t�%���M!��[����C��S��#�Ә>~�;��GnǙ��8<�w�w���|NR��x&�?[D���`#�������?GX�@6[@��I�h��'�ǋI�k���qҩAznah|N��}]x�ч��k��L��+��5̚:Yu��B	��'"�l�4���'QY����9]�/�b���h��}�k��זP���Hd����V��S�_!6��~ _:�K���8��g� Z qI8�ݻ�b$�hId�d��CYy�q�x��s�l�K���v�w���w�/�z�ހ�C�����\��b��ѿ���I���D���!�
�XI�;�?܈sN|7���S��)���#�KK��0�>"6��(J\E x�c�p�#`'t�5�1hP��Ϩ��jiW͡��`:Ĕ*I�gG�B��W�{'Vt����%�4�����T}� �N�Q��뺁��\��Ģ��b~~�]Ȍ> �L+�r��������|��`+h��U�&�ږ|Cuf0�k$ ��%�~��cx��/�w,{a	�~��f,8�4��}��D�0#i��x��]�`�r\J�lΈQ�8z�4�����*@ M�sYys�s�L����Dq�*_{R��A����&tƋ7ߎg�}g��|�s��W����]Wu-<vߧޮ�,��Ų-L�tB���Jh		BI���%@�JĀ�������]�,�꺺����?�\k�{e��>I�;�O�v��k�s����q)�+5�Fo�Ɖ;�yaL�����hS\�]'������G>��ݵ���^��(�ZRpae�ѹA��S��QT�)��j�Ku{B�6A���0����I�dĆ�%%|�;�b�k_�/��u�<l\�\ P*y%vw�7�;�ށ{[�^s#�s��(��7�����ٛ�z.*5<���HH�}!�(?if\�,����$�wJ%���p	���:.����j9�rɥxʦ��r�z��J`�к�4睻���\����ߺ�I���hK?�)��H��[$d"�4��s���C��L�8��I��M	��#q��!&��U�ܶg/.��a����k�z�Z���e$q"�kP�Dmx�9�)xʊ��:!�R*���D�����sɢ�hw�T����B�O�ϊ�I���ؠ�BYrUW9����w��������#������NCo�Fo������]nF��(�g�Re���4�?�#e|��ox=���Іjmռ�D.�J��as��sz��J7ٻĺ��%&F|�p���-��(�<��}r��rJhC��*���|�c��i*y!��R�_�z%���v���,^��3H�Q��?.�0�'�G��4$�E����0�Po1/&FC���]~��t��Ø�R�A��r����mbo9�+�����6����v�&q{��.��xM,��$���'�=_�yW����Z����-��C䊓B�@��z0�5�uI֖�ui�L:���X�I<_�[,אv#S�x�!Z��]J�gE�����������J��-o�mW].շ�����qcǮ�x����g��0�lR2H2hZ7��Ќ�kԂa��,m5��-����Z�N�6<n�7�G�f�$��@�6������9�-�c!��p�7.©o5.�̧���}?V�Y+<�(���F�W�7z�7��q̙`�"l�G^.,NN�;w����3�6#��h�:�)��3Sbh�f��(V�iK)����$��1f*!��L6�SǕ�\b/�W��"f�*_���!�XƝ�wag�O^�Z�u�(�}*�H����A�����`��������Bκ?/r�rC���J$-��ʶ��b}T·u"e\���a��Ta=�g�����0m����ҿ~Z�<<�ED�X�����C&������q�����t���=D� �zM�l�E��*M��X�jc`7E  ��\��Z��(PQsE ��028�;�=~��O÷��X�z�<.�P'�@��y���.$�M:Ԙ��>'���8�%�i�Je�@�	e��@�NL9g+�@+j{w%���̀ž��FS�y��C@pl�,Xt�Y0ԏC�ކs�n����\Stg�hB�A�7z�����v�ʕ�ubB)��2�m�Ri�ۢ�a��*�{�/��B]ܝ�	��Tks�Q�r�ؕr!�T��
xr��sDi��
�V^i�X���˿�T#�� �H3��M��j���D�7ܛ)�%�9�D��rQ?��Ѓ��2�DH̆�Hs�~L�YFt�HXʯ�t��ȑ)lٲ@_E��U��V�n=��n��^"l� z%ro���7�B�	*�fH���QU���$��Fft��YD��b�{���4_[����T[݇�-4�	z���]�N;��ϗ�F���g�$������ ��6C�mF?ۮ'cQnan)ͼ��l��sCϱň��G:Uf�B ��}��0L��<�{��U�n��˪�1J�G@��=��s�����V���8��q������Ϯv'g.���Mt���7[�Z0.Vna�3���%�qx"��Z��0�!w-���ˋ�1����)�E��Ual�!���1�|3����Y��p��5�A�����d���Qy=��q��iH�eXm��]��0�,�1�A"Z��u�Ã�%�:\���ӽ�J(<�V�=Wg���TJҁ"�B�WcS�'V�n�Fk�uڨ��*4�����Vfަ��*���X E�Km�l�/�G���k&��-������1ܨ��Ο?�^$?�� ��ӡ�>�*P��Y�F\�� ��k}�g���^�P�jq_$�Ͳ"1���IAS٭̅�����A�iI�>�g��ο��[�l��Z ��Jh�3��Mo�Fo��A�Xx���Q$�J%b ��y�
Ae�";R���]�e� 	;�V3�=�矵�J�8B��o�~=�a9�_��Q����zrB�F��y�V9K)��8d�TQ��C��l��on���>=���
V͙'�n�Y�0��fr�����wa����Sq�K>0�[��K�<?f�r8�=x�O%����U�f���C��Q�) ��ӬUZ���p�0��Q<v��ظC�FVlb����k���"�ĠM�gzf�V�
P�kSby��Mizo�Ǝ(�j���Çh����K�8Ni��	xˮ�3�º3���7k)+�}&Ə�������qR���KMő��;�֩ٚ$@T�.��D�֒�&�Sr�g��������]��I|G�bUh������];^)og=R��$6Q1i�ڏ�O]��V/�����xY���P��r�r���}���d�ͭ`�<��U��c@d��_���$<XvaM�p�@g�4_¶)��� �c�h�� �y���š	�gba�6θ���k�\U���^:.�q��f�o���K�2R�>�$�P5��s�H���Lg����T	����ꆇ�D�FG���}��	�-���j�uQ�[b�!��%~U�s���i�#��t����rA�*�����9S�ؤ1i����'ǜ�W�o��r$6m�� �F'�T�0����<�����_Œ�a�U�"$n$�U���ąU��N&ͧ�j� ��~N��DuK�W�£=�^��7z�Q�=�M�7n�.�ç�X@��`���/��K J\X'�T6�\��l`!=��5+`7���:\F �a�9@��O�\ڟ��r�'�Bs�Bނ8�T��M�+,B�}�8f6�V��o�Gi�n�GQ��X'8��8��a��X`�����S�1;hq[��8!s�&�Y���enj��*R�U|�U92d��M K�as�_,���b�Յݧ����>=��u|[�.�S�o!�g��]c�{z���3J�UBXv0���N���~���-B���)���=MC5m�ţh������Z>�4�����l�KS��nܠwD�3����`���0ͣ㹴��5�'� N��W<�� w^v�N��L��"�ǀ��"��1υ�����-�k������L���jO�U8�^�|���6,�i��&�V���jz~��&���?>ez��ݻ�q�:zX(M򅻻�15u�N
j5?$f(\L�?��%�7?ֹ�ry	�2cM3S3�>R+E_Y�+��w �]w+��013C6��#)[�Й�0�ȴaIi���U{n��[��@�Z��h6�
E�R���j�%�RD��d!a[�C�aNM�y�y&J�w?4�K���	H���J;ai#GC\�M��S��R�,�#9���ݖ��3�Z���&`���r���JU��Ó� r�"0��"3�P+��p�u]i��<p_��Gq2�۸C+F�ܚ�Dߺuxޅ�C�����w��e,>i=:�MNuX��WL�2X@�֛ �i���<�vO�(>Ұo۽�`o��q>�{&X��%=˺�"��bM�(E٩ h��T,8%��ˊ]���O]��5{GG�0m��6b���isK�9Z�531�5��ZN��|�ץ�M�E17�!P�󡯜O�#�%���zw&-\�jDLL����(��F��gPG�J~�ڝ����]�?��^��p�a�( �ciu��-���^�0$6DL���I���<qQg�7����O|<�8G���sW���%Ra�<M_�/.�a�ńm�Dhۥ�6�C�(�T�6�p� e���\k�S���ɁB��?��$��c�����oɆ�I�)C�$ ��!V-D�D���:�}7ߍ��>�NOe�e:;������lZ�+p�2�-)�o�D]�G�?��@�0z����Gi���i��|����F(��,B69>��@M�4Z�C߹���j��_{֬Z�CcG�t�]� (X`��b������� �"�a���t���q	?z�ĸJ�>L-�Z�yzl}�>ڀi�f����}��9��6V�bҙV|�@9���b��_48 �ѻ��Aid.����"��b"��5��Kt(�jQm5D�]�2�=�����s�-/H�F1�e�C3Qn��s��*l�O>�w�j�G�Ya'&vۑ��K�z�o�P@.� ����@�1P�����|�L�n��l60���:t��
�VD'xb2���x�k^���n���yd�6�1gx.����f����v;֒�]{�|��1��d3TH��2v�7����^��T��re��6o�R��d�	��ٜ����{oƼ�;t��K�����������*���}��m~�$��7�u���ptU�X�X�#��@�}�>}�,ZK~�P�!������[�1��YI��T"��C�#�T}����S_{��f�}uL�gc��al�7��!��cbl+!��Qm����a��T�%Kы���5-����'��]A�:��f$����$�({J� &�x^n��Ë�p6m��c��]�ì�es��Lz�$|B�]Xҵu*�;�V����%�Cjy"U8Qô���:T�ph������w�˯�g^'�P��d�D�
���?҅JR��Af�Y�[URmY`՜��*�N0~x?�-ـ'�ڀZ�'�H�@���n�M�23\aQ��6!nU��}��*�*\y�8*�h���͞�j����J��"��@������w��R��Q��
���WcŚ5�􉛮��W��~٧FC��-[݌f��/������{�7N�q�3A�k��#F,z�m�\ԑLO`��A��r�4���:�� �<,�b�
����."��=^����������d��	0�I�XYf�I�V����l�^:� .��O�ͷ݋� �� �P����	x�z�1�	0c���z&RUb�6xC�s$RldH����|T:��g�Y�ǜz��ص� �K���z�q鍷��}G���蹞(�<���2`*�_���>�[o,�#���|� �HlT#���@s�ƫ���0�,b�ӭ�@{�#s1��.���_��Ϯ��J�X��oK�<�D"���As�W������8�A0����������hO�z�T~޴�>�rüe`�R�C,��Y���b��F���(,yd1��{��Ε�ժ���4���I�%L�j>@@�^�܁Ũ�e<�̵�s\�k?l�.!F�����4�Y9�Dȕg��G2u,���@�u�$ <�����n㶟߈���0gdgm܌����o=��Oqw�A��QÓ�3oi@)ܓ�*��ٿ�43ϵN���P��4Y��L�t �,����W�1�{2b������"��B�R@�'t�(��Ӽ[-TO�T��_=c�Qy���{�7�qB��ltI�Z���PU�$�
Y�0�?c��~p������op �F��ۤ�72�v.z���p�%���_q�G�D�6�Nga��wߏ6�SgQoָl3܅a�>��q��&b[�l\�>(.��+8�?���hʄu�$����Dp �Z!qaI&�m�j�g'	�ll�u�0�|�5�/XJ�2���~��񎗽
+����+���oB��ۗYpS�@ʑ�sd�����J�+}��L�31Aˋ�����vW|��XJLu���дx�J,ظ�[Va�)+p�E��?��!����RX0�%���2����K����8��1A#��%�~#�/�~��QBӐ<�lH"���K�iM�O�R���U6�t�g�]	#h��� >���A��&�,��o�@�Ԟ��*#'��s%#=���\������gVN�����0���g�W]��c��@ߋ�Tp8�ǫeD~?��R++�R�<�Ac4���xV=�,�4���V�[�B�o@�rȫ�R�_�1*MUn�0[�����<��*�E�41��Rǒ����Ų�2�LI��a#J��|��[�M�_��XIřc��q�شl!�;�*�@�\���b.yB�K�z:���"�*N��L�O�(��Ƌ{��7��bbjwx6J6�嵧p���#�0*e4� q�����^���F��{��1p����Q��J829�j���T�Jej��\{*�Fo�Ɖ;�)�����B�X�zT��7Nv�03O7V'R�D�T�i%�6��~<�Yυ�h�?���_�VJX��(B����[�Gl�%��D�ڏmc��=Ց�~���,�eʳn�N'Ոf!����oy�v�guVdP������*ZtU�my�4#q��ze�AG��ى>6jh�.<q� :\��Ĩ�9�FB����`�½ �k����S�ΰ\i�ta	ݻ �B�D3΁%���rJHb�G��)b:̑�}84}&@,ӑf��iI>�G�De�rt��e���5 0��(�� _��~>� ؙ�t~��{Z��V��輶�!�p�ٍ��jI�Q��~!dؾ�Dk��<L�O��5*��74gMW���'�;��wl�z�V�������2���Q13a�����,4"i�`W~nb��cz�{�7N�q������M9��>53���P�,]Q�	S��9ڮ�Fk�6)e/d9>������aC
��Y��a�JV�owP��p���q�6������цX�X�H��Z��̄��f��=rE
�R8����3g22[�r������؅� JTJض��^�4��E�h-d��K���M�s1��f��r���a�"��=u�����E�Z�]=;��p�����=!`�����*)� .1�� ���*6��oc:j"�����ԕ&ys6�ϕ�w�١�e���:�Z[տX�d�Ф��
��d�E�~���a�vH`�w:݆;'#��u��簾�`7/9^�TI���>Zl��.:"�l���B�ff�_)��m��5��Fo<j㘇CS�(=7����	t����У�z�*JH�\M�� ;�[��f�v�'ptbCĖ�4��|����V`�cc�`Ǒ	L9U��,��9q��>�B��`�&�9+����m���+3��X�3ayE�(�P��{1�=v���ML7ZhҋZ%C�@Ō��X���l����`&&#إ>��/6H�oҬ$C�I��8�������,f���U��z�K9`p΋���ա�6��q����1g��`3�9˗a����cv�,�>4�I��d�'��X*6� �*`�2��T;����C�ug1X�"䜪�� �{Q�=�gm����@�l�D`�����0Zb���8q��.��h����Y��C�}��]���j��c����q���ɪ=�3j����GoS̍��y�����#U,
����8�X�1k(y�8=I�����@�&�Z��$�C;���1<�q�`d�L���%�������C{%b;"���ŝ{�� 3,��ԁЮeS⛧5H�[��������ի�6hq3w�#�bhː��Oqgv���{�^O����}0K%�q& ��d�F�C��:XD�:�#� ����S�z|��Δߟ	S��D�K$)�;��^�'&�w,��t�8{��~�5�_�C�٧W�޻+�tF������-�A�]RuE1��
�.���6�����{ݥ���#�<]�M�3q�a3�iy8� �<���w���OPF�+k�>�n�%�}������{���@?��� H�sh�E(���J�D������'�8��ƭ�c:,�Ae���r�T���A��R_F�!���<~uA�Cc	^�$����H�*��eg�Љ����"��A9�B�uM�8�;1|��:�TϜ���]�
�''��R+���1�e�(�7yS���>�VO�zV#zh׽�}|?�LO@-��󶞂��q9�]{c��A�}sQuk�p9����7f�i��[�-�1�����sU�bg�f�T�#O�@�u[@h*9:3�<#CKp�w`���c�e��<�_+-&C�u����������q�x�(����6awy�e�&��QE-<"��9�nS<rt[,e� އ�އ����EKA�&g�7I �VG!�El��q�Z���}��IZ���rx>��~-�����wc�w/ǆ+РC�[*�ƌc)��Ŝ���r�O$�i�0�7z��SR�1���좪�`_���T2�pRCK�ebF�$�=���l���R ���9������!p��	;M�L=q�k��K" .���ǅ�q�P���4�g�_+�mu��r2�I�����&%����9!.�ߏ�����0Ņ�UzZ=T�=w>�/]�ËQ�CҤM�6kf*V^�U�"��|V�j��˱T��V���
�0�\��F,)�;)���>:5�Զ�ЁQܴc6._�u�a�ehp���C���<���r�����U�U�c��V�����'��;�잼�w��l��*A"�ƌ�i%����=w���A,}�+���f��Rm�0�5�\4�_{�{q��e�+%���@�1��Tc��DZ$���8��1/�)o*��7tU�a	�q���R��R��Uz��q{C�+Y�L��1:��<i�&�H���/c_�`G#Ɓ��&�o~�����TAæ���9+[LvS(�X�P�δ}��v���M)����Py�b�2C��+�O�M;v�X�p���^��34=�o�����u��Ei�r��>LM�iJ(��`D�270�e�no	��|?�� �$�����gʅ�� 8����b̌<QMiӚ�}}����q��6������I�w�]�ݍ��H�:]ģÅ's�Djb9�M��*/������Fw�EaT��l�q��p����
�6��=�Cz[r�/�Ѻ�>����ߤI
`�F�_��5�q����+~�u�#��.M�ҁɅ��b��A��:i�
�r�^���{�7z��ǉv�n%�o5а���hS�v���#h���+U��4[�}��ϒ�X�����K��r�]���n!@�­��f�A�X�È+�q�aZ��1Z�
1�f�-2O����Y1;�@�!WGR��N_��*QS3��Rm v���,�~�����L_B�	1v1ω)Z�:�s���a�UzN�ખ\�L8���ZT����'��z��Fvt�4[�fٹ�b
�1jb�Ķڴ�)�&v[�L�;1�{~r�0Y���b�
�С��'��6ϋ�b����D��`j�g��B>[�S�+ן�ܘaډn�WybS,���6������.�<�M����b»6j�	�EG`BX�@���%l]�9+�$� }����RD�"]�s/'�jɺ%���Fo�Fo���W�,�H��yv��B,gń�62ިX-s\�Q��E�'Ǥ�u�w��:�*l�?qS7T�Y��i�:,b)qQ`�q^-6)Ra,�[�#��*.��Z���1X���c����¯o���8C��1�.�r�) �a�}h{J�4f��vmN�n��{L+Ӛ��$�qh��:	��P!��i],u �jUSX03�<k�vt.K{�Y�-�}G<�hI�`(�v %�k[7:M�*ea���օ��Pƈ�X�W��F�Ė��S�c�Fn��y��r]A�.b�le	5��	��$FhƩ4�3^�1�!����ڦ	�8�z�i�D��+��#~�LV��{�9��������)�
{�2u�*��a���3��ǟ>�,L���=��5�ZT���#}�ܞ3�:T�(3e@>�lE�����8�L�(�/�
i�΋�K!�@O���p	m>-bns���X�S|¬Y7|�|�̣�̊��0Mr�P7GD�|�CT<b��2�f��`d.m��MN	?�-�sQF�adpSĎ���js�{�3���:+�x�����]�Vn��{�T�$b�=� ���6<iX/�)5���M,�#��!�h
^��Jbe��p����7�2�e�n�Z�`"o�ٚB��=5����9�v � ����z7����*�G	F窏0ղe��F��#f�B�\y�2��A�t	Y��u�@�T+#�쀋3ø�xa�*�F�F�Ç����csC���Z�J?(�{���h���z�`��/�$�o�6��NeΪw3��.<�{�]�c;�mc'��ƍ�۶m4���Ic';hl��y��s����k>�c�1G=&�],����a��V�"[ʷ�ԯ
	Æƍc`.�K@����Cۀ�i������z����:{kI��!�^�_��5o�1�x�ѠQD��>�+���4�%�:O��Jv??'�����U�(�Y�B�2�m�eB!�����n�����B&���/�4Ⱦ����%�\~���UX�$�K���hf����J��?�_�vVL,�'4���f;QS�S��s��3f�gМ�а���[�K{w0�u����BΚ_`��]B���-���G��(�k�l�z��e���r��Ko*�G*��!+ �!UWU�d*ģ���ё+k,��˂��=�6�@��n
i��>xo�h�J��V��@��|I������SuϨY�d�����ȇ�vշn�X%����]ב~V'4�>WG���4&����c!EM��+-id"%���}��9EG�d�{�E�I@��7�N�v���]�C�s`������3#0����v|�3&F�`�n,�bS'��%�<=`���<L�!��ƪg8�=��V2R�3M�����C��~��h�/�qJ���}l�hf��}�h�$_�2��:ڽN�vC��v~ņ�Β��ʥ�{����cTh�|�s��;��bf�D>M8�
%ݩF��K4� ��rM���Bt���V�hb�	�@jg�i#��?���_��e5Z�p>��_1j�低�#4�1@�5�6p�=&��j��fow�&�����P�Z���1q���X:C��c�i0cH)��T��Ewh�Դ�H�ZA�>����5�1ceZ]��<��
�N�����:��bFkH�Q7�s�^���~{Ч��Q^�������NFLe{ %N�N߯ba
�S,]s��{��YZ�ˊ�8�^6)=5�$����@�}��3����(?���] ��]� jQ�J�*E^ȹ�jSoŹ��)�f��V���<�v]8�񰊒j"�0�,Ɍ�O6ȣE��n��(Tk�N�e5�`M̈́���:4��p���Y�["���pqz�>4{|�iI��`���!f�������?�ׯ���n��O���
�Q�$���'�k�e�j����qw즬� �ۖ��ʈ�ɺ�`�Ŝ<�N�P=G-�l��|#���z�~��D\��:pR����!,l��F6zD�y|Q�98��Np���4��3��iiiXh�Q��@*ڬr/+�vg�,�8�e>Z!Yk��K��P*�R��u�~��'��Wȭ���$4��1��� ��e�Q_|���������|���m���.�2�:�9���f��g�"���Z[�v�,`;\������������-N"�C�m�Ӆ�����	7�u��ëe�[��b��Ȑ���?�aϙЙ:� l�kJۈ�S���f3B���ey3�����@���E�$!}�-W�w��H�A[��^�5��u�N]�Y���MV���b���=��K��P��fL����VC�>C��2��q��ݨ�蛾?>��oMG;�^Ȃ�'�"�IP��MG���X�!C�����*�:�5������:�a�@�&f��X��HD��)��,b�hfK�_���{̹6_��Z�paV�Ӆ�d4;d�;�DE[�	�<��ds>E�,��!��w����nLjF�s��H&N6|��\1�2%�����Y����u�>����^����f������n�s��yVS�7j�q�X�4�[u$h�|@�����6x��<
Z��Ȳ�^���!]�N��2�ȜLt=�PG�n�!/{�=�������V(��O�A�db�� l�l�?m���~��G��ij��[���(�{����!{�o��y�{�H���C)JY���FY�MM/=D��p����/��]���S��`�fwe8�ߗ�0>�#�>�~[�1,8��K��8D���"aDk�S��m�B��{��p΍f_�]"�B����F�=�/h��{��R�p�+7�dÑ�s�־���롈 ��0pEЧj���jPb���]����U���X��%T�}VR�o�b�،_5�
���e���ȋ��k���Hrd�M�e�
98��]�/jg��ܣ1x^a-FCh������U�C�����Ǚ��L��,�/밟���5�*��4��*̤Z�X�������-��*�F5�0iO��e,�;*�rUR��m�DD�r-eJU(�wwPP�6�]V�]���"�V�jo\��2>7W�d�)�	bw@�4�+�֮�D�sJ�{�]T�nC��L\	=?�#�!�)�!%��
v)�������/.a���~(��4ҔX�F��Lg( ��Fr��ê��q.C�q�Jɥ#��n�zF���	E��V�P�R�g��t�HFI����B�_-�������Ic����]����_���Yyo�
[u"��u5*�,K��?Kgb3H���stg7\$\����/��GL�z����[ӫ g�����y�8�B�H
�s$�@�Ϡ�k����T��JA!�����\���%�I_h��l�#���*��ɻ��#���n�۱AH�%7"�>���1�un��ڂ��k{W����Ð�nW��G�
\�*FT�.$�T�G����!hZS��
��ԕ'j�[�u�׃�ǒ�T��lM��ѐ����*k�_�>�l귰8���ö�D!��S�W���7yX�KX���p�CY��k�{��"��XS"J'�����.�Z��=�9
�i�g]�v��s�Q� �r�%Q�u�.��;b��t����b�Ūr����>z���>��!3�N�ȡ�@x2��h�1���za��}����j��t�-����V�)���@DOh�|��"�a�Ӄ��z�s���Mp֒9"�⃄�<V�X��!�i��z[�Q���:Gt1#���1#E��#��=*'Y�{a��(.�j�=]N9�@�I7Jt6��t���g���3����|����iZ' G�/C������J�k�a��8j��3G�uV��{8�ZATe����Ý+��b��7�#�!^��g\L�rdhk�Z?:#�O9Ѧ��5"�~�G�޹y��D�(W륨����O(�S������Z��u9,�[��,=�g?��9 "-s�)e��0��˂�x��H��Y���}�y6�g5�-�ml�?x�E���(�1�)���^�J]^��7R��b`_��I��3�so��dl�#l�~,��x�U4���bzZ��[�%�2��n�P�q���899��'ٛd]-6΄�rT݉-�KY�؟���O�����x�����4%rC��: !����8��Y��(���ӟl&v������,���U�<:��'�?�{d���v���ń5eu�V�8��J�����h!ڒߗ?���K�&dN�n>r�.�y<�����4y��G�ҭ��)�4]��D��=�?�R3����@��	��<��w֚��Ѻ{:vTB��%�қGf�t���>�Q<�r�L�N ���W~���p�?ax�1�#a�X#�E�W.������ιKIig��َ�~��%1�D.����!��ؖ�y�Ոd��	��"U�S�#ȭx돑�=C��6N;���Ũ�k�̳E���J�RG�"�N�Tv���/p��PM.����PTtG=)L)c���=m \��v��!��eü�(�눟�|o~f_c-GQ�Q�j�C�b�)�s�������Ɏ�3?e�j��`�M6Rj�os!�r��p5'0V�V'�=c6AsZ�pm�������%�2��<r'z������q/���=��MBq-�/���WPx5z/f���U^�af�ZB2�ߤ����~	81��J�Q�ښ#@��dE������y���B��Ԧ?��U���Ӂ�!�����c��q
֬�>
�(g%�m��	��k8:��t�w|M�!�ҦP[�������ڢP��1�`RY�N�N��Xr��ш҄0am;�#��-T�
�*?֧����j�-{�v�uW9< m�A��ZP�`�Z�^UA�x�L�3IY��.�Sn�kq�e�d��پ��)p�rͰ�C�++ըΜ�X�1�J�������S�Rա��"j8u����_Z��u�֬�꣑���̝+N������iZ�z�1B`L+Ɍ&���)���#�l�>!�,^=�6����Zp@�����;�q�U%u*{�2%��7�F�|9f��7^� w��T}LE���N��t���NDխA3zkMWon� ��@H(e���m>� `D ��]e�Ey8��hk�����֨ˎ߷�!0gG0l�.	!Z�:�d��4B3Y#}k�'?�&�}D�ޓ㴋�蟍�~�Dݺ6��V�[V�� �ԫ[��NLv������������^�"�����J�����l�6�8�����c
$��AM�GE񐵋��G�5 �	��F.��+��hR,+�������jJ=F�&N![��vLC�6ν/?{2}H��Y��v�g�5��#�¬�Z����l.����^�^�U�G�ڀ��O�OҠ;�m5�_7��%���t5>!�;������o9"j���67?�h�C'�g��z�h-�k:?�u�.����6�2s�΃h�ւ����E���fɚ}�cJ�Y��4����!�i���Q���Ք�p�����bF�ة�a���7�7��%�B�S_�ԣ�S`� �8�������М�G"��4�G��x�y���{7����'�)qA��/Kշ,XO�O�u����Cz��)���I�����_L�N��6b����_���>_n�M���JCf	�uE�>.��G��[-+��x�}�<�'�Ї��u��W��H�EF��j��1%�9�RJE�^���H��i������x��7Ww�^��>�F��Q9���Z��W��b#�3�O�MW"�n��g�eJ"�	�H���B�G�ӌ�d�"��/��pa\�R��b�e�Te�p^v�	f��_w�� 2,U�G}�@���#� �7�w>�q�,2-�o��l����gȺ���(��m�����>Ve���3��K~x�?���G��M+pJ�=�8R�i���C�}�}�s+(���I�5@�!ƤȽSJ��V�G��8���m�*���+����xd�jt7�@��N��fX@��py\"�Aބ�Û���m�;a���(��C>K���]0��#�*�_Ɖ�����P8�0�D�h�К};�P׭�s�/�G�.1~��>�&�O*�v,Γ=�8�٬3����(�%�
����}�<�R(��ppP����Gdzys�F`�W�t9�~��M��Rh�Z|v�]��y� �\m>:�f�K4{�}Z��]:�=�Pp�(ũV7����(1E]��ʴ
WD��f�r5x���k�0�9NI����E/<:�N�8y�J��q��V�ƻ�=�<0������o*Mf�&�F�3mi�t�?���ֲ�-B��mh�E��&ʀt Rp�A�^���^�/�u��U�+S��x��=A}ђ�k:�J#���E���9@e�jBt�iO�ӻ4T*�u�����*R���<������а�c�Pp���%�]�	Ҡg��c�=����J ���&�ݔ�E�ؕ�q���wN��9��Z�k���k� ��� ����z�'(��2��G�'�P��=�T[�oHFW��w�T�~N�̳�?��~����_P��G�֨��`��lH#��j�(�N�<��iȸ\��+P�c #�]��b�wx���^GPw�4���4�,����1�o:����Q��4?��J�8���@�1���v;r����$#��4B�E��ϫ�R�[�2Ƥ�{|��.�tH�!���{m��	��"7�N���Y<���zDlt;uW)t���Mbe2Mb9 �7)G�C��W�-H��<{/�_�O�T�^ ݒ�I���e�1���.��w��+�A�L�g#�t�ߓЌ����<���T��F.f}q�ۏ)�e�z��2-ɻ�PN��rs��6��`=����`Qc�Tkg�t�X������
�l���^b�E՛ȏ���D~���˩1iD�J,	|����2\o.� s�o;!���6�<]r~D�x�芌�t^u�EJ� =��ؼ}�q0���IйI6���&�1'�S}�u1k�u²��h��S�ͨ��~�Bj��<�z_�D��G�P�����t֑F��?������j�����W��&����'�����2���xHH��%D/H��ז+N���UJM3#��p�mv���v�Zf_ǆ�S6����9h��~$w�o�z���������: �"���I.scI����R�����Lzi�XuE0 ���m��!���]�Ȁ�>���v���w�m�����h6�iS�m��X�D��a���C*+�C��3A�"<��!��f%���w�7���zӚ�U���)[���E�e?$w���{]$� 儂h�zn��l���u?�d2�y�2�17��R�|Ih������ N5�L��]��H������_h�h3�N y�#�d�z�E��G�AXV�]f�Q���Qn8M�f`#�������}j���k�Y�#����%݂F�*M�3�lЙ����6X����L8��F��L��e�Ղ��suv����c�������d���2�|����ON�)�!�xΔ5�.���}|]�+Aݗ�5%�B�V��Ƣ� 2f�������~�a�#���l�n*�i�9�e�U0��΃���/H�y��>_��5���PDRyl��,����t����e��_*Q���J��.O���Л���6������8ح�)Un�����q�KzCl�Y�A59�o��RW��^t�����5�ጽM���-K�e�T��~�m|��۴<%I
-��r���y���庝���Y�~1�F�O��iOU�v	����5:�ګ�P�}5:)��D�n�_���
L��
���c'Ѱ��$�f�7���d�ōj��\�{v�a3�����Cx�{FPos��]�|=�Z��J�������7�ȩGA��)� zq��)s�Y9�P
����/��2��aa)����+�Y��h>�Z�4q�1,����M��/\�k��l�ߥ��?�go�����}�P
�|�W��C� >����Z����� �\E}�R����0	�1�|�TT��Hm��?Xwu��W�sl�C�<��
a��$����7���0zz���o�&A���S�%�#��0�n���y�6jk&!T��ٍ>���E����(fU�!��G�RJ�r��NÓ�Y3��#�8�@Ь�G"dd�\���7}@�I�ݑ�!G���
��vb�I�Pj��L��>�����:g�͒?��CDox�N�6�EyoY�+��3�}&s��g���<=GDw�F{X�&�V�VP�Ǫj�Zn )�f�v��|�ci�}z�<�,�g����pX�����'�c�i3bL�y���|2�DFFA���g(U�ݲv�i���*�H�x�/��O�Q:�ct���:�ث!v�������o����q�����������D#���{x�5�����=z���E���/�0��AJ[�ޡ���K��m/tC�?5��^-�O�íIHOA��>��j�C��o��3��Co v≍�5�鉀n˘ŭw�h�x��2ۀ��v����y�J�="t&��w�}��l�'��g����>���"_,<��D�O�>���ĀZ����8�O���r�~D�I�I��u�s��8 ��BO*KX�1P���F��*C��NFv�(61{�,n=|>�9�=��t�dE+ۢ�*z}��<�>@>ұ�6�����R�匎�I�#+~�@7�2��ǈ�+�R����OY�y��(h�.7�� ����Zll��H���׾?r�YX��I�����m�6z�#�*���i�DEݙ�(�9��I��Nz�æ�׳���i������w݁�jT�����{�|Ȥ�����iղ���l{�|`6o6�
��. 2�����F�4&4F��Ž�󃳫�d���C�<���W�%��q�z�?	������؁�d����N\M�j'Q�u�h��c4j(Aa��*��Pl{m�d�w���c����7�u��&9Dz���>�n
�w:��`[�R㣓OՠDL�%�@������mH��b=;m�~	N���t�{ya�HF0�nѼ��I�K���X�{�G�4!`��q����V|�+��	3
1ċ�E�@�F���g�ǡJn�F�b���2f�d����֍P�����cKyY��p�yӸ��1����g����yt&��j�a�<�kv�� ��_��7x�����/F���36��ODs�n���^_v1�����F�P�� ����z�(��d�#�TN�'C�bKn{�,Ծ�SK���q�c�k+mt�V1��SS�>ٛ�->�.W��yMc�=O����pf��)zϓ�����KC������I�4�$��aᤍK�;9�4���6H�¼Zc�
�ߗ���0����Z���$C��ݨ{��C2T~ػ���ӗ�U�4�X�����Ŋ�cR��2;�e��_[�!^�L�9��nDģњ
2����1
�����ccq+0�M���8O��q}}}���X�(�Ӿ�9��MN�fN�����k ����mI�4$���j	�KC~|���
1��6�~�)�:��\C���fmd�L�_6��8����E�~*����r�;����Ղ��*0\����ɮ�ԧ��A#�l�ડ*�
��1&�����IG�}�w��P �l���<���`X�b-�%fF��`;6�(��>3/��Z_�zU1�5��'vlf���-B���S��ES�^&~�1W�����'js��J��!-K��<���_��$�\�L�4"嚸� �2M�zX��#��B ���W"{[f���=0n�&����c��mM�|@b���C0�ey]���3-]/��d�['��B�I1MAD#�|�#ob`�~�l��o��{e�3:�/B"_ GpC
���,u ��ʇ�{�T2@��>����슯�f?�,-�e�_�P�Bq��<�:4-���G�L�:�ȼ���+g�n�i��5APvt���t��i�Ԟ !��|2f�+��5*3��Ԅ|<���OQ�ɨ"��~�|��fd��������ʀA?����[	��ě�{��J��� �;�����-�f|�ߵe��ꉸ�@���8�e��(z^�Z=I�o<퉔�烱Q$��
}F����?�㸽�}�|F.�<�-1���V���e�WF<�*ч��SВ�+F�"�p���w�+7�{م_
ydë�Rpv39�� �]av��;/`�������L�;����<^��A��bZ��#V�C�=79��j*J��F̝�+?��B	��I�Gfk��D�	<�2t�Em�6g
�:s��);[Hev�=�n�P��	�����
�&������>�ccr.80 VI����paNfЧn������x�؍������ �-�P3�a���l]���]}��XdGcO8Q��+{3%4cr��U>w��B��eL2�u2l(�-뢎���_�9��� ��(�ՁJ��z�ր2%�g��w֞.T�0TL��dk�=�j��+9��x���$���#��-R���4�#� �t��JN�';��L5 �ˬ�<"An�(zHz"6����o�m诳+�S
G��Z%c��@[�Y�\x ��=?��k�g�V�B��"PEGE�m�83l�(U넧~qG���vhEmC�7�2A�#D�q&�~�kF�$��6g[$~�\C�wK����f�&"[D% 0V��<�����U��	�TP��)�;���0O<��V�jt:�t�P4�:B���X>�|	������Ҁ�y3�r�5��o����ϳU9:����`�p�6(�Z��R��1ǻ�z�/EvԗJ�m<��=���+V)O6�>n�݁Y�n
7S��j(�*G��/C�r�~�+R�jUiD�\�k�3�R'E�|���`z��c�f�1�7�z��b|:a_�D��4��^'6�q���c�I7.�����2G�U;�(8i{s�x-��m��BJ�@��4�xLX:
��=��⬗l5D�~����fۑQ�ݖ���|��T�!-��g�_��/�@�.�v��Zk�p�yg?AMi��~G�¤y!�z)9V����F�@�'Y0W���jf�1��^%�?6<2���f)Z, ��V��p~F{����w�+��gΒb��H�í�ZW<I�67�`�B�Ѳ =���ٕ���V��|Z/�xc��r-��ߑ+��$v��rh~ZKQ_0��~9���59�D9��,�������F�0T Dn��߿�Z'���wI`������Hq�>_G�kk����?����^��_���������֝�6"�?~,?�ԇ�f�%Kg��(��ܲ�r�;�r�R%���f�mksA˴�m�uA�w��C��	5sdⲦ�<���O��DF�'c_4o����.����W�ѕ�!{�b5����X�d��W����|�W��a����&�n�T�bc�~Qj�&�?Y�Dv�K�g�)L���!-��kTI�la�'_44�s����̓%5�?�I��(Y�r�7o�^`n�XK��w��-��>�·Yt�Z�����o]n	D�3�p��~��d�d�|����Dgƙu��sze�`���l)j�͊��I�o��#��DB�}��x�^�ڱ��e��q����:��¹3��H���`�H��mًf�!����B&�8�����ċ�Cj7�nB[��Xt���C�%ǚ��<�w{p1��#3U"�M:$�4�m�V��W����t��F�(�����{���Fb@�^6yT�N�}�9�+��b��4Bq���Z�R!��\��+
B��8��ͺ	�߃v�-,��?�~X�<��:��`���͝�d�=W�����hJ��S��-UP�b	)�M�Y�H���xy�	�̘�.7�F�)��6oEZP�`R��[�^�AH��G�K�i|B������	:����8���Y�2p��aאӑ�og�������6nˈo8gt0��4��vXz�ڼ��#���dU��L�d^���C_n��qRA����2��Xv��ћO1��){R2.*+:�2�-xA��N�bi
�;I��t�4�U��J�Nz����?��D�Z�U`<�n͏d��.�<]�!�p-LU�!+���br��Aꄶ��&�s-���������)��̽��j}7��2X=p�<$O)3pQ������(}�71��Zy�pૺ]�{����#����HP�	Cӻ�^�ج\����`լv�i���Z��/���PȆB&,**���~��w��k��FX������v>�<:�����عi�a06oe��M���1���K�?���o��Ԇ�x�xR]����E� �����7��gx�d��t�p`2����G��4��99��l$0��j��A/u]�-[.i�2ǲ��O>�xkE�P��x8D*:����g��sjLf����:��A���]d�>���{�(�N= Z��neܶ@+��9I�9ɜ+����������hJ����xCezF"�z��"B=vn�z�c���c`r���|��MFaK�NK������z\hc���o[}�����1��P�%fT.������J*%K�4�����>���ý��
�ƨ��T��	R��1W�:d
������)B`
�m*EOek�%`wf����XJI'Zxo���*p�@�8�I��)�6rBPa�Ի����E]aiR�EkEmxS�A� ��?ŋ�(��Uۑ�P���Zg�e ��^���R����C9���XN�1!�v�:B��X6��ΑUC������x���5�:<p.��~?8���҉�YŪ�jc�Q�K��Ӧ���u]�����k(����6���zWoV��uZg}
^?$��]�Y߸��j���aK��С�B�T�h��>�egΫ9��3-�^���(��4�,���u$=�;�9\�30X-��Fś���x�Cn�0�-_Cձ������J������aj�.D\�:dt�8빗=����%�ʮg�%d�^�U3yy/e��&���-���6?�W'.��:�6��7��P§�Ϸa�k��Dq7���b�~D6�'�_���	���H"��q�����(����[Na��'�����B,KE��y��w�>�v����`_>�k�.r��	y�Dג6ŃH�[�ֻ}��e%��qu����dJ�txY�NY��#-8�X@i��Y�s�YĽQ�ِ֬��]�{gB�{�խu6���ޗК�X�M��X��b�����5���n���� ��x�<^�m�FQ`SNrM�bF�<Tf�rM��ы�A[Q�<�P!�
6���8_����:���bBUta<7�{�&ݘ^����l�Y�$�p�Iv��[��)�3�� Q?�v�$�`��d��WVk?�^�=�J#b�jx��C�liX ��I�s���
��mz	H�W�����<��g�u�n�1rF|�:�z݆W(��S��Ӧ=( �/\k2�{�⌕gt))T��3��U������c�io�egP�8F��ءa�FJy��J7o���C�*i6G����L�-�b�D�BEԊ�P� ��	)n*-�Uٹ��:���K���r�]�|�--6���	s�k���4�>!)�\H&��o��� �5ڷ�	�k�F]d �RLCh�:��K|�ߢdH�p&���6d�v����>�gs�����8o#��Z$�ja�o���N���y.R<�0�w�Ml�gُb�5��H���s.`��.?���/�>�Y�l�{J�k�͐�kʋe���G��B��!Q�nܷ���3l�5_����X��C��ݡt�?$�󽛾L��wg��X����fYX�f�j�� ]palVs���+C-N3[�G8��p'e�*��2�Y�7���6�]���Q��1f이���h^�o��� ���&g�J����C ���9�F�.��5��G������_u���FzĜ{�)���4��y{�sԨ���Z��.x%t�+gb\1UB����O�m���)�U�8��׾mu�j� �	g�����Q���j��	j�Msz�?�P���b��1a�7Ȍ�}r	J�b����DuL9ԋ7��2pC��Zh�=�_i9�ӕ������ꝼH���-(e6���e�.�-����Z�ϻ����-���x�]Y�݄���Ɉye�bM����@ɺl�I�4Ԋ���	��H9X��yĒ�����\~�@&�v��w"EC.T�t�χכ�!6C]tM�b>�=���,2Q�eb�eZ�di!�wB	uuI3OՃ0���������e'�Z�����?/�D�Q�����D}u�p����(��݈�0Ru.�Э��J�P��Q?4����1��\���b�c�3RO3���⯉�����		�֌TӉH|P��`t\Z�7��� �W�J[�RŢ*��̗V���;��i:v�����0p�p��W�QEU�ى��u���e�o0 �̈���Q�e�\���
��ے�#;zc��ى;~|�K����29�\��+�`�+Lՠ^�;W�i���ë��ɦj��h�s���±��t ����Lij��7:T���2��u|����OY��r� ��2��F'6
�rh�����D�F/��e��eLjH�$�2�ZQ�M�g	�5$��ZO�4��5Hy����B��	��!���b�=X�^����c��������N�K�R!AR�d��?�t�(�H>��Qˤ�l`1|�fO�����72���;>�a3�p���{J�|_Fϊ3�<U��{g^�L��Ӫũ�go"Z�ޜ�rj ���;��h���{P̻c�װ��P��eV��eH��Y�:�����G�Y���*<�u�F�>}�S��X��މb�k�(J$��UdAJ�����]�t��LǺI����"(GN��R�
��$z�����iA�v�B|8h(��&������0fyt��q_��[��.�(%����Mu�Wr��U��Ơ�����n�S �D�^��O5�C�(���xin���c#{���A�F?��h����c��n�k9�s�ӡ�އ�+}�?Ҝy�8騺x�bB���6:&!��譃%a��^E������/8��b�)�k"Ep�r�����c�I�#f����?N�����ߩR��J�ܰ�]���5��@���ֻ#ş�!-�CC
ꎤ�jB���)��(�υ�-ș;	G2�e����=Z�%H>�Y���Z���w.7=U�X!�M4*nE\�S|��}+Su�d<����>����{��IV?�]�7�Aa1L_n���
��UV�9���Ie��3�8�hy�K�ps�t����1��ZЇ����$qF�{[�x
o}s�\��A`3۷{��� T/��A� &�-�JJ(*�����tG\B��� e{�&��}ؘ�e�˵�3��¢��_�ϔ�]!��7i����� �|HZܙ���=�<����f�ޏR5
%�p�2����g�a&�_�+�V ��s��C�K��7��%�kc�>�&��ѧ.FͿjAdgr4��&�TB�.�+���q�sN�G�
$6:	�HgW�6����@t��O���� �a�E�9��Y�d�:�f�S�ʡ�Љ�?z� ���e��-^�4Ø����΅��5${�P���l�D	0�᷽��hrrÎ0��":O�>�8����U�yk;/Z-`���$<� �&#][�
���}0FaH�[�WJm�@�M՞��%'.p�x�)��n7X�� �@Bv�-��Ԝoo��!Q9����z=Nxh2k1�0�Z���ȁ=#��z@C%f���wŉp�G�������F�@-�(
L�]N!b	܌6����r��C$Gx�,���O�J�Z�T��2D�4���"\$��\?j��p,O���]���3=E���׋��'V�%������7����4��`q�T���4NΘ��Cj4�Mӄ��|��:Q���LA4���f�vx%�1в"�o//�%���.WFAws��4y]̦�"��3=d]J8^��c�F���{��$�76�׆�~�8;E�a�ڤ��,�^����>�P�3V�Ft�"Ka��>a$�&j�i�p�k��y'���i����6Y���yL�*��������"����TV�����>ֿ�u�ʳ[d\v�w�JH5����ͷFZi,�T^'����/a;ED(\�s��[,�C8���T�`zt@�2�9[���x��.�<j;�1�?��Q�3�ӛ�X������
|��=m'�z��ƕr�;���H��|�.۳p��+n�<�� �����RǕ�x�˴є��<�;�m��y���,=��s%��*�H��L�Rp\Ͷ�L:�`b#e�$���,�9_�Ҋ��1�d?,�8����$2dѿ��	����&��6�NJ���8�*|''�������G�)*����4.���1��=�=vj��۩L�,&�zf����d�?�`<^��;dpjA���6�U�4b���.�M��9IƵH�o^'r��ԫ1Y��
�B�W��L���,��j�'�_(~��aF��'�PU��M��#���p��4$�/���d�	�jWa���3�
�	�ԓ�Ū:
�Ѝ�z��)�$ܜ�#�ݱ�b#rd+��+����̪�Q�9ݢ�q�͔��u�2�:�����|qR-�-*���ZY�&E���.��<����_P���L�+_8EUM;_-�-~�L�v�]$}q"L�٣�QZ���әտ��V�7��c���`g������t�[��a=��s�x#R����$�@#���ě�`Np�ߠ�>����%n)?)����L��[�Aa���tj�s7�	�%�a-���W�*�e�܃r�4�;ꋿ��rO#T���E��왉VC��~� E
�k�RM��K|�~��F
(n����xc=n�r��9�Ty���)5Z�s��*}��t�g�g�֩��%�(ϋ�н�f�a�����߸��uTK��aN�g(a0ܭ�r>%��&���S���r��k#�h�UcAP���~s]�"'O��?D�c&��5۶m[۶m۶=�m'<�m�����>�=����Z]�֪��v=Er�En��De@�J�2�w Hጃf��r�跹��N��������D�qSɒ���eҡ��� `��;�Ytc%�eg��.��\b���a�K�C���3�%�󫃧����d��c�R��/�l�vl�D��i��n� "9q^���n]��%�4I��R\�xC�4�H�M�d�M+�H1�1T%C�!����_���]�1L���AT��p��s<��� {�ɇ��K��@�˧lr�pL�,P�b�1�,�G�h���Oр��Ȗ�
� 9Ф	'e6��d�z;�U.���Ů�c&q5*�0��G(w��IK	;-�~�(ͤ�ڀ�J�ȕ�x�d��f��C��H�a�:��A��~���&ba�ю�C�#�@4�=4��h;�M��"#����II��f��	��@[եVJ����l]߈�l�N��D��%���F�1,x�4&�����['K�(1��,5�(
�F��$~EyۉE���Ѩp��fLsj��e1�F� Ἇt�pɍawւ�	]C��u�^�e��_��P|�q(Ld)�c��h�(]Ë�>P�İQX�M�WȽϯWOih��N	 jw�
�X�ہ]Aڶ�Gy�\WfK���s�v=?nIU�X����ގoQ#{4;q5�����t��jA�ؗ�IѨ�г?s
������Hi�f�4l AdB+U���?��ʟ�J�,%�V��9XD֗����
}n��6ςk�;��/(�ű�[
I��V�p�����T�#X"�Z拖�B�F��(�ߤMJ��we� �O�C`�]���ѿ�~.{����p�r`���7�q~_a�.����<h��5��H}�i��~D�l`���n$�܈ߘJ�\��t��i/�D�	5�b��"��g(r�#Y ���O4i����9cԸ[���c��^�@@�l���#�{����Y�	f�B��a�I��^��׍
98������	�n���A>:��ړ�X�n� ��.%#�t/�1�Ie�G�~\����h9��0�6 ̷S�.��}K�.���$x�öɤ�	�i#|�ʁ�(�ҭ��K� �֎5s�U��]�Z��e?�#�Vv��.ʩ���G�y�@er�M {�����x���6�a)�"�4�15Aʧ�3���x��-w���e�4�=�)��x��2,ơI�D��3]ՅL̃�,�˷%�P��|-@NM�6j�՝�G�^V˾��:�\�0z�X�H���8@�U���o�9�q0��W>L�`�}U7!��>0�ұ�T�Nྜྷ�+��_c��ℵ�b��؜ơz\�����*� (�nV�<QfX0ǃ�^a@Hv�Kj,]J�"�'4��dA�E�`�Nr��h��J�8����V�w�c����������<�� ����:��B��*a��g�M!
G��@b�5����|�&!Ȁia.���ǥ�����[4���,l>O��u��M
�?��������B0�X&�p�xE�v:��k�p�}��s����s�kU�[gSh�$�|!��>�DH��S�B��d&��:��s/�?�q&F֟�2�NB ���O�ͤhӠ�s}k����Z5��=(��$!HfG�u���#�C���?K�!���-1�C7�T�BLH88���IϛQ?�a�鞇QB�:"��+(!�1%�c��/��E贖\o�x��'$;�k��d�'�
�&5���\:�R��ΗZ�=��������v�wp�lV��!��x-V� ��י��L�@�����.G:Ns�$�<\��P)Ù�hX~��)�	�k5����
���w����$F��\.�TmQ񞔕I���^B��x~n��W\͑wZ{��-�$9�.������ϗ��݉�j�;_; I֘�����jdP5j'�Gc��` ����`������h"A �VD�R�gOR�_�p��ye ���p��'j}	�!�R�Dm��t!��R����J��Fy��U�~&Q?�^�r��Px�s|¦���Yxy�-7�d蜤X�b���$����M��Y8�z�M\F�hq�o\Spk��_���������]���IG�9����[�_̅�^�}v6�������d�qMu&q7s��(����t��kt"K�^7��!�werU�"{_��i��EU
WZY��z���Y�V�8+y=�(�V�������0��.������evU����o�Z���v����5��S�����)�X�1��J�fL�Ċto��i��ʥTJ���f��
%�Đ8�8�*�E����4a@�P�߃~�7m���q�<�5�` ̨L�r[%�r��RL�ʻ1���|?�����}yfl���LN���eM3݇�Ԉ������<Ŭ@�,9�iׄ~4���]eB��*�&Q-y��Lܵ��ϼ��K^X�7�^��e�8�!��zQ)Qm�}�/"������/fA7%��%H��$&�=����⨃� ��|ƶGLC�e�Ќݲ��5'ݺ�,� ���8�ו"�v�̈́_�ߪ{�ȥ��<��s���D+�qb�I�z�*m�y��H
ȯ��9�-kzV?/V��f���h5��q���{@��N�l�e�Z�f�b^ޞe>���,�EW��Y�C<��Y�$��U�*�8XY���\n߽h���i��V^�'^�76�>R�^J�s�.��@�������� w������7֏���"1�d��;Hr��I�P�zV���X�o}*|�Jt&��PM`CpͶ;��u^�S�P��s��G(UO�T��=>|�*.�3�m'�������v��������˶��[�v&�ƴ��<r��uW��,>�Кj�Rt�5�R�J�a���s�<^���}xO����w��a���:A3fΊ�'u�^�Y������w�=�ǜ�~����E��F�C����\�����+ԣu���Bծ���R���8;nO41�x�¦��a�>���v}oꛎ Xq�tv~����m�^��b�ؤw?�.p��
b�>��OC%�m��wa�����׻F��V��Z�-���7�,��C�h�Ɯ �,U:q��
^u��b?�~�s�O(��;u�^/��}��K$h��:�>�c�8�M���U��p�h������}�H
��h�sK�fa	d��Y<7��:���n��A����Ǔ5{�����1����c�(�!��,��Ύa72�I�i۔M:�õ0�7}�����U� a5�����d��]'
�W�ИV�mq,���~j��6|��>�����.�N�v�s���:���z��>U�c� �ݧ���:;�o*0�;4%?�E����r� ���-�@���v}Lh��9�kVTY%Z��{skژ�A���̓��� �&��g�>��Ǯ3�<.7�,��w0���v�;����Yп_����i>/�6w� ��J�'Y��mč����'��<,uyG�G�ĵ�ɱP��Y��d5^��#kW���!�12��R˛B��c���N�؋�yE8�ˍ9����0�V�Y�����чؽ7>2�{zF���A�s����W�ˬ�9N�4�u*�j@�An�Im����v�eaW��GZ�q�a��:��������P0iP�ƍg�,��B���o��s�s�ݛ{����oo4_Nz����s<�q��>˃�)�V75p�� H���k*��9v��5�jՔ)�3���I(������p�GX��u��Xk���i?�p~l��b�z�Ln��ͶA��wu�:�P���o�<i�՚�|8eLM����U�qU~�c��xZ��Y���s`o,�&�d~���9Cۗ��{D������}||�ߖ ��M^��##B�^����91��{Sv�aE���N���>r��Ӳ���ϓ����T��s��-G�r�$΅]�=sq��W�#��,>t|<���ɝ���)Y��f��xW֨��A��m�ߓ��k�ygc�@� /~��ْ���7>����n�,�_����S��B���TQ9֝��+�%�L�I'�{\������S�$�g�23�+E����GLY�%q��77C˷���Sx-G:c�D+�H�Uk�>\e�} ��5>@0��h�#<����P��U?'��,�@ZHՉ� �@@0جWr*P*�]Q'�������:���%����Q�(���;��J�jXq.��]M�����J�t	@<S����⌄/Ӗ�8S���Oí�n� K�S�����"��U,d��=��pd�؅��?���%�Rx5��~���Ƙ��\�tl�'��+l�u�G"�b�F�����K�Y欗��!`�r-�W.�3�T�{�wh�b�������:ҏ�3����:��������	�+�b���V�F��*�[O���?.MO�:�+f�c�4�]�bgZ�Z�>"0��B�=O%��`#'Jv̥�q����{@W,2�D��*A�)�`ҋb�$���ZIZ�7MO��
�g+X��ЕM�X� �p�W��#�G���6�+s;T^�&&Y��䖭z�Zv��~���8[�EQ;��r�:N���~�=��9U�
_�����������`/�L_ ��������9Cy��7�Ft�����"k��5N�#����A�k�s/�9��g�Ƴ�����T/l
��h�R���l~.g�}2Np��p�+��WŜv�T�s�d�x�/���sh$𞓚���# Y�S�[K$��`�e+@�W��u��>�3�9��07�D�f�n���AUX�8�Q���a-�S=&�7�UkG=kE�r}�[�O��:#�i
�$��S���(�B��O��ϱ*�M�Q�GK(!���G"����V�e�K�9|ڢC���$O�Б�'�]g���2R��߱��J�<�n��ڙ��N<8񩛑�҄Q��gӖ{���p��je����sZ��8F]7�y�ׅ�I���6����8����aj����t"���&��$O�t��Z!s�8Z�o���������r��W�BG���w��3�]ؘ�ԠST��J'�]��wPߥJm���Z`;ՂZ`�k� ��=J�0�Tԕ<�v,�C١L���ۑ_�Ҿ��*�p��: ������Z�Jty(Z8ІK�j\`��u��B��CF(d�kΎΚ��Uk�i��hC�JK�>K�� �<�&�zEqKnfq��)����5QlotutElJU�5m7�;w�Uf�M�<$��mKm��B�ɪ���.o���{ROv9:ǊG�N�td���;������Ŕ�Y^}M�%�	���(�Af�F)(B-!c��͚��v,�;��#��;��X6k��vK�k#��q����ڻ)�t�Z�z� &��S#R�YV�`-]�qK�ݹ:v穚(p5�F̣��!b"�ϭ8⿶w�����${���`G��fq�AwտA����wDb8dB����:U���hg�4M{�׃��9���M�S@��oc�r@�:��=�a�M�Sq���a0#h8	��odZ�ZD�W�M�9���oX�OD(k��o�{\cK(��$z\6�[$�{뇇�BO������(�H�C<����=�S�V_ވ�H�\�\�q���	0s��NX$�,��a�!���33c�v��.^�A��Q��a<Y� ���X��#F9��UK	j����#��&�^��M'��h��`D�S�
Zh�TK�/aʸ!�4�@���)ܒ�
e"�t�j(�Lv��D��x^f��N?¥�n�)�ʡ��ڍ~�x�S]Y^�G�*��L�/�P�g��9�È�&�'�Y��Y���h�ŁEb*����$b�}�|�o��̀�8����$7�pE<i�>��t=����q��뮨����;T%0��z�[�e ��Y�?�[qv,s�A�y��s��jl���~��`���r�;5���p�kq{8�H<P<T��֐�$x�g��P��v)��4z��m����xx5eWG�S�%�ERґ���X���	���YN�w��C2��.�P=����v�c��ܯi��]���a7AҁOO�4����@�BǴ4�>V �[|���[R�.�išɿ���'~�I�G�*
�4dM�ׯ8T/mЇ�p��DUs�?�6�_�@	?�@�W&ܶ&�'�\�ZV��74��i���k\�5���VK�d���P�>�a\oG)��8��B��f�g�g�S��+��W�c.3Bs�R�0~�w	�
I��yQ����������[�l�����'�y��i�e��Y�͈>A�}�����3
i�#fV��ښ�[�֌��7�C��<N�m�NF5ݶ���FǷ��\����5O�2e��Y���yv�M�U�������œ~��R�7%�O��q_� ����R#�.
�L&hu��Þ(���0���'��xux��}L�Y��)�]��8�n�	��֬�7s�_�	������Bք9Cu���:�����u�>���0�Y�}����_�Mʴ(��[��P�@���U�.��y���܏��c��gT�QE�Ǭ�&>^ڱ#�-(��>j���c��
���$���&3?e��	\/-�a����w�C��χi�H��l��&@�雏��SK銰괜l���yb��p�G��Z*X*?�*|)����x������Ņ�5��"�Y3�şv�{��:K�7EyX��qۅ>��(���3(i&��.!�J
4{�f�%#�!8V��W�YfA�O���Ԣ!��ރm��]>o�<��v;���΃��)dp�n��k�@	�[eU=�^Y����/��2��)�kU�������njy�g/���o��cU:�}��oQ�F���y�q"a��ٚX���=��HH[�G�?v��l\��B������4/�N�F��H�����U����/����1�vg�AN��f�w��W����m��ѫ g�rr���h0��:�]L���&��/���C=�2�>|>�~h�۽9j1.�"si��Je@K��E�2��7�����"��_�	�qz��F�{Ç������}j����mɼ4�p�%LcNH�@9�����<�t�MR�~gۺf<�P��;&B�� rD���C�@��짒K+[��uZ��ړ�X�i�����E�C	��>�����ξ��v�����I��S�=�R���d��������(;��	�-8� ���-��~���d���qQv��U{�s����+a��´��!$�b3:������ؼ�L0KM�Ȳ�X���G��J�F�K&��B��W�n�py^��(^�y���p����^.~&�����~{s���9�c~��+ x�3�t�Tto"��걟���}Gڭ1ʙ�f4=�k,b�y[}��яԾ@wU��~(2G\�}��v��9����e������,�����F��U*d�ޯ�v�Y�U�
�=���ȧ���~<MX:U;4��IE/���Q5�|�#�������RI�:$�leR�)�)�o?��1K��u���#�'#�0�g*�_U.��9y�Է�m9���}/�\V�<�����=� q�ߜ�2�ecobBƣH޻�k��4\=�B�k�%�������_Ɉ���%�V`�k��#�h?]��S=p��͓Ɯ~Xo�bW]%�M]�Lh�ߤN���=1(�FӜ��v�����]���s3�������s^�)E!��o�IG��%ɶ��-�J+�j�\!Z8�X�(�R�g�YK�0@�2�ۋs�������}o��Q�a�@̫!�=c^�\b����:��>��?�{}�C�=5/�'���� �<�oL�y��Y�,E�2�T� �dg�K��A��
{̛�$�U�G�Jl�f�$TZ
},�s�l�?�����Y�nP&�b�A�� ��\�&?|�ي��;���n�#������ �`���,#NX&�\=�x�to��	�|ǎ�aWY~���H|p�\�T&;Bzm��,�I�H����K�}x��)����J�����D�a��n�\}��<>��y.�8��ʱ�s ��̆�f<cW71��Ϭ'��;��J��~jy8]�\1"F�Q�S�hG˓{I��9 ^Y-�|*�6�&�|��	qoc��c� ������qt~�@�0x��6v\�1���|�u���wa��)����N`���0A/�^D;a'f��H��;�ז��bf�9�f���t��2z���d���R2Hz��X�߭���~2�y��N.�s�����}F�^�[� 	�ޞBz�z���J�Ճ�an�]|@7F�����H��F��O��}�h�&XM�J�)����1���EE5�)۵G��&V�6�c���Md<c�}�g�*߷h����I�6_��D�Nɒ�$=��aơ�;-:�ߤ❠__k���T�U�Au7q������rㅥ$<\p�QD�5=)���)2p���^�3���j85��A?OE��9����\�Wa�NBʑSk�+��9�B��� %s�:�K�S��y�c�Y/Ѿ�_8U����*�n!�/Q�j4��=�e��Ι��(�d]���|� 3���
}��=�o���o{���=�,n��Gm�������k�"S�U8�֚����x�B~?�����C�K�HT���Y�*5�R���а3j���N�� R�I�fE�[4������SB]J�*��?��堿�������W��Y_�q�����l�.��ٯg �~��x�a�!d�+@ ֭�����2�r�l���2^�xQy�Sc@�"�؈>��{�t�^b��V��q�pu"� ��z�H�/R|	�x�vž��y9p������K��ݣ�`���t���V��1Hv��a�i��\fwc"�l$lM�U���*��1�,w>��2Ms�K�M/�ye1��O�b<�8o��򺇡�wBp@-�\*�2��r�K�bZ�s3g'|��X�Ǿ�^��z�SWj�h�W�0�e�6����=Oϸ�]���um�6cu)��)���+}��Y#@}�/\�����G��u(���E��2g�'0��??S$���0Q�c�A��I*�&(��$���Lg�`'^(��`pʹ�b��HI����뗴t��s�GTC��b��ആm�]��Ϗl���d�� ��d�L�q+���3��L�/d�P��d��� ���3*�)5��~�FY���;1��/VN�\�F6�չ���0�`�P]x:J�Ö�ˍ��˥�|�H:�!
�Cn.4����U��ر����|��#�Q�e���th�߇��;���ς�$.^��L��׍�Ԍ�Peľ��X���.������ˠ�f�R#�;�����F�m�H�(�wU_*�����aC�Iil�J�0i�[:ڲ�qL�xW�9��y��8�@M�0q��'A�׾�R�u��v^�z"��<��ź�aF�e�WO�j���Jj���' �+���W(�:۹�d� ���w��˻��ޅ�� F���SSG�]��.1��7UЫ3FS�7����?��?��4J��R�ҕ�#�e)-Q˜��y���FҍS{D��hL;u��R$���W��S����+a����P�dxwy��礪�F;Db��=l������Q���dj��+�iW�RgU+}dbG+&�Ev?��.F!�޵�>�@���[�r��Ht�$-� �u�����)d��
䘇_���{�t1GhF"�Aa�wO�RA�`RE``,e����<[�������@�H��Y�$}�
�,��6
C�D˥�Т~���>��Q�����PB�DH�w�����h:`���p5�Xb�/�!f��^����J��fl�b�G�e� �,��	��c�X�4��� ���^�P�����<�`3p����>7����Cq�C�	�xrnF�'%�^��~�W	UZX����Y'Wm+j!@��DI�:�������T2?�!��3+�~����F�k��ȕ�!�k�ӀX��Y���E��m�z��;��(a����n�:��ǒ?�|4���+g�[GW�M�!Ø>gg�v : �����'��ge:,T��+��D��#=���aĬ7���P�@`w�@Pw=�s��&	WGꝇ��G���#c��=nI�t^�^��Y�td&jq�w�E)~H���;<��=��<x��������AQg�\F��'l"_dh&�.��P�o���g��&�$�	�N������W~��0���;��d58�w�
a4:ў�$�0�����W0@H)��p�f;>�FP�
>К�Q%�z&q��9(�K�eܳIvX���c��7l��7�G����<����{?W�x�>
M;(q��sq.������B�%�1�\iV��4O'կ��&��Gh#2�lj�9#��֚4z�{I��am�87���v>���7�E���n+��O�K�X�Ď��L7&Gu:���~��%e&P���i՗!j~��u;}�*��$)�	�x�)���ch���v��j����3���q�ᢐ���>�鸵E��Gd�_���\��2��)���^��0�C�x��R�7:e�k)o�4��/h$K
0���y�Td%P{G�:^"�]��䈕�>�o�q5^
�\1��f ��&0��ad���i�������m�F�P"��Y����g3�ȣ�k�O1��_ܹ�W��������Q����з�w�����re�&�l�I����@d˩�����x�/��j���9j���ƟO8f�}�3*�ٔ]��*���.�D8�7� C�~�\���]��<������%�Yf76��6�)c��N������;T�ps�s�zڀ�n��� Q�Z#��I'��7�+ɫy8�52�sGv��/�tqꆱ����(Lua1���-�B�ۖl������ƺ13��Aْ��ǆ���-�����E�`Uc�J�����^G�����8�q�z��s�X�l@�ns��ف�1�9;�1N��F��`���<�Q�ܑ�׹
q�I�Rs�u3��� �l�F��l����8�lr�\��"4״����M�����!��9����m�' 3��H�,�Ԯ�Z4%S0}��B*���52�JɃ� d��^7ܑ�u������7\�u!M�w�.�_��l8<���h�'X9JqW�NB��tiR(�( 5��D�
�F�xa}j��{�3�#�G��kJ�����|V%��V�E�UP8�Нf�(�/�^��Z�r/>���#�k��A��h1���f�;~�4�B%E���w[���q��<�ٕ����D�� ��a���v��?#3�3y���˛��"���pK�I���.Ǯ��F�ˌ'�x���X�cH�b+a�~��Vgߑ�	�����K?")B�#.+:2���mgE�9F]������u���S[,Lk�xU5Yv�3Bh\V�w�`�[�y�	��5��$��	�A���ċ�r�9���+ቧ��YWGV��jQd	S�5d�K��rV��La�j,�E��Xа��ԆU��*7�d�`dj I����*I"��媇�h��	R
��Ԝ��0���i��D3� >��c �v-�u�V0	�p]�{3�&M�;�6.���ή����#�B��A�wu���j� 7D֜*�.�YU��7Z�2�V��n�
�3�)���d ��L#�y��^�:���8���{k��#f��Q�ρx��U%��Fl���Lc<n$�Y`��?=�#����iR�Za���_\��Hg�����h�D�J���呭|sjf��~�0�Xt��b�0� �/%�<�Q�緑#�`�B��㲦@yp�I�N�<�"�$�W����p����Xs����)�jT������Exyf�Ǵ`R����ݤl�]ZP8И��xo��DM���K��,Jd�l(�k��3:f�R�������c'lIF�Y�ذ۫�3y塕X�(�k�%H���̒��Zt����U���ĦhXͽ�6wc"�B3��z�0��po?�F1��Q�U���GƟ��?��ޛ�Ȫ2\�E�O�� >1���P�]4��_��at=��`9�.��YBx�Р�>=�]AV3f�r����I~VԼ��1%�_+!�[�ܒ�D3?�!�G��z�.%0��\D]��צ�'��֦Hp[�|�	\Ng��/� %��*���S���$�|��;�:k��,���\�.�H4S��ӥ���>d��Zl�ˈ/#q�Fu��~0bӁ�C�������)K�K���{��
�Γ�M�^�:�d�^	�*M�oG�Q��)ݤ�@S����S��EB}��H��ے���;�A�R�n��!z����p� Fc��3BQ�$���V��vթ�S��
��CΎV��P�]���=R@K�P�m���%"&���Ҽ�~�C�WR���3ew�^a�&���l�:�K��ڛ��'H�>�иg�Y��=ӵ�'��\}�'�t�l&�f^�X���.x;7�S2��l�d\&U�P::�D_=a"$�wf�V@MZ�?���p��}GA���"^�����7�iAR��#K�[�兿	�5�^$(3F�9����"�cB�8��h�ʎ�f�)�! ���,�fg��1��=l�
^�p8{Jo٢�.3�q:2��Q�PNX_�3��6�Z�ͪux5�8m$�CX�H�tubY(��U����Y-\k�m�ڱ�b,+��"9�Nis�G��LG���W��$��0RG�=G�du������m��cF/lu�W.����a?�~�{�f�aW�|�m�F��q�a�S0`�)UcK�U�V_I�$��EU�ݱ�g(��P#V�b���3�i���VrW{	���'m�wYQ(._i:yQ�� 	�➋�|�Og�j�����L��Y<�<B�ns�̉&Y*�n���X�	"0��լ�Z�S_�<���Gj7c(����n8�x$rO(N���M�<�Q�G�v��;�
��e
M��|� ,'�x���^���a�7�זʍ��f�(���#���]�t��K^�N�ǲ:
���ǎ�D���L����t�Dl�2�Di���9w�0x��=���*	��FV�{Y��P��(�sv�0�E?�,�fY0M-���YZ�/�i+*�"(X��h��AEM\�"M@�H!��\>�n3貳�um�lȺ]f�f�EE�/t�)��ț\�/Z��TV���4�&U/	w[*}b�-qT�F�����"&�H�Z���&]AX�5E8����z���8��y������
�s~?b�I�uO��G�tA�.��r�Lڽ��"��0v�{"s캱Ʈ���F�x5�&6����sue��
��B������KV���/0�>`xcU���h__��)�|�:X���H�8���c�e[B�9�k^���7V�����f����{�Gaek,W����ĩ��}�%�0��#��;��G�{�
����"x�J[>��G{�'�u����y�PlQ&����"���Ş�y����{�vJJxmؾ��}�ԅ��z�W0/�K�Bta4cP� dtv�)ض�����w8����,�����E-�Un9G�u��M�s

F��}5`tE.�i��h���J�ah��/Nn��&s�S��q�X��	c�0q��r�&8��͂�T?��a.���n��l���3�y{YGV���`����8`�[�:��)��J_xr�s�v!_�Zu|����$���y^�<�ä�ۡ��3H���h��Ѽ��E�!�?�c(��@��K  ��\��۱贼�BՕY��	�$4&+ǥ�&`����J�=�Ju��sIlP�,�R�Ҟ3���{�����<S��J�j�Rn����C�����;���7�C�wc쫆����P�����4y��M��T��X�l��3<C��\���ۑޙ�U�qx��Sř4!�s���Q+.��M:u%!��2j=ҫ�5���ddcS�YF9���� f�����Ց���L:�L��%�~U�i��>cr��%����V�l�u�J�E
�[8��[%��A=�M�dW>����������K4�S�F� S��R��F��eWSg�J|�t��/�`��9�Ƴ�r�UoT4y~{ ����ﲞ���������X��{����$�WU��qI{�921���,��UP�Ӵ#h�hzc�|)��F�?�@jvX�ƚ�I8�d�Eӝ'-�`|�+��;��@���D��&(��x��]�
P] ��s�5�L4���w,�s#Q���ck��&�8�{+N��OU�da�B���Iq���u�׀���цl	�S��n�kN:6^7�LE�T��CL
27.d�44��7&���S�;�|�tطd��U�e�?iN�PaVO�52S7}�չ��;8")a5��E_p�a��d�P��u��k;�ț10��H�6	�Q���фx%�\�W��s�1�W��.}n� _�P��uq����:7룑�]j�=��`<�h-Rݰ��N��H�D��h�M3�e�k�y<p�ɲ�cY=��e�APc/�sO��ĥ>�ju&�p�32I�c���xo�V&��R��V�gM�@����� Rq�P���J��Ł���)7̒*n�{y�m��@x��Bbݴ�O
(�&�_�moOx���ܜ\�&�㾼!F�"P��mD,���Ie������zG��On�� ��fal�ׁ
?�D�}]�Ul�eS~�[x7ȗ�ђ��<�L�}��=m�+I��x�&��2���dZX�J$��~hQug�,�3�C�S�ٿ�j�H(�l�>D*��#��Q����ѩ7�E����yp�tD���X��>O�B⿂����k�m�:������q�u�w��E�eZ�����/c�g���V6��LFw��d(M�
C옷ӌ�r���}\ҥ$�6w}EZ�eiT�?��S��`dz�.�}�I�<ɗi��tֶb��M�eW�}�����V��_��S��i��;ɜ@�=��HN%��@��t@xz�Jm|w���9qw���ht�)��+�+�D��X�$�/ó�6���i �*?崎���P�
o�R������֑p�g+���ۙ�� ���hީ
�e<�$/[?�t/�Wy{G�2�C���Bf�"�+W�`&i!���{NpwG�z�^�t�Q��$�#����a���h��H�kUs���?b�4�W��TN����3YN�пY�^&n*�Ċ9ϼ�&��:<}lS�pƀ�5���N�V{��S���k�M�gXǡ��t�?����@V;�'RE�֑�a!�'�FJ
e���!^�L���bw,�al�m�:ـ�&�ť/3<��ڔ���#����{�t�?S,�k-��|�P�����VG�Ƒ��`�:ͩP)q@����� �9U�?Ql�����y�\Bjb�e�}�"�A�+���j�\M@����.��?�h1ҏ�v�F򕁞���F����#�� v ���v ���i4��\~�N����ۊ/���F:h���Gxa|�l�4�^��3M����Z��f��	߈ V�Rt���t@�q��;k8+�i *����4���q#|A��ҟ?���K�_r��~M�]&g���Y���5�e͌���I�D��K9�˓�r��E-�<��g�f[M����}d��|ã�	���m�ڀTcLi���-�����4�M�#�軐񀃾��;4#Tk���S@ �~�<u�۝c"�`�ٻ��rU�J��/"F\E�s�f��,�"�5;����l&A�G-��3UfC��G��^
L��.� '���H���lWTaʶR�Ĩx2>>F�i���jBE�4�-�E�
�%*���P����x�b#FN��2�`�
=& V�����G� �S�Av|}��e��KV��M�?�+v�q�������[�����O6܆l��?/�l*�i�J��e+D����˕m��y��"��
\���)�i ��go7b/r;+�R�O���B{��aX�8��l�|�_{\��^M����X����gXQ�������ur��w�g#R�
����Ӣ7�m���bM�B�7�+]5�l�mK���#�H�fD��i2{�H!�n�}}�g�[���ţ�Q�RapOYK]���;$���m��A������-�'�Dp�3����S�t�����0:lJ���\6�jK�6�Ůi.NW��j%�&��G�w5��!c�~����V+�8��;�圌�|�E���,+
��O7Ӿ�7Մ�Y�e���O����{䘺��f�����lks�څJ�@q��.�����]�)ŽHqww����Kq	��˺ﵟw��}<�\c�y�s�ɑ�qW4^|B��`ǭ�.*%]_o�ړ�㼘��]�@�k$��R	gY�6���<�`�:
�o��u����a�'�Y��>�R��rډ��;2	���
��k{RV��2Ĉ�P��ȕ��]�s�I�'yK�du�tUo�Q
��ri/K�M���
NX��5I���L�I��s&��p{~����w�.IB�/:��K>��X,�JK,p�6�#�70���+})�70��Z��dR�4b��qA(!u�&��O4�B'F��'��L��u�e|~[��9�l(���3?v��O�CkZ��._[U�/��Q��ǖPH��kѨcs8rG]�{=L��҃�;tխK8��l+��JW�q�Xj�m�M'|�W3BG4~qG�=C�i/���r�.���M#��!������F�����ˎ	��N\	�]M2�e2s󷾪Oz��2���c���1�F�ܳ6�&a��3��E�������TU꿳}�h+YA��ؑ�mr�7�.E�����N�iz�q��%*cT(��6��1Z&�lм|��R�TP��@f4��{�[��'�(������m��W���|h��(��Zٳtɷs�ԣ'o��V�# �S�Zn��P��b�}��C�W���8���97���(��	^�a@���#��E�R.i�w]ZS�S��6vxhԅ�鿞�܉���Ի�3���D> >�~�<��"$��,��@�X�6
���u��`I�g��SjE/�&u� 5����m��<�x���d�F�@��s�����zzj��z�X}ch��Hg�kʑ�h��[s��ν�c������/P+͸v8���V�\ݗ�ĊA]8MS�~'��K�,	
oY�P[��-��ϝ��!�h��dy�F�r��������N���N�)�R����SR�����W0I|E
�c^@���e�f��E���$�6�Sn˂
�*J퀣o�@e��y�"p��������ox���V�|�
n��[��8Q;�ZEa[ð�=��Jq@J,� �-�D�b	����^�ZjD쏳:C*�%l���{�2;���B�����jǶ�rm
��ɝvi�
[�O�UH����46쬅�A�|�E����ҫ�Ԇ���*�YU
&3�.��gSx���<����f��.]�i�Z�"HV��*�
���eӨ�D�p��Sf�Ҟ��<jGb��	ۈ���va5�Ek9�󯱩�o��*��7K��{ �$7Z���L��V���T=�ER^��x}cp�& Z��'�H��R͒/G�����E��p-Z��K�L#ĺ1���I�CN������b3V���<�u����Jf��MZ���i�I29��l��ڳ6j�/4� IB��8E���p9#�Z.�p���$�fĸN��w|�i�c���@V�Z��M�FY���^�:���/\�h�A��x�h�+�q+6�U��-�M�l_< �������z�|�M��j�u'��{$uiU�q��3v	��Z�&Q�_,ux���V�tc��hf,'�_`3o�Sfg�*e��
b����<k�$�ʎ0��	�Ah6h�E�J�K!�p�.��2)��eAQw�*�����spm�s��Km���x �qL�Ȉ@��Wy�(?���͡���1���QL��?1��B�e�^��'pԁ��u�Rpv0����X�e�֍�ue&��W������3
O�@:��%��TG譎|N(աu<d��a���4h#E���R���
�U���%�<FX�8|�s�HSW����ʨ'��u	�{�t�����cx��6�S�����x��ß����nB��Ӊ��|��n�V�j����eǃ��7�����?�#�R��4<�x�r��������Md)LNt��Oψ:�O�+awx�̐8L��%���c5K���&i�u�=��v�D)�᳏�M����J8� 4Wqqd������u���Yd\�{��<#M!��=��X����'����)v�C��pY6�}i�W^)h��S�v�L"�6�gƻ�R��qh�m ޜ��)�ù@�����+�t,�}�Xiz�TI�����dQ�u�]G:��[����O��#������X.G�q��*RǶ޴�f:G�_��~>�V{~� �/��!��\�L�e���{9t}�h 2c1��B���� w}���ԉ�T�m�@!k�*tR9�>��aI/�U�6��	�'i��?�ԟr�a�B�5_���"��z�y�>R�a(E�tR4`{�j^!�沄���ߣ#W�%�v7�{0���u�IW�>����T��R|ơFZ��O���m(t�<���=��'��m	�x�1����Fp/�[�u��hLk��%1iIe�Ӥ�����6�2��@|���@����$�~g�SϜΆq�������~z��R>���SR{�u�X ���*d(V�!;Lo�3PȐ��e�M����o]E	����@ܙ���-V1ضؾ��d7�G߻��|�?y{�ء.���t���׎o~,�;��EO�8�[6r_]�"̩�!���q}x���:���u�\�ɼ^+f��_�u��0�j��e�*k���/;u9f�&|#���^%K�F�˙;�ž jbW~��>Frl�8�l���xქ�o�1��-�RZ��_�x���B��gXBG�;��v���_�.qT�$���2�����6�nSa�$v�g|^w(�����:<���)R���áW�R9�.9�]�-�^�~�9�����ɟ���9b��Ŗm0]�M�m *Y��uw�-q_���A?m�G�Q��hI�����J9�j���뵌��$�W�2���-�z�����	/8��|��<��J.3���|�Zx�F���d
7;>܇a�k�=�(*��0�樥xg��뮞mMއ�g<��>��T���t�AtSə/�Ks�O�Q��>Ym�3؆2L�C��TU]w�Ed2ggra'*��w]�}2��Ф$g����1D�$C�{�59�j�t�O�O[v\���-g`��>z��V<�4�!�}g��U��cD\�	<����IC���d+���u��=[����R�k����"W�O�<���^J�g|��Τ��?�9�#�Ow�ڃ��4A�f��λu=s�1W�a̠)*F��SR�����ω�	N&�$燔�^����{�����Q���G�Ʃ�q�_���g�����2�^�J�<3���Y�gئ�U�|�w��Rg*.�q'����`����7���H7I��5�&��ou9'�8�c^�L���}�n�����B�������a;��/���NVk&�W�f��?-�͈�"�9�� �����]������抉R�^n���+��LA2ѩ���|hߟ���S���y|�f,2��%1��W��#�Yf��7R.$R�����>d�:$9r,&_	�|J{�Þ���y|�떕� ҉O�uO֓e}3���X��rh�e����B��'Ә\�=ۍ���|��o�s۫��h��tw�� �����'�
BV0�z��^�z1%>����k?�hr+59vI�#B:;a�g��q@:! �3�Uw�a�N����N��K��`��u���|H�������r�W=o�V���Sk�����]�꟡M�@ꉘ(��\	"�����"��m������X}�*Q��������B4�E�Y��hvh@�lXt���<��( �����S�k� n���l���O�c�p\���U�B��X�b�iGpV�<�ݍJ�d!&HF��&��+GF����p����A��5��47�q��8~8Ѣy��s�,�ؙ�����n�7,���rN�1a���{B�<�H��e�����J�c�ͪ�0C��66�U���OHjQ�gZ@�����ZxB':�6���?���e��>ҵ[�%���R��u��f�^Q�wK�xw���M���USޞ�t%�$��ģ�4%Icbk�0��O����Y3=8��Ӄ|��}N+��@���z�]����|����zH�K�+�~�/�x�	��7,��7:�0��5{��7�ӣ��ķ~�������� b��;MF�	x]m��S��ȶ�����i�%_��P:�5��鬡Y�,�f�rҢr��>�fP1l10�=ӛ&��&E���t�V�d8�<9�8ݛ0�j^����Wr�H�w]Y���}�l�ְ�q�����<�r��y:�s����wxҊD�$5�dg����Kf\�>-"��{�H9�ެ�:�w
�}�:��~b��
*���-��?�B����ϝg�g:���	��Kd�O=�M����o�$���B.��k ��zy�_1C'�,�ei�M_�D*�����K1$h%^i� �vE v�bʠ}��䵲9S�+K��)>��D��kG-KZ,�ũ�(�����9b�;۠#����d�>g�D��~���9�����<Nz�%�|����as~!�ȠyX�_�zJ�Ǫ�5@�v>gc[T�ֿE�3�<�`�[.f��� B�9*��A�o�(鬒�%���&Օq�5�x"0h����`��PjVNb�F�%�������8Ӧ/�������3��{�UmMn�'Gg�퉾Z�!�W���^1)jD2Gԋi��=O�,�p`�L���4GP��	D�F�&�+X/1Lif�w�Q������N4�W㏷�`��m���u��4Lzc
�ϸ���_"���"K�D_�rbPd��z5�GL/:�S�����8**�.A�76��i�p[7��EE�PT�"�] ����k/Y6um�E�ʲ<�q2��]�IL=y��H����L��SY����	�y���{
O^��жj�}���GDIn¬�4$1��x�!��Y}:�Z�J�4�*5�����p��x|9������1����m�j�6�^w�ـ�_(I��Kx��}*`��Ӫ�p�1�0����-Qnj���އ�G!��֕a�K�aԥCgVB����W����L|W/M��+�+�S���x�+5�����:�3��)E�d��� ���%B��Ujv�����b�bg�[��&��W]"_����UH�;E�k�Q�AP�e��T26���)L+��Q4v��'��w=f�ĕ�_y$py��$��*h�A.���q�ZS2��tι�I;v<�!*�&�[�K����w��cb:kh/��(pu�Ԓ+Fl�#t��r8{�^l��Q��R����7Id�(B�z�-�h;����7-9v\p�@��C��@X'!�~�-�E��#����u��	!�l�q?�4$�GG��g���]Rb�q��۳r�<Zb&h����X&��?qpp���C��q����/&4��VF��qw�|��%���ʎ�������#$��}U�@x㾟��A;���ڡ/7�4mze@�T�I���v,^h��;$�2{̆�WzB�mZ�Ky��A���}Vƿ��S|sH��'����Ǳ��D���=�ޑ0���a[��o��g����Ft{r�#���*��C����QZ��rh׉l	�Xdq�c��zB��؟�>)�D7��&�����4�ޱv��ꦮ�����j�E6d��2�gI��Y��KK~v�my"�֡Tæ������¨��eg��E}r�M� �CgD�lzC�|�xE��"q�I92蕙�ٌ
0ʮ�r��G��w�k�:�/5���Z�o��:���\�t?���z,7٧G���ța�;$Ӓa�z8meF������#9�&	����|K%����\�dhľ/�����%a�J��0�B+P�T�rY�U�U�K�xs z�~�i��PkbB�7�GN-5�r� s�~���$QV�Ѳ���Ԕ\6��fF0Y/jW��lBQ��q�PE�>�ڄ�Q�,c��ӟ��):�H?v'y��N���>c��J�ּbz� �2���z��D�>����(���Ӽ���ў�k?��-�.|NޡT;��>�R�c�O>;;+��M� �0�s:�.����D���K�=�<�ut]�#�:����O����){7!��r&ā=�_�u�O+��ZA�47���)���D��`�N&��V��SLA�F�!�&[�b��"_%��īI�r!!�Z<�+S��:e�Ҙ�D�z���Y,Nu�=�@��T���tz�H�H0�l�G�о_�m򦼷�Z���'���uCd�/>���%G�(Y��h��{�Kԍ�§��t�z�����3l���c��N�&����㬸�{����?/��z:JV�:�4��;z�3thu����E`^/M�i�b/n���K�[�-�S���֙��.����M=�9���6��F2��	�=Lؒg>��t\��\u���S��LJSe��3��E�'�㯶�D������W23fe뵃��u��[w#Y��]�C�Rwp�S�(`��AHԳgJ7��-�[�M՚��Ba2A��:�m�M�$�5���s���[�j��|�����.�Ol���e�h��YVL)��v���rJ	�DU����}��]+��W�9�����-]>�U��67d�ɧ���%*����}_b}j~��E�x��62z������mA�O�_'fK�P����V��?8�&y�*K�� O�:s^�,��)��cP��[�t�4<):�ԫ�P|D]R�M��=����n<�K>N�ĉ"+�����Jk���{����]l��!}�mdU� �|/eY��ɋ�?�t-�u��Ǳ����̦��ɖ�(�9r�A?�'��<�1�!F���3�<�v�����|HkF�:-˘d�NI��1�q
�'�/$%E�y??;|bIqP-���_��D�OQKI�cU���>B��\��a�Y�`.�u��n�%t�0��=�1�Yo�15���$�.���noVr��x`�l�O�׏�D\�a���� �RF�T�������~��K���×#�7��~�{峖yT^}��~6_��˩��y�������q(������\��A~l�������������kpNZ#q*3v9Q��ˠk۾!�@[>'J$��_�A�k���S+�4�$�T�'�Q�b����n�^U�XE��qF�>���~,�oSI`'j�J��]z ������c?�L4Zt'.+j����4�d+��������!��|RGhH�wh��#m�M�����O���2E�8�A�h���a� ]�-�ɰj%~#�Cs�i��o31��
p���T��G�G:���h�|=��7 ����8  A�r 9GA됾�n�w}=���
&$�a��85�'fJ{j�o��t�=��Z�ֿ&L�oQ���1�Mc�����`5�R���k|�1�%��Y��]��R��h��,���΄����ÄG1���[�ƵkX�k�SM?����y�Q���T�3����2O�%ޝ,���:�n�ExJ�E���MРZHDuY~U\�/u��Up<�˔,�۠�~"�~�*�蹄�x;�Bt��a�_�y�
_/by����t�y�<oa�c�u����lL�@t7ڔ\�����hL�l�
OV�m��%�J��5*��."��ɶ��|6)�<?�/7H��ƙ`�����`>���>������:���e�tbx���O@|
G���;��M�d�����/�Ogp}��V:qP@wL���|t멦x��C�=?�$:����8�Y����w��W��f�1B�.<�M�pޮ�l�;��F-�%.��<��3��cx�ʼ������7�*��s�9��.����-�T��헑-�o���m#�Ns�2C�s�����@E����k��(�,��t�mxVݲ� N�����e�Gd����0���⎷C���X���È�B�;3�L���ǃ�����
ʑ�.�R~d�����r��)�b?)���;.Z�m` ����گt�Â'���2��~��������~�W4�!��~7�SGs�s[��.��4ٯ���r7[$��(��N_�V�~ة� N"���<��I&�zh䔭~��X���Y:A	��۬Ԟ.���F&��>�$9����\�o�� �}�,�i�Lp�gdW�4��s��m��g��V�IM�G�||\�_+sN�zD�$�G8��ω��,U�O�B
����H��<*j���؄��L���4���Qy��F �����)��	�?�rv]D�ư�����
�J6c�����=��ѱ���|G�}8e7b�&G5X�Ac��"���8U�I�<�~ޡ�>���7�	Co]���2v^�<�B����F�1\�+�m�r����Ji=P�sbΆX�~	��پ�K��oď����
�?H�����l��'��ݳ<�z��O��D�ɫ���m/�;�&��Eq�	s>��8	�V�S��6�QZچ��0Sޫ=�cZ��݊�W�۾|j�� ���iB��J���IGF�K)r��Ȁ?�a&PÎ�'�n�1�>�{��y8��1|[���9
�I�^fS��d$t>��s��ݕ#�QJB6t�F ^�β�gRn'��fT.}�֐I\!n��Qx��/�N�<��1xg*�*��v;�#M����^�ܵR'#���q|���p�����Xt"�#��R��"o��yqW�t*G�j
�iI&� ���؄L�U�ڞ5]�^�����=����Ӿ�v˶��iЭ}���&�ʓf�՝�[�軜��n��*�?���c�!P|���h+���!�6"C�I�!��{�5�m��������h��@	��g���ݺ�.���0�n� �̡�G�N~��ӀؒH�`�`�7 8y�Y�7�𻡽���C+P�Ӱq涡��������;��O_��Q?��m�n$��[������O��ɬ���Z��H��A0�� ��0-�l�ʬF(�S�o3}@�á��c)v�_���t�	t:&_�����/��գ�=̷�t؈�RZt�uy���_��n�*@U����_-U�Y�O";Q�������Y��#|/�ښ������T���<�����a#�K�����Oڋ����M�	Z��0��{�o �Ǩ�Z�:�߈����Մ�[�{Q Ո�p�j^>�z�4$�t�,"�������F%�i���-���QZ�Dڵ����o�Cod�̮�.�ݨ~XC;�ȴ4�2���.V�'��?~E�m삊=���[�._������#��M�9�#6^o���\��Va�` \5ǚ�d��A���1)�ۂy����a'!*�;��m��FG&�5�j؞�ʩX$OY�J��W����1f�%8?/���aM�]_�t��5KPk��u��J�yJ�yƕ�eg�NW+I_�t�'������h�s�=���'�:���Fd�8���s���|L�!���g=��=���!m�Նo��]W����?<�n�@�i����Ny8��R'߳OX9F��T�+ uܢ�Ū�וu�c�cF�vW�e�H���AW��r[����#�bȤ�W�KUĹtZ0�,&9j�I-�f��A0��ߏYW�zn�4�v�P� ![�e���TԑB�BS�wEx���d�{{��zk��'�����y�"������)a���h���y��L1K�q���YW�N_ٴ���'h9T�Z��AB�p�a�
�4����a�	��4�%0Kl�mY��,F�afJT�[�}6��hlT����1Zp����"Vb��&���x��]�L�-_UL�R�$^0�>���/�zl$\QN��4���vlH��v`!JP���ĸОX
 ��p>De�d�,ﯷX����t�_��Xwc�Q��p�>c�sź$�{����d�b����ϯg��޷��;vZ.v� V(:x^����#���;��$+pc��c��k���!�!�TI�0��{�4;n�BѦ��[�!�֖��-^p�F�qW)f��L������k}#K��Y�:|b�W��?�� �K-U�%��`_̕%����1xv�L����b6����$�����2g.�dw�|:v�n:o���d<�@V� ����l�S!�����K|ѥ:�%��J�x-z��#FCZzFLZ�ݔRg�˙����9҈L`RD��u���H���&��A��z�p0�a���YqM]�\�L�Y��`�1�ocw۩dqI:�e���gn�z���nR�k1-T��ixf�e$�FV#@�I�0� ���E�ݳ�N�3�"s��3�E�^���������? W����Pӌ75�x�	�"Xo���4��x[`z����L)�;��_�s8�fzܫ�I�.W��ZZ��v���7|�	 � �7�,�Z��\�<�X� B�Шv,v�cҟu�G����9����&.^�>G:�pJa����M$!#0[�/�Jc����[
� h��҃���,���8U� Xɒuo������_d��JJ7��p�p���e�tː&$>���Z	BT�t�f�*�p�m��������X���IG5�����:ڰ#��J�6 N>�����r����@��w�nᄑ r|߱fr����9A�	�u>�� �����P�ix��(V��5d��ui����S��xߚ��ybN\�<�K*>�E^��]A��F�-0��J�]��QL����wZ�ua�0���qۼ�p��QB�8>C8}��
��N�w����#��G�Krą`te���]��
 p�f� Ё�������/2,  �}{`�S(4@(2 ��H+�=W����~'��m1&� _z�Y*RE���+��lN�����kC�!L8-�?�6~"�L���k����@8�r���(��?��|J���lz�?Q�Փj���&pJi*�&4��<�+F��&Ꮇ\��.zՙ�U!�g�O�^u���)��l��V�ߌu默�7T�����I_�p�$L7�1�X�c���������xe1�#�
�����fv�������A�s�5mr����u$Y}��ߓ�^�=_)w��xc�!OG^s���?s/	{�:AW;	��ԣ)��R��g��DE�K�&�:e������k;'_cE�ֺ�BK�n+��(��S5���8|�d�錢"X��yw�	���[!#!�*�����a4��oO�Wq�X�l7'^���o��(b*�%��أ����ڦ��Qr����w.��u��6��ԯ�#VN��G�S�I[���A�[�M�8�g�~�O��g���q��),���Z����JE�T�$#�a5���.r���U{�]J��!B�հ�8}{#�p�,>:S�����������$���;*G	h���r�Wi��b�tH�b�D��^���F�=���4*�v���!~p���A��.HH���%�5�|Qi���Yq�Xb��f�f?�����B(�ưW��\ ����[஛7߉Bp�:���C}�
C�=�e|��Z܇��cC���)a
vbr0s���h�0�=�AIX�����֜UV|�n���ζ��פ�3�蝩���N�/k���&���.��z�ⴟ�͸g�=1p�\�����IrD�1��Բ���Mb�鶿��ۤ=�%��l���Z'���{
��zv�J7��gC��ʱ��_���-�v�j'r��f�;l��W&67=y�~Wψ[�&��vb�Ah��^n�,����E-�/e$e�&�(��a�]�T[(���XƠ�6�|��B��AH��%��[�U��V?��Z�1S�y��%F0�`54�xnZ62����XU�T�\R��9�[U!�X�� f��������8W5���|���l��l���]eke����Z�XE�:�F��V,;��B~�V��x�DK�7�7C�;� �J�G9����K��6�[H:o�G �3�8����礨R��X�z�M�ʑ��� ۑFz�����%J6�{W��J��3�H̦�q�,r��F�Jiu-�t����iu��M��3�r�j<��ol�O���2d2�n�n��6	��&̍��/�FͲ^{.mn��";$��1�:�����{��{����^�d�߬���ۈ��(8Q����حw��Y�g���{b���c�H�3kW�V}�m�\u�g���6K;�Y���7��M
 �ZF�^1����xv������nl/#]?�������0Б�n�Ѯ������,���]�7������i��df�N�)��a�-�Q�X�����zf��������\q�ߣ�{
1�= Ƒ��Gad1J�Uq�:Z�"U�X��Si7�����j��9������4,�L����^�D�N-2�>��^]i�Oi��YN�`\�^,��:�Н>"��2���d?���b������0;TD��>z�q��6'��J�/%�Eh���A	�<v�	���	�V�|$Z�Z������oB ����.�Yxy	��YZqq�\]$�tiN��aC�ytٮ��w4��¨oDY [ST)�����gM�(񰐩���#���VJ��GZf�&�pu	��{�0K�8@���5
jJ5ۉ����Afx�uݸ�)d�42.�ﷴD%o�Yd�&�("�e��(+��)��0C*Ea`�;�ƨ�Fؼס�2�%�<R��Ns>���!����s.����="H���ʱ�K)Ɠ;7�E��&L2s i�K�O��ɠwm@�b�*�����24���Bq���B!��;�'�%4��Y�ZLknȚ�	��D�}�x�)�(DsTu�>R��� ���p�a�L��Z�&X�p�#�TR�)D�WM'�
U���"TU���7m����͚pP�?|��}6�H0f���Kv�獇0�ٷ�l�i��1R�T��Q��#�c��������0VC�s:�/4c�f+�mH��V��m�Ƣe[%#�v��(���=��9��J��ʬC�8�+x�k����q�m��������Bqr��(�@��Z'?h�0u}8îXmP=39�3��e�x�I�����d8�������z����O�\Њ�?�#�L0ɯ��A�! ��H�C�Yl�l����aB��r�짩�"	����s5Z�w�1�e�9,H<��=��1�S��D �L�`P�Y-(��;<����pi�1��|���W�}��d�����e=���cK���ǅ��<������n��f����ʎڙ+�F�s.����t�n���'�sv����y]��"��Ϸ����~<�-�E�*�JbJ����3�� �������i�#~�v�,>�9�z��(gš]�Ql��8������t�x�W��J�i������B B��g�`��^�~�9��~;�%ʣQ-*!q�&��G����R�E�naw��]D���UHjW��ZE3$�E�{�?Q�����&��3���l�Z�)d��P�HO��w?��\O���`����a$˽O��Rh���C�Q�.%t�ۉf]UK�8��k&}],��6!G+�v��&r���-6��k��eJw	;�|�V�+s� �=�ө�e��a7\m�&R���)��d�d�i�v�0�5T���Š�n�y�Vk����T��_����YML����^2=��yn�A�*�W�w%a�g�oބo+����#ZV=�3�0Ȫ�3�Ĝ*��P9<Ì���2uUr�7a����KB#|�l�V!��My4(KY�{t+��]��	S�����f�Xc��>� ���H�V�E��ݥ	����Ţ���W���$�j�t�Q��X�I���a����e4♧a��2�F6�_��{.hK�Z���b
��e^�h&���z�+q���-Z��~�����Z�5�5A���J̃�n1� �_���i�9���B�cT��[�:�C����<������`��i�<G{�(��aK5ʋ��zA��Z�ڰ��CKl�`o��h�Z��3ՆQ�1�~�{Ǭ�'m�/�َ�Ɋ�U.j����4|}��g��~�x�aM27˲�p�A��J��Ns-����S�#0ن��o��+g��h���wI����$��ŝz�m�u����W���n��V
���$�[�?�{����87��7��&�W�����=��z p�ּ�*|�f0++�h�"Ȋ���j��VZ
1M��4tk������5onS��C���� tҘ� SK�i0�p���4)�Dɾ%���[p"�����kaa|��(Y�Ԝ�Q���-�j�t압QN6��=|�A��'��D��
��wk�L�rbS֡����P�wYѴ2]p�;%J�3��VO�ą��+�-b�
'3?�^OڭF�:^�
d��~����DK�r�t�IEV�֤Qt�n�'M6���Mfz���x��p +t���8�&F���$+�A�y��%��S��R�k`��#�`�q�o1�{V7�u�f,Gsd�R��U]:~��G�I���/?��ṷ�@�j��:�GRi=�����0~ڽ�Ju�#A~��+�S�H��ꅩ�XA�i���7��fw����Ln�?J����ձ�j�o����8�\�՘8,9�s�� yr�x=�&I&��<��@�,܉=I'P^���O��[qH�'S��JN�*�5���uQ�N�@��\ml;����}M[$�]K[�-��1��$�ݗ�CVb�BP|�E{�v}��vF�(��	���Ŀ�DH��Y��n���ik��~��c�F�G��ӆa������@B�1��n�.�q����:	`��N|*/�Jlec�W�|/�n������Wi�5�$�+z5L�<�9������|9}��a�D7�y��[7P���A*��u0�oz����i�{
���"�:�%Z_mؽ^��)P�r�{G(	��8{lHݯ:����:;����/��2�	��-���v;s?��r���^�@��$׿"���wư�O���3v6at���$X䖻�I��r�ܠ����VA��Łc�ID0����애�GT+��<�T(�-mv�dײ��C8�S,Ii�2e)Ԯ��vu��D��l�}gD�}�.�u�0�=S+9���i���D�jc�FoR7!QͤUC\b����3:��=(D���t�j_��u����$�'8�V�I#Ez�!�I��!E�^�j45r�$:��{.�֤�8:�V-����\T��*�t�F���T׌ec�+~��F�G@(���q('RJ&�`Y$a9�x�z3��̸��0��$@/B@5�f�&a���xb"DFvh�#8]wz�9�al�|���
��:_T35�|�l��x���˾���&8���I>�pt��.�2�ɗ}@u�
��ꑰ_;�x?����*�Db��Z�|�����W�=eL�Q�O���)���=ȄA�I;]�c������ռ����m�����/2<��.�p�,��ƟK�a���^̑�,d���K
Ha���;J��YGX�+L���O�񈈋���OP�'�>�~�'j��w�G_ky�ÐTG�^��jc'�:���7O���M�$J���'��$���6M�����W��X:�9�Y�V�n�f���>�#��'����lAkL�T�q3��9��;����H���yO͌��\K��+�1���V��9��W��w<�C|�h��&��+�~'[��)J*o2�k!�*��mK@y�M�F�Ԏ{�k|R&�8m�Z��bih�|EC���L��J�F�l_����������9�+�����W�{��y��1�@�?G�P�xm�\y `���lS���ݶ̫kgP�g�g�M�A�[Y����N7s,C��\Zk��]��ɒ�W�=ҫ��׮ɲ6�"��bШ����6���Z���[�����R�i� �΍�IG^�렲m�q��fvg��O�L�M�b]V�����>��MI����&=�֙R��
�׿�G�n�LJG�ھ�R1q�!���O�"S���)�_���j*��>?��s}��幝��%7@g��|�'Cv�b�Ł��w$�=k���ɳsł���6J@�A�*H�p*�̟rD�u�)Ԃ��ql�3g�aƆ,]��z��h�(���_��=�m�y�9���F�������a��*}!TTm��7�c����YF������a���c.�NW�O�B��G�7��c����^������v�	g�S�^u��r>u��)�s�;^=f�p͌����#ry�$��vx.7|��mR��x�%& �Lߓ �]�x��!$���aݸ|��RqE���x��ڀ��������a=��͏ܓ���a��X�T���s�Vw~���n%��p ���e4I�?�� 3�0  ` ��&	z`E� Y��Q�A��U�_��U�_��'�.ߠ�b�q9��E ��
bU"FA�PK   [��X��D>  ?>  /   images/b521c326-5f2a-4e46-b9c4-2671f5fb6bf2.png?>���PNG

   IHDR   d   �   (�-F   	pHYs  ��  �����   tEXtSoftware www.inkscape.org��<  =�IDATx��}x�u�?3��ŢW�;ER%QT�:-Q�r��{�{lŶ�����;Q���ʲ;J,ٲ��%J�D�)���lߙy�3�X� � Rrx���3;3���Ϲ�����6Y�H���K��W�৯� �� M�m[�/���%���q�?�o\W�eeAܳw �n��-�Ć�����߄������x�=�]�q�N�<,|�
�ǎ^ܱ��H���P���ڃ�T��>�����R���`wW#㺤.���_�i�}^U���룿oD����?Z�C}1lk���4>�6���˱q� ��B'.^P�Ｅ^��?f�}�(j�eM9n{�	[[G��˪q��R�b{݁SʲqaM>��H��6 a����m�l.JJ'W/*�W���gj�ֶ(���Q�0zQ��T:GS��LbOw����͈���{����rܷߺ�߹��!�:2��܃=�yZ���,Ë�a������\���X+�m
��7�"����>�'���a���c�o�`4��ҧ&��2�no.�y]5�ws=��a���](Т��>��>75���o���\��է���������a��"L��B �[F��&�z��De�$�f`���\|��E��CMH�l��YA�r}:��Z|���jB�俄+CB�y!tE�1�?߱BQ�uK
q��-YC�5�i�]�.�h�U�|����P+H�_����&�;�� ?A���J�z�
|��fv��t6�ޟ�ׄ�$?�����������|��||c�Ɵ�=�5����|h4qW�*���6�qmF	���G���/ .綍��W��	!��en��6�]y;p]�>���<]����S��ѵ�������DU� ����s02�C��g-|���p˹e�������g!l~a�p����$��;+;q�M�CqYZ������Q��ޥ�]}
��l�[VUa�5�nx��!�m�{��p������0ޟ�7\}��}£�����ۼ�/����й�7�&\}ӧQ>o!ښw!��_H���~]8���y	oY^����,�� v�|?��6�߬w�+O���T�bx�9�t�z�u���EFP��O0��
�_������`+�]����	̫Y�ζ(|�5�Gె�����꺕���� ���W���/nT���#��G|f۲B��@"y�u�W_�Ҋ:un��uX��,�ۊ&}|B��ZKs��z��#�d[��f�ڷ�!te"�5�i�XTQ�kެ�)(����Ê֍��_M�[��ҳ.BE�bu��Ek�x�
,}��Z��F1,�uK?��P���7aϞ���GԨ i��{��4+/� �c ����ވ�ͿV N	2`�X�&,Yv��P�"З,=˷6a��P��h k.܀��buݚ��������t��f1��Den4<4�|<��e�sK�MJ8"ajB}�n��&Yjʄ}�lg�	yV<C2W��	ʳ|���,[�/�t�5���J]�-}
p�Ȩ�?v��K�L��H��5!�%!b*� �[0֧���aZT�p��g�}�w�)���F2���&�	d�4&���G۴ �Z�q��'��W����hܻ;ۇ��Z(Tm�T,��Q/'�b�3w��7��Ϗ][6b[�Vc!*B:bb}JV�~���pɵ�����a�y���a�XoGGLl�Va��G�W�QQj�����҅��:4y>��H��X��=�̔pf>vo} ���q�,KK�t�#�Jl
���;�K�Gx�OD����y����i�}�ī�Y��� 
6�Vqdk�v�j<��[�%8��/z%�����)�K^��8�AA��2�%��,y`$ea$n���[/%�+q��Pd<�6�%7`��ÿ�X���d�ȽG���|$;Dw�w7(E����(��"�����&���k�Ϣעg�,<p"����ǖ��V�����}Q���`�Ǹ�^A��:�B<��]f�ym5޲���	���[î~�fbj>�_�,'�N��н��El=����w"f��OEW���y�R����M�g�Z4���[^B����Rע9Y��^=�?�_x����FF���o'W�$/��ɸ~��C��,��|�)|�YQ�w�c���w_�I�u¼)D� �b��-�1,H��#-b�/��n�}m�I�\e��
����S1-��b���w�+���؛�J~GL�[]�O]T����_��_�\�7E,�K�"GP����u���	�*���u���O����5x�X��P�Y'\��w,�Ϸ�� G�/�Y���_F�F��Tb*,}�uy�xy5n���]<���*|��P�f1Ɠ"�Đ���ը-��C�k��lӻq��A�JhWq�޾���bp������B1�I��s?|�B\/�m8�(+[�U���v1��"f1mn��o�P�va�4��u�ů 2����J) ��-E�x|uѢ����}Gā��֍G��7/ă�D���|4������GZ���m��lX��pRܱ�/�'���R������o߿D8t�O��hRN�m=��1d�C��>�����m6cT�r�b��Ou�5�h�i
��kg/~(�mȟ=2�F��P�`,%�u�~w���qyM9M���A��K���k�*/�Q�~�S�hPy��x]����hJ]IXʳ'G�	�}
!�A���^�����I��}���#quۏ�u���!E�v�u��I�>�%p3�����q�Kyݾ�(>p�a�����$�bB ��t�1-���e�Fz��!�y���`�PSf��߼�|C-���^�����Lѧ6�gO$��p��g��rC� ��>Ǯ#a��)���<���I8�"=��S�C++��.۟��Ag1�l�<|��u�'a1C�Oڦ��3mn����Z!TJI�	�Ol41����&k�i�7�"�27�sK�	�ØM��o&����/�;��9n
!I[Ǌ�!|��&�-��@���0O2C��M����芕�P��h6�q��;ѧ>����o
ꎃG�9���>�rs���4)�N� 	�\��W'ě�g�6�R�ki���k��I<�>��ӌ��ަ�(N�l��(,Y
� ���JA�S��?��]�M	��u`�у�f9V}�nV�b�(�K�c���O-��<�Z����Tr1��7���u��4�P?�s�1fF�4��V�P]~nB99j�9�"�D\�4�g�jB���p�h�|�BL_/�z?L1<�i�>�!31� �TH}ک^��Q����S>h2';'�?��L���RB�<3�^|6M!��-�G�w��<�'0�8Y]�|�DW�1Rם�&V����|�Zl�1�r�E�"�r��O�Y?��/�)��O>s�
rst�KnAϊ����969c^��]��(ׇ��a��\}�C��
!\n����H�}�twU.�&�\�^C;�<"@��F��"����tw�'sޱ�#N��g.9�f��@�f�����!������̜T݇���c"K��D�1n��y�5�$��i�N�Q;��=�S��^I�R(��Wˮ�4��J��u�=Iy�֗��M87E���644�Dr)#'cٵq�:��4�"���7d���K�:��2�! 9I�h�̈́�x�_���>+��r�ײD,������Y&S>W�O�Vݸ¿���*������9�"�%�){*���x�g@��Y��/��c��wc�]���H&x�;ߊ��K���� �^W��'k{q�]w�A��/++ŵ��>�9���5c'��p�9/R@%�n�0������s�0����AH�7.���?�H$� LĿ�������@_��=����J�Al��B���X]Bii	��[P�O O�*WK�di!P9��Dm���E\͛��d?a; ��,6�#�IB!8i�K��;��'Ї�s�g6<����E��]
��s�X*��v�8���\|��O�8h`0Ǔ[��x�I�\�
����^���$�`$U��@}�J���̿��yf��L��4���k����-7Ll|������h�r]<1RRf*�%C�`�I,��c��DLh��-�����iCi�����[<�қ1�v}����n��⊍ruOo_�o��$#z�D��'%��]V� b��!>)*�� Em� ���Y���1T�ּ1}�eSLL��1�}��]�cV�fFyY��5*V�Z��#��(��8,��!�J;P��t�ir�7�?	��.��".bӢ�5>)(�[�<7�坐C<��	A/X>��"�|�䖧2f�Ī�Y������2���C���˗�I5�e�I�,���>��#ibT�S6f�\�S��0��(�8��z��N��23m����K�8S�*�R�H�$(��d�>$������"�D��V�Àf�H����s�z�ODD�^�-P�)'l�G���R`pUy)"9�hL�)�ז5�ׇq�����P0�E�cǠ������&�p�,�nj*�8{b���ߜ�^�#� ���ڢj�n���◝�t	�Gr0��f)c~�@���}~3^���8f�����T\�zi�>�{�,+Kt�I�Q�������\�b�����񛿄����x0�=X�>�*�G�>�E!���Q��ڑ4�D))$�� ��ea|��w"�`������Ư��ʰo�L|O�?�����9C��@;�'����.�}Ǆ���b~]bb�����N&�J��ʠ[��!~���A�rJV��1���B�WU�$FOw�*�p�D��.'�ru�v~���G�1|��a�~d+�Ǭ,z�@��á*�~�|I����q�?�6���gPG�U�����)*).�֣�%3$�L�_���2�T�oSot!��B3�O�������Z�"ĺ�
9��
�D��c�L?%C���P��ʪą@��Y�ɢ�BS�_��d��sޜ���A�pL��1G��r����Ю��;�E(h�az�3�l�)�����$g ��j�V:Ru�<!2�/{c6�z��%���?��0D�O�~����$���4r�B�AX�Ō���+͘p��N�����a�ј9M�n1%�Z��a�f����b�-�5`�Y�v� ;�5a�l�oj {�?�H���9^������sވx���8v|P����Б�*��/~�Z��!;2]�P�$�I�� J������?��ؙ�"�!�8��ԩ�h��˜����b�מ2�=��Ԧ����̞d���B9/��D8��?֯_�b�!ñ6��5����� FlACc���L�k�C{�Y��p4h^��̇���'�N�,����.cbIk�U*�G�`^n���m&�A���ƺ^9�'�<[S�V��D6��>P3�{�W-���@ ��������B��v���9�^z�c�D
�ΰ�qg�o�ch�� ����	(?dCQ=���xC�B̻��S��yQ��2-��jq}�����"8��RN,'9��{tM���oR'�Q�P��a4Z%X.��^����kUb�ރb�3ڕa����#�eH�8'��9�B6Mž:�W��+zȱ:�C�DpU�[�@�����VN��m|m�h:�'�Чh���d�=��c�4��v��$�M9�h�Zu���\�Ԉ��/��M�b��S�Q��pj�5�R�Q/T�/��ADcLr� �T�6L��'SɄ_y���3��t�$�]i�PGܳoV��u7�W�s�38��rǮ�������}�oN��C�·6w��Zx���l���zm�pF���D���>q�"f=��\<l.��<�I��s�|�p��X�<��ʩ���4���F$D�)+����,�O����1�Hg� �χ=�Pk��Β	z-���M��訍_�T���:�e?�]I���x#@�S����6��g�JS���N��G���H�8Q�=a�n�������"�����m:���t˩5�(i�`��b�%!�X���Z`~�K=�ŵ���k��R�5�b�7����F {~É>}�gڔg�=#�K��&�I�H����BW���ocK��2a2%�8�0TpAA߸��ԕ+��VC� ��y����tI��n��m�c��z��n��*�H庖�Ѣ�]A�_�|��+?����=��+)�,#��ǅ�ˌ8�����cݝ_6�)l�Ϳ9����n������:���@�>)�s�8��`4�k� ����'B
w���R_�aw����2|z^����ӥ�i�p_�kꃂ�E��K�j�Εa��� ,��U����w��]��PQQ�?�)|�8�������Q����-�s����yJ���m�����&��\K$�tA�%�㐑n� >r�"�d�&50�YV]GU-�.�NUO,�,�5P�V,LS�X�GI.�B#$JC>Ya��ExA=����˔:�A?�+K����8��b5�ŕ���>~�1�.fm�p4�$��&��b�gOmc$iT��MmL=�/:�}�#2��	�'BGR��WL~�`�D�<V�|;<$@�ca�9GC1��;��:���z��dO"+>����=τ��^�F�Z����>��;�o�o�0�O��������v�����&��w�����D�ﮰ�SÝ�\����Z_$�O�߄��Ѵ����΃�zƠ�ht8z�-��;�9�vv������X\��/��	��϶��av|���l�q���;�Z��pT�S3H��Q��4Co�v�s�4��}����Ǖ��/����a�M�'�$�)=�$~(X%��hW{�a�)od ���\����ҏp��c�n:!^��Z��s*u�hg�0���-�&b���qaNu��9�\��
�{���Ԇ�i3k�ge���j<�,z
�?�RW��y�*Kh��j��A�����8�-�o*y�,�����\R��s�)d���ˢ
��֧~|C�
��3��XW$�����Y	���7���}��(
jxZ8�p�`��Ѥ�m��V���Z������+D���b��AΞK}���ۈ$m������f�����5����)�����j/
īX-�a4aco���i�Q�4��*�q��H��"b�K>��L��yȑAK))C�b��2�~�s������d ~�=tRq�{4��S�M41�n2O%��{�L��&�s�EE:�_�����E��g	#���L�	�.$qϵaC�!pk��6����zC=|(ncG��t���R��s��X���y�e�AQrHwvD�v�X�q���ɅE�mn���s����AT��{��ykX;�=�gy���s��cخ
j4T�bs���H/�O�]�(��2]Z��&��Ԍ��-:���	Ǻ"R�%D�&�!�/�)�gT ��!����&��z�==��=`_�D�ʪr�YGGt��q8	81�����7�wb}e�e�Z�h�B��	|���?��%U��/Oq��rϕI���-)4�^-DMvOJ�ab��a|�r���C��j-Q���E�g�m*����/��a�r����]A}��HSz��A���(\A��ȡ�!�A���}x�1��;��P""O��C��8�T��.�=�!���,�(s8e�tB��O0�rv��L��?���m���u7�W�De�t����~+��� ���:�Ƣy�1�i��=���z��8U�v�ݏ�<��o[�J���P���w⎧~���G�kQt�`yr�����PW�T'��Y`D�3�2A�N�Q<]\#��d��VS��Ǵb���m�	�u��y��*!��4���U�w��8r�D������h��9 s�l/|G�O��ǯ	�>�K��2�x�m�{2�E�I��w��&XPU��V�1'j^���M�5u�C�t�vFhJ���7��v�O�V=�B��WҎ	PfWH=Uʋ�pѰ��
Ȫ�E��!�4�ISe:��@�ꛓi:���8��@ �J_�	�����g3�v��椒2�<��we�݉c���ZR��[e��jqi
�@wa��h
�)��$w�j���Y�s�C@o�J��J��r�;�˰4�:s�rm�ǚ���4l��N����UY^.�k�����\g��)�U_A~��,Q\���҈��	`ѢE�$�R���=�d���k�z��\�%�O`�h��Ԝm;<��mV7��� ��v�U���ը^yeV[Jq]qI).���*,�1��9&T���q�57�yN��mC0;R����I��g��R���q��KǛF`��QYQ]�7��3J����"Y�����#l�<Vxм���Nۮ�d��w$���BZ�/]D�?I_����z�櫉�N���'��}X��G[=17�I�kb���Q�%�4c�]�m���e���H����h���6�=����f�r�U�or�{�e�!1��Cfڴc�L�[��Ox�v��NQ��SiDؙǎQsf#�S��:c:x����{�������:ӎߴ����9Ӳo�:$�!�BNe��DV:�z�C�����0�������v<�׳�� �7o��t��K3� �4�t+C�x�"��Xy#5o�|6��,�{��O�R��Jr4�.�Fj�AM-����A
�ׁ�K*cJ�znL!������m���v��F-�<{�aym<�80�N���eN�=�[���"�By��z=��ziF\�~��ě�j�/3j&�YNM�xJ�O�RW���:��L����U�kX/�G�^WU���r�d"�y�Id����c�Z;���2�
?�}p��9HL�p�'���:��Wj�^��\7��d2 �5����
a�SEH�%BXL��k�f"��D��T�DdqAhe��2+�I�Mgc�y�R΂?�yU��i��^�3D�v8	m���b�H$	�CnZ�S����'�%* ڸ���!��T,*�r�T�~�F!��)Lv9�t��\Q<�LW��ϴ���^<j�A ESxhR�\0��e����1S��~����9A��V.���uRr��iX)�&u1�Z#��)�p�ٹƴ�NE�24�u��
'͓ ��+��3�:l���C�O��y�7ݖ�D=qs&�8AV]Ѳ"Փh��/�F��I�-(d*��-m&��8��:��I����<��"���d��\q�g��,���<�$saKqs�Y�A�BΟ.�d&���{�d?&�J!k��,zL�1�\�a2�i�J#h����N�ua�m��=�Q�ٽ��r�7�Rp��A��>M���Q[���ݖ���_f*�t�S1-{�L�!i+��}V���
�i��1WO�Xw��&3I�\���1����.�ud3�uo���/�m����P4DW����XK��4ԫ��#�c�<�)N1�R�.����O��%<O�we��Rf9'"���0`)r:\�L�L2A���U7К��eG��
�暽�r᠝2qN���ɱ�������EL���x@5-[�ɯ,b����|r��7y���t�a ��}1������9f�3�s� �O���1i��Ǐ�\g�RB�E""��L.f�,Eke���=�#d2�Ho�鞛]�%_ �AJ�gˁR��"�R��ĸT�+�h�Pw<�2fyёd�Q�3���9�x~*�|
q���!S�n��CrsI���|?j��s��-,}��H#�Ф����� �>5���Q�B������wY�D�E��1j��wf�OD�bXs�*q僢6:R��E�W��4ʤ����g�L)>�V��ZG�QD��
�"A+����U[R�Mބ89����VV�q�B�v��J�SD߇���ŮO��6
�P�6;ʛ\q�<��t	q� � ǩ k��^Z����Ŗ6Ag&[{m�b�^8)���b��$b��sj)<qV)ȣb}�)��g��ٮ�B3�I��q� 㒺|����Q��:���2��L�,ۇꯡ$���c]MH]�rۨ�~0�J0S�J�����E�>�����1��j("�;b	W��s�{8+4���2EU���U���"@�}8���G�cǬu�*�E�-����e�N���>����/���<��g���PL鄩^�̳�o�dTXb��"\P��A�+��5˅�m�{ЍSqL4.X����� �PLq�Dȁ~��(�V.D�8����4�dr�\9��k6E:��I��$����3:Y:�ku�1G�QܱP�ѕѼ߯�JL�=X<d�;�1oymO$�g�Fpò"��g��$�6R�cx2z��M�)��@�&�Ϸ?@�k+D���5J�X� ,��Enp�	���B��R4E���Gt����58��XC��:Ǵ�X'���%y�8���ܱ�<U��Z��#:�}����犕��쿂1v��Ek�i�$n�D�D�p޿�&g�n���~��Jr��^���:z%A]�G�� � V(���K[H|Ur/7�<ѫ
'[��R�^0+�8p��#I�5/J"[�D^��p�]1$e�3F\����(8I�?�\�TL["��Έ�X������e�6�]�OR2p���P�:{[��}=1�U�g�`wWT=/��*"l�CQ�#q4Ct�Kh<��h�Šj	Y�ϗL���3��tp1�Ef�Cl��ܫ;䱪���ci,z���q��<YߡJ�/�m���|"Ǔb�%UM][��Ӎ#h�J�Y�)�V��:�7-�QKq�J���yb�qs�R��M���GY�ٔ��c�1Mn�G�K��s�:A�˩Nv�ɹp��i'�-�g�K1n�5�t8�w<� U��[��c8�W@J��Mм�v�SH���j�yi���\�E%9��$���Y)�O����)�2JP��y�_WN)�+.jq��Q+�a���HH<Jlڎ� ��ߦ�ټz��"f"-sm}֭,O�yΜ'F�u�rNF�Gs�Sn�#c}��ջv�N��bAE�"�"�V��wμ\<rh�Ą70�N�4u��+aE��%��<���ǡ�r�t�`�c�q�Ǘ�f��w���1|'���D�S�b�]id6��F�t"n(�#C)��y��� @����pS��G06���Ή���r�RǱ+���*�Is�C�T�O�ҁC�5|良���F�QSq�����Ն�^���S4�t4��*�	���s����Y�D���W-�w-&o���-6ƊZMkl�����|��hV�~<�C�M�M����M�N��U�&��QtȜ'Z<4�� Ԩgt��ꍕ"��^T��Z:y�-�6�q� �k�S�Җ��/�?+�v�����c�+��p��
X�9�#ӛ�$�g���Z��>v��p��L�s�T�(���o;'*H��4�nB_$���vx̤��(3��C�|M<�8���]+K�v�]by	lDFe�S�~�x弿Wt����;�MX�d�KZw|��e�'�C�&$0��<�7D𞨋 �E�(df��v�5.Ff]d9�P���1������Ds���C��&r)����V8 r6���WWW�b��Q��("��N|���V��B�3�!aE���	���(���(?�A�p�T�X����A @�p��*V�9�D9�9v����0.��shg=�΁r�� ��"�����NiN�3P<2�8��F��GM�!#r��I稩�2w���[oI "��=s��t��c���\���}'R�3�$Rw�����m�=�L�{#�#gcl��ɋ�1ǌ�K�\�&�$��r�5�?{¹9Q�CU�ND�"����8�$��㤽X���}W�s�5Ǝ����8�t��\%��;oS�P��ꓙ&��t�Cd�W�CI3�������&',+uV)��ȭܧ�;�,�$�ވ���c������6#�3M"�'|�ͪBQD�S,1Q�S&wV�Oq�Di/+�9bI��Z^�Sg� �g�jWT�F��)�B�K�T��y�������CD�sD����S!:���/�]����䲑2y��L'j0��r���L��sH��5a=���F��R�e���
*>�q!RS��/#���\�8A���f� �d.1y���u
��{Z��@�&Q
����?���1���*��v6|�)�c��9&9."���=�\��B�k]N���:?C��U_� �+�l���I��r�B���6��f��=��1��+��@�CS�������K\�Y]�E('�ͭS�[�S��Nl�8�H��!��g)T��4��A6�r^�M��8�U>g�a��T�;�˼�C4LΣ���.�r��Tnju�u^Vb��4ƨV��.�A���d�$8�x:-ST͹�N����bל$����b����F7�cE��|�Ikݼ�����&��B�l��+�^��L���$ }�T�л��^���:���"�吺ʔ���R������F�)�8c:,�צ3��I.��M"Ӧ�>':���&��?8�^���cҮ�Xu(�ܱ��@����M��Kk<��&�����2g��U���c8�\A_�B�gd7�r�/�|U�J`�j��r�CYk�:SN@��e���#��*���?a�uF�p>�r��Nv�N�2B<�Ek�J��f{��}*�J.!�Ѽe:�ܦ��2������S%�9�'�E/|Py�cps�|S@�g��	gb�WnL�e�0I��Q��4�i}����;t`��ϝF��Dz'�s*�8Y�WS,Ѭ���p�J�kEC�q3anɤ^CNbZN8�}����309����>�:��aV̳-f�f�	uE���I��.��gPQ5Itq�YGIg��M\�$��A$ЙM�M�_uu?/�6x]�+"f �5ӵ���Q�p�W���!�7��ʞDD�q�%	��8�p����� f�1%�2�43�D@.Qi�}Nu��NG9��Fky&�wv;��J�ce�i��ƴ��P~C-3�d��Y�}b'����l�>17�M�>��P-*/�}���Y��X*	U�C�a�+�G�cU���4���ݦ0��!lTv���(���'�K*���=��R>��X6���袧�T[*��Y���)3A�X��)\1d?,�a��^��,�w���0��^'���E{�#n�ZAE+�����>�vJ8�����z�7WP&S�Ӿ��R<��R_��Ϥk��<��&�TYt�Y��e���z�}�F���ey���	���5ϫ�`}��7=dL��P֩�t'2�P���0}��44ϫ��01c�1񙓝;mY'T�odx͋<�֐���)E�	^��!�v�~�e4�xf����i'nSI���!L�qvR���ʛټ��:�d�g6�}&����x/�"�N2����X��
u�N3�b�ݎ��fI�;nF��+����Dj�Y�S�c+}(W��c�Z�����,�3�����}�U���ѱ5Ь�e�����5�ډ�2KR
����I��5�:�(���LΒ��o�p0�`��NOXR�B�'�SX�o�4��Q��O��y�:�vS�B 3����ދ?�x޵�De�on�Ç�������O��޹X�>�\G���mNb�'�"�/+�W�עs$�����ZT)�?o��Ҳ�Ԏ�~��w�g�Bl�x��y�o^\��\2O!���_��>��o_Y�����ُ;^�QH���$�s�>�G�I��8�R�~�6B�^���ksp��R�r�%TV�7v�Л��w��%�[76�,�x�|�jg
�;n�܉��է�qY�Ƥ6����m�~��* ���*͔!g1�+O��޳T��
��C�L�#gy�/���ۨ�~�X.|�a�)��������}N�$s����� Mu�y'�h�y�K�:��7.��I12�0�\���o�Kp��K���o�FQVЄ[����_��ԃ821W�f�%��"4�Ǖ(��<�L��܅���Fݟ���n��m����D���W�êP���?~�"l�?��)J�)�8^O1ű'��B��_j힥����e(�ĥ�������W����w��l�,��w/���.�'M�՟��^��:���&���&6���P�߾P%��գ�0M'�����
��=�*�g"H��xa25S|X�I@���RE��3G���U9���mQ|Pg}�6����G��j]���S"2���"�&��Ay��/���:9��Ib&�Q���j22�g�7E�p̔Ɓ;�+uK���E�E��t?։{��s��~r\���M�6��x�[��M6��>�)���1��<�>Ӏn ޻o@�R��EG|�:T�����l[%Y?xpI��E?�j��������{Dq
E$�p�菜I�����JI����|*U�D�l"7�B,�o�������v��J�_�����_�E"�9A*рOOo���VP(��T�g����bi����)*�+b�Q��XS�RN?x^9^hUȾ�*{Y��cD7�N���~,���xE5��X���#��gu)>q_�B�gO����`O���l��c%	cgg����-dr�����d�"�ơ㚊�"�8R�CB���I�)��N����$���[*q��P���*��xn8n�<,CD���W��[�T	�o߿L=����̯����O=� �C��j��G���fU�N��ߥO*�|�Emh3Q9���g���˰�����7ԙ5��
���dm�/k��]W��U9�9_�����F�F�����c׿{�MM���\��nb�g^2��_D!�}��Fu�5,#�=�0g��±�:�~�_	 Y���OE]��ͬS'`���#J�(ȉ�W��LGr�i�K���i�q9	ݓ)c��o��5�
���lD֗oU�3ǭ!a�0ӎ���"ޓ<wR�x�2{�a�����٦���?<ێ��ܲ��W�s{�hVb�xm���i��3�9oOs�#uzf�T��[�55�K۸�6�w�"��$m��xjl2]sj\��M֜=SRx�V����Y4�wwG������h�09&r�L��3��YZY^9W���NS�M2Փ����~�w ��7�(<�&�Қ�\�����@��>�s�)K��[�����3ճ&S��-�p�3J��B�D�h�T�P�y�D�ԍ�v�J$�|a^1���W�+�T�����Ɯ)n�}������39#cR��BF>O���@1!-���֜����[3aA�e�)��_81��Q�b� 3z�hl>�i}p���v:B2ݓY�\�$���`��?��+sN*.a�6��^��8A���`v$�Z.�ᆚNQ,� Yv�=!��gU�T���d0&@3��Y����u���@�b���EB��Y������k6kcXf�d�;,%�X��0`N�C&�q77�2c�Il����l{�)VÊ2Mm��}9xn��F�6�-F��,�c�1�2��B��$h�{�Ddn*L�9U��L��@˄+����\��ؘ��N���f�EW��8N��`:-+"����SK��}Y���49x*y��!p	�P+�R�������csӎ���-�BB92�Y��Nuc����2�c��0�6�����lSz�[�MA�yZ(�cL�Ζ��z�Ck��&�0M�������i�\��������2��\    IEND�B`�PK   [��X`�/��1  �P  /   images/bc683665-cba5-4f6d-a6f7-879f54c58290.png�zwT����ke�ā�AADz���F�P�B��5�Q�T�P"��@@�@t�^BK"Aj !-�=�o�[��w�u��ho8����9g?ϳ�w����/��� h���!h�$my��V���vI�����KA4�*����8>T
�s����C�U(44T���~A�?ܸ��Der-�!ht��{簬F��١�+��
�폌�TtXjC����ѷ������o���n�щ}��M�^x�}�uWͶ�ߔ��f�Ǵ�;n�~�Q��W��z�4���xŏ�C������W^�MZEǰ�1�{^��9���Yne[7�A� &��{.���u��}[bwI=�"�<n�l�lܨv��~�i#A77o6���ɆL�1����'MR�%j�&����!�4�UF�u���a��U�(��HNU/�"4���`G��dN������z��7T���9��\Č�ق�=eOu�Z	���Rl�ƚlGXYQ)��oVu����k"qz�g9P�4��x�T�ͳ�5!�U��i����#�-s�.�	�n�#�o�P$|Ek웅ĊKoE���K�-;᫞��H���f���0V^Ϟ
���J~��d�5ۙH�^��Qɿ=�Ƕ�%��V�._�|ǽ*?ͩl���-$n)����.mY�3���j�q�0�6��Ŭ儁��HSH$����m�ȥ�Tխ�'9��U���`�J�G���
w�(S/E�4��j��,�/��ˠl�����1��P//+n@�:�TБjgP1y�q�A�m�Zhs�03S��k~ק���SM����~���)ű��ٕi�A�rr������a��Vi�Y�v�iy-L�KTD0��B ,a<g��~oBnr���`[�R�2|�vQ�%��[��f��x�ӳ�/�D]q���;3�P����̿����b���0�jy>i�N����OX%���D��5�Բ���F���SI;s��Mv�qV��.mۘ�/"�,'��ʸ�\h�.C]�����i�ײ�ͼ�P�x�|FeS���K�f��(
� T#'9��(ٚ#uΈ^M��C6��c�?��1�4b���?/��V�*�c�h����x9�Hˈ2�l�1:f�C��ժ	t.�`���8'rVs��ޱ-x�%�X�_��ZA��>x���5i��©LU�
�{}��X|�H�뾒,���%�U�K���s(�������2}����:Z�+
����*s��,
���Yl�$��F�~۹	�2��	v^׮�s�ά���;5���&�0�+"ѥ+rm�ӑ��1�^J$i��1g��1�n���i=�)�T\?�V5�ęU����(��������öfo��dG�%��mmsk�KW�dii.����N���^�5�x�$���5�Hx7Eֵ��<�w	u2YxC=�~��%���F����	��e)�I��~�w�#"[�u;[g�C��z��ZL^4��Z�V��v�w�㬚{{ Q��/��5�p��_gp�0a��9����b�4S$C2^�x'��DbNg��e�w��I<���I����n�p���ˢ��hsl�W����!o��s�����)|�OѢ�t��؛�a��ţ��U��y�>�GzEN!q��\Z1L���|�O�`$�I�BɆ�������{&T����$x�*����V�dڄ5$�M��Dko�tD��)C����!�5ʘ�@aK|�ׇݓo��.�'�񓪮j�1��6|�x�F����G[C��&e�~�]�R��R�l2��};�b{Q��d<:J��Q�}3����mk�
���8���9��<���~��������o1ϊ6C�n�2g�!E>�GsD�?u�mN�|�1;8����jc֭�p�����Kn|�{�3f�<�SD�7�J�jPZI�Sќ%h�ED�M��+똢��[���,���� t| imj��".�_�iܔ������c��㪐J/��ƻ{m%,�̉Hw`n6+�G�:�NJD�t�U}B�0��Z}#ҍ���q޹y(��!H�'s�6�L
^�zc�#���^	�n�Q'���_�+��W�kƌ��cf����,\�����p��N�[�����I���Ss�?ݵN�I�o��I�I������j#ꪸ����&�m�?�y��)g���|�|?:�+���*�/���8�6�?���J4����SS��5���x�N$V�Q��q�!���s�dǒ1%�48����t���J��0Z�PfbvD�Q����M�"bմG�2R��#R^D��+刾E�Um������uA}�I��
�~�Շ��S�u0�u������!��d�n�Q���7����x�|��r�|�ST��kO�d��pf�G����c�'F��adyH+y;]�Q���$F"���o�ܟ�Y�����ck[\;3�*x�X�d��VDVQ��mz��4����A���0����> Ph#M�h�ī����t��[�pQ}���YY�H��EN�����n�p9�l�Q�t�sݦPM'fc�)@bc�R<�@9�?x-e)^
��-e�^�)մ�{���4� ]y1����"2o�@`7���xZ��R^y����olP��_@[I�W�K�y�)ZNx�����^�W�c�(�����Ʈ�'6�Rf����.�o��
�5!�e(:J���׳��VK�;��`�;0�[�x�aҊKG�V��\p���n[����1z	���z���i����/�Vqke0�J!!⮬�r���CJ2	��QNG�E�_J��l@#��^}���C�]�k[�2����6��]隙�x_��`��$�ʿ�\G$�����X�f��I������Lq�H7�>�D9A��-�G�ٺ�g��Zi㣊�� �3�[5�P'I>�ּ-�s��ӯ'$��0�ϓ���quwg�����j|=g��!��iy�bf|�m��/#��f����M��*	�c�-�=�v�_�R�\�@�+ŧӳ#���=���Zq���#{��	o)

��YK3`G%	�<��2	�6(݋���|tߦHs=��L|��N�>9e-�M�&3���4�C_��쭪
-+���rc(�^$?�Ɵ7w��l��$�T:��{�=G����Ҁ��ŝ�Hn�@·[
_w<��]���%�65פ'��oA��1�&�.E@P��#�ed�u,sǚi4G'�����oWL���}r�Ї;w6ut��R���������T�HGC�_�g�����ltԱZ\�>�tHH�Nir���tq���gE�t���~�������/�o�hfn��~VT gj�������Q��m�����������QGY�S5�z͏b��8�흧���QȂ�/r$����|�x�%7��cR:;��O�<�o����C��jb���y��N���B'?t�Ė]]Jq�R�Ħ�`��_�?���+����b��q������;[��ߚ���*�:g��[��(EB��f���dXF�iA_mT�w�ؙ�&~,�p����	^�8a���^��뿽ɥ�X��(�;�`l�-匬�O�X�H*|�������[��~�S�b0�{�g�ϸ����%3˧��wZ�U_�ѵ��df��pE�����K��e�]c��>��N�2e~�B	��,�Z��ב�2�����쮦�K0E�3���/�D2��������/�w���>ы���˾�j֮[:^�����9�~�{f��d��������A�����wj~Y6��-�jlg�[/,���覹�<ԛ�U.��V�t��W�(ڱ�
LyP�N�����H:�`W�?Om^5=Ë�P粤U�
�JŷJ��4¥�)޶TbK饇�⏌��h��ԔR@P���w������k�[oę��R�8;��+Vѣ��?VYG,Q[���ϟ?G�]�啜CU>\��͢5��S	����LϺ��U��uz;a?�Ϩ���L�Is :j���c�SzM����`xDطXJ��J���J�\"�
�
�ʋ�C�#k��FY~��v��k4�p���ƛU�¬v]w�IVV����Wf�/��������t�ʼ;���ã�-;���|	�OXg��r��9^^�d�Ou\�6О\S�=j�.ѻ���B�ط$n�9ԫ�ѝ*���B
������H�ۙ�vmrM�k?�L����[��k�}Q2����i%�����������A����L8&�Kg�f$�4��2n^�'�\]�z��q�ODw����vd�eK��t�ҵ����l����o����)��̋I9�sM�&'�$<�����F6z�.l�|V$s�2Z����u�k[��6�u��ٳ�S"C1h�����_t��A,n����Ξ�R��Wk��<�_����r�y#m��� �:��2^GHq�ձ�y��H*9-9E���:�ʚKM�VH�J\t��N�#Cflo;<ߐ�r��Z��~3�e���i�u�C�+����a�^&��@���c���4�'������nW7hx��I�*�ek�p1�y\ޣ�Zrڥ����SW9�fy�{���#l�	�a���ʍGV�Ը�m��T��jL�O��4f����w`���4���'"���S��B%׵	�j����{���J	O��:'6�|�|*���h	̧��o�c�I}�֥1��*a=�?�#�}7=5�1���f��v���h�0��1��t�_'�5��jd[�^g����N�H%W���D�U��=�=�S6A7�\@�S^��I����X�5�u��.'\�G=���x"��w��n9�|��-j����ʫOfٝ�3Q#�l�9DW��	J�lX�����'�N��7|L���K���)5*��S��蜜����$؛�ܹ6�A'�ezx���Z�m-��z-;�&G-`�A����� ��*�Ls�M�����U�cA7߸��R8�Jyl�B��Cc̺�W�r@���/���G��FKo	�<���? ��N�E��H��E!��V�XZ���<ҏ	\Y��x<j?�n�ˠ�	A1��BZر�y���ň�	Y��<�%	)i�w؉z��B@؉)�����W	5���@�*n��@m�@t��%>pu��Z+��ɐ�����Y�G��t�Z.s�5�I�Þ�/�{%�h���ex�Y���cd��w@�$&'[E��a�*H��fyT~.P��" 3��"e׷��PE��J�eI=�{t�r��'�Z8$.����!�^��Ō4a��&"��d��if/L��h���W���8��9��݂9���0�)(�r׏��?m�v�ݲ��E��_�f԰D.�g�;E�z]��w^
�u�W�'�=0M/D���%����э�v�y5Ń�p�	�'�WVW�Y�R�GF`?�SޖLXP$|�2��%ZWO���C��6����.KKyM����[S��t�];lj�rkm������K�RX�Yʪ�oR���,���Z}�'���RO�ϕ^�I���s�;���.�ai��A�LJ�)����%��[��T��QG��z�)ޗ2�>�c�.�.El�>��;T.��=IaHlfȒX�賌\J%�|�ر2?zi���t��홨��G�����s;��ǉ����d �w��R �DDKaYʨk!R�蚋nM��q�vOI��`�IE��דR�p�X�p���)�-����B �{!<�yƯ�;#�H�aEP�tU>�{�	�i=[n,�n{�0�5��4������Ŗ�8#T���;?<�Q����{P�3h`:l�񢽓ࣝ
��"���J��W|��K����O�!g�9I�^M��s�h/�|c-սz���;"Pc�ia��x‒Zk[W��wQ�fۧ��h=� ȣ��h<���lA7ԱjF5�a�O}�x��@u=��س���@�(W}ҧ�U����?선,��a܈�^��� �J85sc6���[�*�D�nw�1�wow".CMA�q�I��'O�Վ��i��Lt
����h %��M��`���o�N��c"��;� ��:1Y0q���gtw�6X��]ǖ��ɹ���e�g���\�{������+
����2��o��,���9���z3V����VB��sf'��p�L�����b[� �U�iX��u�X�ɓ�+���Q<���O�RY����<P,�>�X�Щou���_��Ck��.KY��ڠ�sM##�X����b�?��yJ	�{`E�/��w���X�D�X�����U��w�{�ck<%4�V
K�י^-E8酿�yȾI�5@Ғ��8�]���R5&
����A -%��bK\�����|�SL���Fe��Wn�c���� �{��+v�1ɝ�2�Sz�/�X���i?>sʲ*+V�/�$*rXK]t�O8vD���X�z&;�7��!���f��.�����k��,ż�lj�\;��x0f�X�+a�{�$��Bҁ �������@	*q��ɤ�t������l�~K�r9�4��*0ˁ� ���%i9�,<���p������[�1��S���^_\21�&���a+��)�y�;��]����(�'?7�R���]��&BL�N��e���K��x�����O8]^]k5V�����U2����N:���չ�yف9k��)H|l�;�H>���%�ef�`Z���9���3�����X7G�����9]ζ�J?�X*�}|&�N�)��7�bvqq@4ڍ���ݤP�����;�j�S ~�@QUUZ�&HV�*�][��u�D_y�@f0�B���'���T�'F?_H�ZX�Y�t�\8��R���u,o��U�p���t���U�cj6���ܖ���V5�1+��C߂i�.%��%����n���E�	�t�[,�s:��'�� e۪fJ�KV�&��Z1R��T�}�Դa^�r����7����҃r�:��X�R3i*��d��vRZ
[g6�Q���5���D����޽����u����6���|�ٲ�G�Q:Z��^�����eC�7Mͱ�a�K� �� ��	x����,\]�r��/�ݪ�9��e,v�����^���R,sY/E5�<lAa�f ��@�u&G�gG,��`O '���ݍ��x��b�~2I���?Q��M}��8e����'۽�J�h�������-!f���*���ˮ�bl�����(��=}�
װN�5��r��l�ky�HHb~8���
A:O.�|+�a��I~�����&��[{��B��u.�3��j��+f<�\և�Ù���έ�G|�yWu
h)I�sO��$Өw��C����;����ѡ�{c���;'����uc�5)��Vs53������\X�y�HZ@������:!�����5v;�L�I6Y�u+�9ft�̦\s��\��잘l�*�T��>�	-���B �����#�&G��>�������v�l̮xR��ǆ����K_Ձ�}+���W�U�������@�NYQ��k�j`E�WZK�1=i��q:RN)n����H�tiJ:P�zᣑ/P�y�G7����u�ER���I�N,E�Geh�/R�~��v�����P�S���h��	����*}��Q� ��I�̉���2u�ku�O�e��6�ͫ�/���I��O���{���Ԍf�ϥ��D�$y6y�G\A0������ӧ��"b<r���^��J������aAu���8H@NZ��+���� �4��Ҥ�ZM�2�K��-���:iR�n�4v@���˽�v��*���o~�0���%б'ݽ�/�[�&�o��������}19s0�+���@YSZ@�E�7��oR��Ջ9$��L�C��f
�'2������6�vxmM�vi�4�������%�H!\sŃ�.��f�M,|B�̶y��}���ie��>�{�.�|y��yـ���
�}�.)��w���������n��ݳq����P������$
�Zᦙ�HOOWR#�Ck��ټ�Pu�]܏3m-�j�9�,��\�]>�_����4���R��(�^,4G'�>15�1��p����\�n����?�y
w��O�a���rכ�G�7��-�?n�%k��-d����L�矒��w��t��y ��� /����3>\��4�����5<������r�o���+�w_sv/�/,,$�v��w�y�\�����/z}{�`���7C�A��w��őQ��R�B����O�U5.�*m��L��N\$M}j��i5�� �k׮�GԖi<�%b?�^�����.��'LMM�Q`ʣ_��˫��K[F�yuȃ�ѡ~����1/iSK��>}�Ժ�;<Mxu�c{;-NNk��#wi���� IÏ�*���T

¶+V�������g�AѬ��N9�F�8:������դ?��&�:l�mh����k,SX�ۧ/���iɽ��7�`��r�jK�̥d;�%v�_ĩ�Pa|�?sͅRр��PTJ��:t֏�@��嵐���$z���RU)w���|�Kr]�k��1v��,"����fP��B_�mM����R��r���ɨWI��T��Vg---�_"E>�K�*{�����i��(7%��`<�{���Ҿ����x�yf�'�O�0���?r�i�:�J��_Gg�C X��-T�ڰ�:/�q���tqk~���a�E�o�˫4�u�~�����d%uV�����z\�sx� ��Pf���SeQʴ>�x��ȣ'qu
��x��iuӣ��u��yt�/Ru;��0Am�[����蝣�(&�|�Ė�zV�'�y3"qwl[������VC��^�.�|�PVy鵵k�"_�~�S�Q���dy!lg~2���A��v]}b޸��D�L��7 Rs����@a�ֈb��Y�)���o�[�o��)C��1��kT�(_o�nn�;J�'u��v<v���Nm���Y���(iDl{U�]9�-ă%	���(48����W~a	���Qתr!��ƌ�8��'��a��/�3g����QC�ݸ�Z���Á��*��<�v�ك�bǢƧ	�͉ւ�V2���f�0^!�V�w ��~�k9��վ��n!K}d��+*��C�p@���L��Y�9b��+� ���)��i9f��rv�.ʔZ�`�3�+�E��l�Jw�^E���R�}�U�)X���:���c���؀3��8�/�`��d��{'�>��b��s�E���˴��V��XB
�͏t�6`fڭ@�M�q~Fz�<���2-V����5;),��K���Z^z��	�sj߱h�Tܝ��P�(����\���$�4x�}F�L�t8����=b*�޿Ֆw�����H��+'''u���à+3++ѥ�-�%��%w�{�'x�V���6<z�r!H={���~���#hgyo03�L-���@��������*�	5_3���:��dL h�O�Ȫ'R"�} g�*(lY5;u��L?m�`z�ժ�N����(<�<�i��XϮ��a��6���^q#�c���,u.E��A����R����;? 	y��sCS��v���k��ʾ��-�Z���9�RNHH���8t�;�G��0�2�^DzBJS��t�k�/��������GX�M�¡Y�ʡ�ȭ�=�E���:����h8���6��>�Z��l~5r(�~@���z(�/��HMi �j���K��̕3�c�w�O�TK�Ǻ�v冗���RPaNmS0��sr6���1��Ws��X����|Z�b��<8c�3B�@�^��M޿Ȥ�R/dG�Ǭ�?9�ә3M��hl�� �or��,���T;���|>�x�"\�\��C!Y�U�l-2����_|{������s'���.��`��*)ͮE�����~;w2xHp�d%!"!{�(�j����DZVا��h��ﶤ�X�-*��������U�a�t#��8�ؤ�ac��A���M��;����?b�P���k��{�2�O�c��J���P�.S�#:�Ԍ�XL���X�^`�]̈���~X�V����M�7=��3QD�Ejǌ�����������Ld�q�C0�D3�ٛ���!I�^薁��9  ��U�2�%pN1�o{~�1�K&�$d��k�m^]�����<Cty�����N������CX^܀!Z����%d�	X�e����4����@��9�S�@��I��7�y岄x�Y�p-��XC�-5ԩ�6r�����zf�3p? CF��G�&�������t�����6 ݳ�a�����/%Le�7����C��D^.�w�9�P����q-a�����+��Y9�\�+�뛱0#6$��M����f�L$� �h�0(��I��g�I� gdU9`���6�3�3�T�}�6�i�z�����YE?j��,���x�I�����N��y 0�	5�K�VaQV�ʠ�(�XRu~Nzhw|���Vlt2�b�J��o:�N�uБlI��s*Ɣ�?_<i�*bn!�2�d"����X�K�m-O>��1PPk��/? W��|�d����ڮ��Y�92)��lڿ{ҿG0��	',5�6{c��vO���\b_�KYf���DN�� ��S�fQ^����oVf<�II$� �T�bK(|��#���sY�¦P[R�Y�*���:f'�Dz�(K��ULx��Eu8ڮ�m�	�l�r���$|.FY�ʪ�n����\_�3��3/�'�V$u�B�M*{@���Y��$`,)����0N�j�
��s;���0�S�`n:Ժ�U�ܮE}�����/~�Y�i�2�d�����I}��V��n�bq�
~�=s�&M���`� �-4�r=]*�</Mb����$�h�uNZ����;9E�]C�&��e�*F�O�]��C脻�Nt�.�Db��D.�S.��Q��k�ǧ�V��,pN0~�N�@����b�I*VBsC��ЕϏ����K� ���Xz��
��dR��L��3M?+�x`�}���׾����C�J�$dΏH`��7.0�!�^Qꤐ|nU�ݲw�L��sC9��Q�;�^�uk�3���:=�/ǝ���Z��m6Έ�|X�-H�7�$��� rg���M/
B7�>�-9;Sw�0û�=�d��HR`�/
�?
�Փ�y�B��{ǆ�R�`�x����=<����fƎ��M���3 ����[4Z���HϟM�y@K\.2q3x����Q����������F��I���EL~��5l=źl����%�I�4ԕ��U`8�z�5w��d�&��S�%Xܳ�Q79}�js�5��h��U�aI�-:y-'����܃D��g�Y�����[�"j�s�|�Gm+��nH5���;D",���9JC���h����Kp���Hm���Ǟ¬��w�mB�����c� ��4[JFrl�e8��͒@�z�r�F�\XR���ӧ��K-$t]�	�P�hiJ�l��u�jz{\)�������q1ۂ�q���c�=�5!t�Е�,���f�ұ�R"�@�"i��_3��氊p��L��Ͻ\] ��t�֧^Z���mP-`����9�a���{l�����v�_�\�~[u7F�`�خ�3�b7�������� %D��;t��xy}�j
.
��Y�.�)$�D��	�s�޳=?��ޓ��M=C�7����F�-���̯)E��)��
�j����R�Y�Z!NE��?j�-�R�����6�� S��ݰ��;1+*83OIV㉹���)�v;g��ˢ� -�`h��al���X���Ě��o~��t�,Rrè����|7B�~^L7�/KV~�YՋY|^�eچ��h�[���`��������^�"���|*��V��l��R�a�W�\�mT[�A����y���ݓ=/��"Mv#�nq[�K�GӴ�Ն/u�������z���J��]ޭW�Z�_��K�6<�M��b�����>�#k�r�y����$8�f�M H%W�dns@?r��D�N�n���R���+#jX��\��� �lv �z���@}������a�X{"Iu_� 1�<0�<�7j�=�5�tr�z���|�6Qh%7,s�Z���?��/�k���c�Y�3de������-�^K<��\��s�-�M1F;P�5�t��h���p0�_�V���������}	ݜ%�R����QG4�\ON�ͷ�<�A�}�lk5ā��{`ƶT1�	�$9|�&dV��(s���	�/#��g�s����I��I|���y��p��+T;�O6.v�g�IۑC_w�8_�p��sM�$��ݻ7���4!����Mv�\;�_"8������f7��d�)��+�����NIJ�孫�e�1�h��"i���T���F��diV2#8;�)WF��x^/����d���%*%�B��}u� �y����>�1����L�1�����%#��r	r2��������}6�_���g�CohyyY��|�.��w�b��Ws�u�kM�3�Ctʆ�EҊ&��'���L�1�i�,q���&��O�	�3����r�PK   \��XvO�XM�  Ի  /   images/c0f01ec9-b7bd-429b-a997-759c27a1505b.png��S��=LHA��eq'�%������!�5�[,��.\��	��%���_x~{�jj���L�۷�t���� ����g	T�g)�^>=�/z��t���ꄂ����|�ȊC���,-Vs��o��B]���Bu�+<���ǹ�c������%���E���?$4���['J�W��]7Ë�3bq6M>��7��`�њB���*sO���b����炗=Q�ȁ����s��ǽ�ɩU�ͩ��T[^
�Q�+�o����4�R���Ď�׿�W����I����0d��]_$�s�h\��@����UK�_7.���)^l���W.����Dh([���8�<����kn'�������������K�)��|K�pZ�3I�m:i���E�䩩���Yh�| �<E�4E�7N�9��0��l�gng�2��6Z�z��D&i�A�TQ�R�3j��\o�-U���@���.�e`�!I�z�j�V*�Á#�[>��B�J�k���+r�e��x�.�2���i�V�� [�w�,�i�6��{_�G���M�fruq���N$�ɦ�B�r����{�}������/>��W�o,��㹡�������'r��Ƀ�^X�]��T�]*6�����r���+��ʙ5�9���n�jҊL⯻�N*��j�-�:!�#� �=�gO�Eʡ��V��]�,�o�F�ڹ��z::�@���L��r%_W�UB%	�^�I��i2��CT �I0�lܩ�y�;�O���ѽ�u���zr�&?�Yg���LJPKx/�IP���ߛ8�F�!o�Yh_z�/V+.7x��i�y"�+{4���.{@�ÿ��;��P�����gC$vn�g5�To)(��ڢ'ssseJ\̮޿�.1vMw�2�l���˳R;W�Y��~��Y\�h�����V]vP���Y�O�q�kQ?�Ҹ;Azo�
t�V�6t�,\s�S�N\��O�5c���yʼ�"ܛ?�Ve��R�؊����ؽn�E�v�� {G�o��lk �ZD-,"rG�)6H��������0kKKkR�,�����s��kۦ��^���7ͅ3ss� O�Ȝ�y���Y�<����\���0�c�����L����|�_�	쨒�1E�������_���N�]�A��ӽ��:K|�Ͱ#�����<�B��+�����d��k�co��)w��'l����f���~������"&+t��o���c{V�.���G�&�u�����g5���K�1���b�>����Pb	z�/�_�_\�-��{��	���ֵ����K�������p20I��:"�i{�y0e�i��n��e����Y��:xΣ^'E�=�*��/�(�(T1�̋��YeL�ރ0QPjXx���VL_T}zݤ_��ET��:��NO<Fwl00��iHt����}�r�����D�Qډ�l�	�4Y<�rq'�q�]͏�Ȫ|#\��1e[?��[||��Y+��O���V��@4�*h�Ěb��ǅ!�h��Ӓ��NjE�1��,u_;5C�s]^�5p-Z���t�;���V�x@���/\<כ�x����K�;�w�߯2f�z/"�M��r����)X@�+*��#��W�m
s���P�eS��8=�nC�{���i�t��a�p�'�*���1/�x�������o#w�sV��֩�����ۋ$kyd��F�|[\���@�G�eoݾ�����z6���ٲbU����H�Y���Ƕ(��DC�Ԏ"���B{c��_��K��z������*�U\�"F���M��p��* ���XH���^��޷X���'kD:,���1�i��U���e�A(����;�)�����c7��Q�0^�S�c��}^��FmVJ��l��n�$�n�x�;�&빷*z,�_1�9+uU���q��xB�䮋1e]Waӑ�ز�@�F�Ć���
�4;n�"x��C�.Pz!���u�^� ^lD;2���

��21����'p%M��s/w<�d3���f�����M>²�s�#|G�c\�g�M���j�r������-�@o�jup�z�_�UX[{Tu,yk"I�˸�5}]����J�.���V.v_�M�8��U��2a(4���s��g7 ־<���܉���S�^2q���|�]l���1$g�;�NS��!�A�cD�ׁ� R�zV��}=̠�����|�q�x��	ZeR3f��������Ud=N���_�ܝ�Ju�3��X���đ�h����ڝ�#��xڙEm����ASK� �ź����}�濥oʻ��G���"��'o��x<0�K��H�ޘYh�[̝���ὲxi;�3ۛ&�K��ҿR@�E#+I	�Z���`�B���S1N��I�㓹<�a=8W�O!_�����`$V��r��d�	�O�������0Qf#p�c�ڛ� Y ���@r����5�^")���7d)Z/E��>f�C����~)�,h!!v��'��p�߼-(�֗k�1z*Poj���]��z0�ΐ�@�(z�O��M�$� h���-���Ը�(��\p\w7&�V�].����_�O�
K0�4�=�Z���r�g�+T؄���Gu�xp�:��^P��Q�Ą_��t�@�#�l#��&.]��qVJ+����e��Bz��=����;����9nȵ��+E�%������.�����_��Y�o&�m��İ����S�ͼW5͇b�r����roJJ�5dh�iN�VJ�`a�X(=~q5Uzq>XU�	�a���D�pdp�Xè7H��w��5D��ʩ����O��5�'�DD|��1��jI{���j�p��y`Ǩ�;w�!I��Y��м.�k	Ҝ�ߢ'��ý�����&ˊ��?w-D�'��������X� 	X!v1��"�n3�(�f�����g��1�l,mKe8���K;F']&�La���:"S_E����TSv�@��6�PE�%�����m���}*�#���RZ�&iC�'k�ff�����F�%�O��r7�,��na��f��5� i��t����;��'�W:�X��w���'J/�t��e��Z{k.���F����N��r�G�5:me��4�V�#O��CN�a����׺S��`�WO�My2l�6U�:T=yܒ�����ĕ����!K���z��V�7�k2^�-vt��-4|�����Eg�>J��$2����/��KW�Zb��@�����C�]����Ϋ<h+�j�B����ɮ���l~/�F��~K���4d�'���o笯!$Ύ���|J�+á��9zL���(��%`�|��f�[Ƨ�!))=�����^k��ym���Ǘ�`2�֋ԑiS]�mG��L�j�-zZ9f� "plP��N4��:3�w������L#�����3�ܞ�bV�����}�2~�Z�Ȼ�P�&��|�/�œMg`���x+x��e�ڱ��̯�D}�?؎d3�rO� ����	nV< ����q��^��y�� ^} ����?Ǥ����Me�Dѣ�I��UY�=���a��)>�.��Ljܐ0uۇm(Nv���l���d\j���krc����h3�[-{a_����mD�����hTUZ�6�׭=j,�UW.D8��u.hWܡ5�r���I��℉�����0�g%��F�Q��#v��~_*��ϡ�ԧR_�jӊF�oE$Go+�;.���lA��ij�,�MmqW�d�X��CYo�rٌ�Tm_��i��_*����ҡ��)4����]���l�������v�D`Fّ"���}^�ܯZ��o�⣷��b2*�52H���bhŨU�m�d�	��K�P���6�4��aٜگ�X��b���M	�	��������Xc��/|�`�F�v?0��ݓ��0�U<)�O�]<�Q�"����h����Мou}�s�����S�^9?����{�]\�$��/���Dτ����=Sl�?;v຿'�Uc��Ң	|ù[*<Vq�2���U�n�5�Ԓ9`��Ӥ�Q�S�"��5����q��-�$.5���i>��g(��L0��6��f=Nc���߮唗�� ����q�:������Y	^Ĭ�E��%h�H`����W;�iBe�dB2�֑�4���g�@,��SML��!�F��a��A���<a�@�W��[=_pȱv��]2Ў�Jͬ'Lk��^Y�;<����j9��q[č"�'P�sm�97�d	{�,�6�>�~��x���U�률?����v0�J!L+�B�BB3VՊ�=d���&N�/	!�|�/�cI�ۀܩ��\)]����
@�#����<g��v�U�Y��)��bHԋ�AW�0L����v�)wN���bI���'�e��HIm�pQи�||s3���ѹ��َ�����f� �79]��M���0�k��6��(�����^��z��͈���٪�=^��{���M,�}��Y+!l�F׀!�d���IR��L�������������mv��Q�wH^m�������<!/�,�Ɋ�d(��#>�18�����6����:h��/���s������R�1� 44d���Եut_L�����>�8�����V9��hiTYfV����C	�;1��^) ���7������S�u�\Ӯ}�s�9�Mޞ��^����2����ʩݲ�&&�ti�w�ّ�N콶�yq,�F��Tz�+dM	�I�$Ǭ�R�s�$�������@���5��>�欍+�d�����
vaAa����1�\��.�)+�Za���j�K���7���B�����]��j�j�63����Wt�Z{=5����t�Nx\V����Ol������l�/p��1�:��"闧�a5oܠM�0�ۄƺ���W�[c����G�E����:Y�;��KF�0���&�o�*��ՙv�}_3S���z�>��&���qhȼ��GmVi�eփv�a�{�b��	�7D�ui�r�g���E���h�[�������枏�'�	;���v'��f�8{F��'0�&ݢQS�����|M[�|�03%e�RZ(�lٶ#//�4?4�؁���W*�j@0���.�T@�Ħ���ZXz���$�H�H�bv����~��J~R&���U3�tי��2&��M��{�J��(̝���e�lm{k��� �\�O�#���>���6���q��R7��5TB��6EPP�>��Z1�jD�uv��Y�����F��RPd��YDC�ݶ�u
Q=�NaP�a�L�xG�\���i6Vm��/����t<�jFl_{��j1 �=�����7'�������������?�ث+��<�Է'54,L��E+yߟ�Hn�$sl��M�5h�+�&Q0�+-𹵱���l�8�$��*���B���Ő�a�tלq+�k�݌��Y<��q2�����e®Y�����X�7�D��$��f%���9@�gb��g�v 8��1,d��y7S�s'B�&<�Z�l�����wbC��DM%�����ykk�8��&�"���A�LFӴ�����+����a���q�QLDt��h���R1>���z�+�k��w�X��*SWӐ�1<*=�c3,z!��E�8y�4f�*�M�#�ܟ5�e���fe����w�Lo'j��+d'�[������t�F�oL2��cx�|;.~���������l c=���n��f�.�͒6��2��t�au�����8L����ʐS� %��@3;f�_���Q������Oq?����l|5��`���<b������3}m��+�����'�a�N�z37ޯdu��m���ܧ�k�m��������@�)l�oyˮ^[�+w�K�����7��&��N�Ek�����U���?�e���ڙN���Ύ{��C���v��[��%��IeW�!����E�'&����3tZJ�F:֟����?-"��Hq$`Nd}	ꗣ�,�����j�m��d���*dF8��UM�|�`@�����HBWҫT$��P䫩�D?�cɪ�ݢP��FZfܾ�F�I�����\g�� q����)����S|����I��BXc����T�����h�쯖r��$`�^�e~�獷�����2����p��=X�����{=�=��3�­(���C�r���.�����7u��j>O��o)T9�é�]xb�Nk���>���L��X���[��[�$x�6����,��)%��$l<o?��t��}��v����o�y���´��Ҩ��X���9-M9�u��kc�%K�d�-�@���݌<�
��<
�x���A�qH9QZ��--U�' ,���S���5�]ͅL[�Ck�tTP<ƣ���/�Mh�眳B�;�W�V�H ��'�AU��c���'�;����s5�����[��㉎LIlļ�bC')�ֵ��SVf#\�%]3��I��l��8=�� %�1�w)����������'UZﲀ��o/o��/��(��Ǘ{{]_��\��	�ͮ�q{D���Lo���Ê�Ϭ`l�{�g#@��a��n��?��D��7S�M�䟂[�a��u@7&O�S�X��-�4D��ZOiy:
���C]�V��B�֢M���@c�Iգ���&��E�e:�M�TN�8Ǥ�fױJ\8���	���[?,,�V#��'s��O0��o��on�Ȏs�o����D�Ld{I���B��e�v<\�R�����ʹ�d��l=e��j���Xp~�$M�w9�T������=�݅$6RN(]	���G&�E[r�=b���+.8�fj��h�c��L}2E���ן 2�2���5s
�F`o��Tk@�+��6�'8�"k"��e�;�l�0Oݎ9E���A���7���
�CG����F
a$�9�0��Ll�� ҳ��,dh�F���=X|��@���1�#5��fb�ޣ��i �_c5tQ��_T�����@��)	:����Is��`z� �j�gxe�3�aS�������1��ZWqO��t���A���a��⦙���
Ą�_��:�M��$�P�M�	�p�^ו9w�ܖ����:B�[�y�Ob?�P�����<6��_l��d_��zoj=�WX;67��(�h(��͘Xx�:��7���+;�ė���Jw��	8�6���~��9�����n�"�h��4{�o�?��#�u��t����� ��[]z:���`�V_���a!�I�nM����W�Q�Nh�9���?mN�$�ׂ�P�����������h�t 5�P��=�V�'��F�v_ �(�����CñϽ��;���f�&�2�k���`���y�4�;I|_(2�'X����^22�]Z6/�|�:qX^Į����G���h��c-XRg隤�c/�:�����0"�"_�Z(����%Jr_�*������L�֮y�}�/��� ����sT�IO!��Ĭ$�������eR�GW��X�6ES�}�@�C������zi��� H&�C�y<Є�R�أ���;2h!�o��. ��w|�2��*e[r({E�}�+3�gwM�y��Z�P[��i+����Zls�"}�p˜5��pk��-�RC!*�|�z��Нt�%�>{���S��#�MQ�v��:���{ykc��_��ō��anE�NX��s o$��vA�ֻ�Y1��t��"�8s���SCv��N!�gDHĒ�)t��E-����L�,�龉���ndD�Fi#�N��z�n�"9�aW��_QV3�>�v"e�^R��Ԫ�[nᑂ�/{X�����Z_����t����-$E��l��3�f�W	�m��e]��m�n��ƭ0RљR��G#Me
��O;|�r�MN�Hw��wl}��"n�x�8�ˑ����:5�ޓ*}���*���:+�y%�^�F����zOt�u���e�tl|j�'�P��=h?�Tc�"4��Ԅ������moݠ
,��=�n��	D
>fP7��Si0�	&����8��O!�#��0Q�Y��a����b�,;/�['���͜;�Kz�G�z�_��s�f��ףp�\�wv%r�?M����ց��_&F�z�D^�h�����c�S��&�Xq�ʦ�aK"�g�-�,3�ںZu��3�
+�m�?��Hڱ�����r���G�a(�}[�Aa�~�h��bt0J=�M�gI��_Sέ���V.qj4�Ό�[;6AG1V�VuF!��e��@̠����P�p�.w��v��N��^��\%&��<9������k�6�N���{g�t���=�4�6W��}OO���@��]�z�SB}�٤6�T�Ti�_��$i�����tXmR)���;�'1U*sC����/�c�mE�z�*y�M|1��]+Qt(��T�.��P�NB��=�n����l�z{��h@I+h��<�\��ښU ��J��3�Y?&M��{�"�D6����c\�`��h-����П���	�2<ݽ֊
����D�:: ��L})�r9*G��Z�8����ڠ� ���>�Ghh<�2$}��d�&��(�����}�w�k�)I���B�:1�eQ#O� _67���p�A����
�dz��$À��W�i�iƆ���<�Ѽ;�wJv�}� ��Gj]�Fi���za�ǝ8�h�X�:��U�S��(hC�wY�aaU2q�v�*ޖ�s[M�/I]m��,ϲ���y��N7wp���걠��o����������{K����_�$F�&f�瓍���(��.��k[1wi%u�xF�U���,�=\���ܣ[�i����w�㌊�w�{Tw� cŝO�A�[���f�@\H�Uy�5Y���i��/�T�[�!�YXtV|�c�$�p����j��䌣9f��^=�Q��:�ztM�H���/�K��������y���hWW��V�?�OG�遽�Wv�8W��Q5�*�5n�&b����������3?|%O���~7��/O���_{'�)�	
0>C�@��� n�J+N��<c/�L�(�N��N���rQ	��o���~��K׬~��ѫ��ⲫ���Ld�ޯ�:��V-��D݄���f'B�C� 規��A�����و�@�Ar�q�N��͙Ru��!V�G�� ��(����~�摒�Պ�g{w�|�Y�/}2��j�~�\��( �q][���oe�o��W�n�N��o����u�\QZIl(��=$M��ۅ(��v����({8Ȝ�GL���R!�f�A���j�z�U
Ly�Ҏ�w��ҋ�~��b�7���(�a����u���6�.���̏,�O.P����w���[�_򶛊�9��٥�G���w��E�D���� s"i�ndw tp�vn���.��qM �m�OD�,5'9���/u�ӒwT�_�g�����\!�O�s���q�En�Y'-�o������q�<
�3�<��'��>*<�K�-U�Y��B��m]�����?|�Q*"�,i�x]�v{�.)�a1�ki6�����W��>��0.G|ݴ��Wt]B�e��spl`��-lg`L��EO�c4�k+<[Yn�
[�;�d߻m��z쥺˭mi1��jm�i;ޤZj0���/}�̋��%�_�wv/vF�z��t�D�W�����H�c� ��kt�����N�V�.��&�K�Nc�r���-1�E��yI�7<g]��`�Uu��E�ZѺRU�(���-���1y�Ma��bL��J/�v�N�ʌ�C�{��Q
Ә1)W��,�X�v -n=�a����[Z�F���:N犚{Tg'�ae�̷Z�o����5N��E�]&5�X&_*җ*5IL������v�1A���O캷"�%<[���������[��Ŋ�B!��G������Tm�/[�O=�C���9p��)G}�f�i�%�ȇ{�-��ݻ���x�"�G��V*�H|��\�6Qo�W�Y��S2�)�g54�����k���Fubs��(*
��������Pݑ��R�r�x�xYn|�9���[w�Z���\���K1\��%�ӡz��T�o�׆� �N��پ�8��[
}Db����%��o|�D^û��[��d�n搤_{�Y�ҩK����g�J[��)���8C�G�(1���z"��5�(�J�n�:����s��	����_� �כ�э�Km��/�~~~{+�����J%ZTj9�������g��Y�_���c,�	�����s}��D��JVt���!�=bTTk������,�2.�v�)���Oz:�SҾ�A�Iw����z΋�,���5�6*�#������#������ˋ�>���Ӿ��k~���E�����{��[\\���{��O��wFE��nvA�z����mT���d�NYO^r�����~�U<�Z��'��t����7��]W���L�xy��|~V���O�l�zᦑ�#eTI<di����Jg�3{%}&u((��E��n��� z^�lŐ�Dׂ�?����^̞n�X��6=�D���U�nn2PRP4����go,���i�f{�������ā�kqIl"�(Wt�a�3����RO��j9��I��4�U&irU{ך���D���"��q$My��I�WOJ�i�[��٫'n����m��=X���蹴�[���X{Xي�����*��"FOY��=����q�$M�s+�46��ZK�<)��L7�hj�(�J~,�7VqKd�e����II����fy^6�x
I1�N��Kym-����ʹ���<U ޻((� c��c����=�F���޽�y��:���P����ߍ�Ø���0���|����\�xG{a�RK�ڳ�+�Z����������S�Я�̠Z��>D�D�k陝7�C���0S�|���*w_�L9�%Q��Ŝ53AJ2j����æ��_�1=̇�_>g�b�9�58�[��fP�Zۺ��s���:�B��͵_�]]9:��Q�NI��j�矈Ѡ���'J�s�>cB��.�0T���֌�t��?ޱ��d�ϰ��98Y�e�lY��,�;X#V������pN�N/�}�2�DU=DAz����`�G�ȋ(T�E�+�U�|L}���(������I�L���/�>��"<C���Q��μ�2�� �c�'s������k�CX���5*п?A�>� <��>����ߍ�
=�G�kU����' ���	dZ��껚���R��K�Kww���x�� 4��/d��eJ�p�}U�I��P��o������nv,�ZF��Q�>m�`�)B+�Yt�*����TY��^��n}x���O��̛%��,��(�v���momYZ0���q��T�ǻ�]#fjU���n5�&�U�O:Q��v���v�f��ux�M���ּO^[ O�R`
�q{#���I}��Dk� s2V�XlM�p+"��o_��SO[�v<^����郍;�����t���P�3hhc1��K T�LM� ������`�Pi�1be����4�I�Ӏ}�yI5����H�槡%��u\��R<%(X�,e��+!��Ћ�0ZENK���x�bPš|��h.bVFF�v�~%������_Og����a�@^��zi�J%�L��i�o9�ت?$���/1��̈́%�r���ib�T�7�V���K����f�wFÌ��dH)̜'����T%#�>4
YN��{��55>Gs�D8����W���
�s_5�a�**e��2�Z��{%���O���wz��ͨ��;Q X�ˍ�Ә�%��.� ����R+I�d�|��12���V��L��ОV���H����T4c�k��NjY`r
q�Su�cB�<[ۤ���1J��~���`�ڊb�H��xj�Y��np��}w>�w�ܓ�(���s%��fD�`��V��}mQ�J"�xR�+�k��U=L�E���l�_�엢��n�Ew��r��⯽��	Â�skV�m'��N�dT���6�jC+�K:�A�gFW�(2��$m����&F�ѽ5<�i!U�<�{�f���W�Cڗ�e5��0��T�N�j��66���(���t͖6�@ ��������.s{u�Hx�L�8�F��+��JB��GGg�����p-�P�;���ǲ��nr]�O���V���C������#'}Q3�&�{��喥<�2i��:�ߵ>���eݜ�5���y~jٺ��i/ܻ[��Gr�T��*�8�	ns���M��G��_�k�
B/�b���;�Բ������kR����*C�a�����턐p��$�/���n�ۡM���s7d��.鬃Z#]���4u�|B��G����ƝOݳV]���ǌ�������k�;�Tbo�kJ��2��*���]��R�ߛ�B��6��r4p������ :K�M�����	��R}������?iU�9�%��ԛA��z����r�Rv̢�aa�ꋁ�t��;͓G�ż�h�Gn��w�='3�o�nZ�3_�LY't7��i�*�@,a�5կ$_ID��g���M$[`z��'���*se0��4����~��А(��M:�:�Ľ!tztf�|n<C�r��d�J�8@y~���Y�FL���*=��v�)��PM��_�D?�$��H������;zz�������Ֆ-�w0#�ѱ~ɡA�M����¿m*�ﭯwi���'~��	
�	�*�%��$»*�?K��-(`��h�J˹Ig�<�U�oD��8ϛ�z�+�4� ��1g!�g�~���H�Y�F�ݘK��,��p�֯�*��{�k�%ٖ�gW|���%\� �w��^�3��Z�4f��꧂�]��5�Hm�N�j�'S��ǂ�'�(ur1�k<��&�6���d�
��Ĉ�PVNXT�E���T�u+оi��X�lv���:0�:+�p��n��c�4m��~cv �ִ�t�����!u�6��}�+q	7�m%iiQB��3=oG�H��p��ܞaax�F�ݤ�k^�V���k`g��:Uz�iJbx�DQ��̵�D%�?����(��&L>4��&�*|4Ts�w�]P9&��9d��1I��^�UWmh%�'���>H�]���n�>3+K��xaE�1�l����vw�e~͵��Y�d}��'~�|Q��[?k UFK�^��M>���o�.�<�H���W*��=PA�o ���Vڮ��I��H�;p��*�ܙ%b�=�a��z���T��=r�w���K�$=�_ޛ7�֮�F@�LpP�f�� �$D�y�e���q��V�+0��-�!�KG)�VK%84H%�x�������_6�����]�:�%*J�*������=�+���j���βC�l�N`��-�������Ό84��Ӧ�F�*R06AE�"Ǧ�{1@��['\�H������^�:�7�+~��;�X>����>>>V���/�D�"-�t4���6�_��s�����7��7Ś�]ϧ��\�7������r:}�?Ҵ�
[�NM�܊��Z�M���{�N�yf��v潇1^� ��@��:w)q��((�L�u�+��f��k|��F���j6A#Γ8)���6p(f�;`�ַG�&M�p���90 ȏ�4X�(3����B������3
��,o��-�1��N?��UJ�G�Uw����Y:�#�p��|M�^�Ve�v`�X+���kĞG`Π�.����X�������F����T�u�rtwgeE���T��U�k$k�.��Ӯ�c-8>Τf!���%9)�l�gy��6�
_��ʬ����9wVK������*�((���7������®����܊:W#'U�MT�M~�T:����3�Ҕ���.�w�yz�d�Y�BW+�*�JM9���9�YS�އ�EP7�w!8\��X �o֜aXV����/-�E�U��b���N�U��bF~�u��������Q��>>�U`�շ*U��3��{~�k�h����j|E$=Z����p�b~�[��p@ā��F�7�7Rb���p�"�%(��[����{��tD�\\4�db˦U��"�ؗg�G�q��`�*��7�ĵ��j��fmp���7Ĝ�r�]G��h�.��>=*�,���W��Y,>��TU��Qv=���:��%o�su��1M�{n<ߦ����oJ����޷��8B�8��{����FN��Į����|4Z�o:O�����Y����g#�QQ���>57�ɖ���Ï77#V�H߫ 1إ�IV�����ăs4W����|����K@�L�*= <ֶ�ݑ{U��������~]w���L*�u�0E�wAg*�v���ſ4pJ!!�
�:5>�,����L��q�ĥ+���!��b���!؞�`��-��ԙd��+���4�c�z��_�vK�H�ծz�~�$*���r܍���2�V2!�b���b*B���-��YRm>%����վ�;�l���/ې�����ϙ����9�_xWƺ���7ec�������&"��.�����Sy�hLg ���te��Y)�lPM���`i.��ƕmp���X ��$f���|w��i�0�De[��k��)�v���P5��r�rο�����g��̘�Yb���6ʲ��,���O&&U�ʁ(=�Y�����b��~��;����-r��)'գ�����(u��p��p����!�hZ���[Py	����!*½��~(�֦�� j�:z=%VD9�� H�B��Ƀ?9u��A�a	��� �.���'��>c�8 ;6���� ���^Q��W��h
vJ1K�|�	"^�'��'���h͙����4�3陭�_ ��AD�T1dd��:�C�:��vw`���[�QɈOGh�ш��jN��j��8�������q��}sQQ4�X��Y��BUl&��4b?����"&T^��"�L�A$�y<���ʵ��=:YP��y���~�s����
�WUK<�p���e�ǸF��Zm_w`(K����(�md�-�Їe֓�L�2:�v� 9��+�qR���p �Lk��5�>��tޓVf0���R'2�{�B}5�G�Z�wV��MC儢�%'��DI�y�0�-�2�Ai}	o6��;�Qƭ74f��,鵞]9fb����^���(���c<��U�w�,�<�-�������N�E3��d�1��;��`��"���j��,���ױ�b�����-8���%�@��6�A�"6�).<�)�$�߶�1����OEm���Fl����v�y���V�q��Kg�勇��u?a��j�~�w�5�9@�:��a�c\U����͖N,��$���F�VW�7�dY�J��܇�һֱf�/�<oi�h�5#�����a��M��v)�)�a]4���RB�l}E*�7��>�W�4t�{xb������υ��˄�iҷ�m�Ya�1�b)�m�tU�vaL���<$���_���1��"�g¹f5��Ő�d�T���FTi���*��x��$̊�4��-`Zu&�Ø\�S�W-�5!V�5>)�Y�'�VL}fV<dA烘���}w:=�N���������A����7:I(_Ѻ�p�fP�N�:�b�L��j18N)�����'���&bqo�&����.����ap~�
�1!�d���������El�ƺ�7D}�Mw��WO��x��ª�uҢ�(`q����I��~�\���+�����q���Sh}�9Ia	��6,�h&!���S�qt�c��H���?T
?@_PXHo�&��[�'@��Þ�����Alr�t��Gpi7����ZP����NIùo��m�7绁z%��q�H�wg#Qx�9�[@�x	�̓�@U��4B���mO�ӯ���0�ı!�qu%�9���V=�4��̂-�?o\��4ݐ1��U�%�;���z�CAx^�\L��V��Ag�j�v$}(��Q�/��)���:�M�57�� /#](�St�)5b���]�|4�Z�c{����͑J4^���#1 �����x�EEz��s�a 01��#����.��mN�(@�cØ��0f�.1�Y?R�����ɬKcP"vC���Mƨ�R�N���慥��/m��>��j.���W�˙[eaN�agN���რzG��62�[�e�~.�����y]p㶘�k���@
�'7�@����D<}�ݨf���F��鏜��K-u���z�Tˌ��u�U��T�����gڟ6K+�����!�.�_#C.~I�Gϡ5���j�#H��H+׹�ԙ{!}�!�0q��c�(�E�f>�&�"H��Rv���&��G��S�/|�.Y~B�>���zn/��ZWW����� uy��X����~'���J�E��e��$����Y�Q�4��*����X�Q�2c�=��^��E�g��#�*�궨 JIwI��� - �ݝC*��P�"����������'�^{����sH1���G�~�@{���9�4�C���A����ȥa��?�&�$=��*�\,9������ma�=,��/	Z�ƞ=��iZ�xM�7�Y�ڪ�)���1�Qg���`�Fa������ë��1�����aVh�j���G|��vƑݿPc=�~D�rj�D��ց�/:/[:72BtUG�wWDM3ޞH�i��4�@�\^����O�!�$�H��NZ�1a[8b����E�MI�g������o<�E��j�V�Xۏ7߰� ��5^�Ӱ�z���1�A�lOG�I|��x�9 �q,�7���7�YJoG�\�Zrb�r~[Г��Hܰ����t���eX	���CC�:^(�AeӋb[��G͑܈�ŀ���2�.�;��o��M��Z�爩e�i#Zce���l����/�^�\�[,���w����OuʹV
1#����Vӄ��go}ԧ���*�46��ȤO@���m�	K;T)�DDD'''ϟ��W����/N{Ènu$�6Ze`���5N`�m���.+s�W���$�f��A��c��K�eh��7?��`���pM��K�8*C��K�1z�ӷ^�6�#��0B��1�%Aq�_jߚ�k���7U���cn�L�g�^J���R�X���]�7�)0���9TTI!$�ā�=� �����IO؃��c���fF�̜�;6�u����!_d9��w�C<b�W��`��|;==�����=���-w��K����҅KlZ�4�X�fK�;Ɇ/z}��B�y.��D�l�r�j�U�U�F5�G��������z]s�&������z�o��Kw՘1����?��l�ї��f/)���2��#�שd^��ȿ����A���!�Wlb��S��>�;4���X{=z�����f(��5HW'����\��� ���C�q�7�$���rK���@ݪB	g�4�cو�����]⸆�
��ƻ�p9yy�	։)����<�5JmI`gw��3���K��	�=�#U
�m�J�o�+��M߁�����^nNbU��U�1�d�z�I�&Ħ��/�$�����A��k�A�8�<Jd_�F��yBif"��*��?�Y��G
�;�]a1֧��3V��y{�y`�zj���diy�P�!��_O��V�K,(ceS����n`�.E�;��P�Nd������L�]	�:	��Jſw���/\a�b�ʅ�R�<�߱~�:˘�<�XTU��Q�
^\��z��}�j���F4r� ��J9����bq�� -wpp�(�U�l�捼�)�8��B�i�s��XB�5����,-�_�8܊�^َ7�Ґ|��a�9����D|�ڴ%e����Os-ˈ�k<���H"�s��)�^�M�vFKG�Ɛ����*����iP�gTmk�̆�j!�z$қ7ma�s���k|�\���#Q
�����b��.*0|�(�=��|�t�_�n�u_��X˃�Ւ��X�M3Ԙ�
$j0a����$�1�5ڐm����O��ɪ�\�K�j�m�JJ��UK{U4S��$D�=P9���Y�po�dg�{sK�A��&c��
��������y�d�Z���ӗi��Ħ�����u1j���
�4S�Z��)Ƈ�}�FӜ�~5N\���V��Isuˤ!�S��ߔG�`"����4u����0���;�׏�J$c�1��-��C���I�j�i�c����e��	���<E�1O:�*�$R6���?�� �_�����ʬ;�	���M�jw1g�:� ��h��Ď7�3�����2���0����EN����PS[K�s��jr�i>���*D*�惤�7�P��цX�}�2���8����~0p��g� ��������B�!���QV�����_|�+<'E^?�$��Ź��n�;��9I��K�r������|��la��ж�T�B��`��l���Hy�߇�/�Δ]���K��
/�޼Y�8KR�������׸u��k�'̵��M+�F�ᤏ_�Ӷ�������;�^kY����yf���J/�s���%Կ~+��@t~Y_{�OaQ������?��'���K�5�_@*f�8]OW��ؿ����mt��q�����ݎ��h��p����#���>�Im~@��.�
�Vf��:��C~�&��c#^4�B���Z��������qީp7����о�{��.@��F[K*�kC�v�w�c�S�U� ƅ+"=�����m@2�/&>l��NV3�m�c����y�.V�ɮ��Q��4�K�^"0����g��P���B���͌�`��0�P�� �x�w��$�OT�aut�
7�^�17 l۪1
g 9-Ē�-��]�5��9\C�X�S�m�*�*���t�_G���Pa�z��t=�&�z��z�p�W`��ޓ����c�O;ls�%\�6e��1k�h��-*K�H1m_�*K�9omp¤��O�o���s���:��@��Qm��[\��c䦫��r!2�sG�,j/�~é?�s�����u�LxV�Z;_�'�Wo�k��	�_{[��J:���q�ޓ>����� �a�hy�2u�[�:P�|���Jq��2��S>jy���r(�01�@Hv��uP�X�~M��%��]�ٚ��w�o��vXo>	l�Rm�k� "!#��o\}b^n�H<Yn����D���f��q3_iZ�V7Uy�������q�)��֔���d��N���4qnZ���9�����P"�A�@��KpQ���	���?гxb����ʟ6ߦ�|��L.����g��~��V���R��yOf�_�'Z�z���k
)�ܳl��s�8¢�w�V�{/Yq��
Ek�������g�؜~1�g΅P�>��&	�T�,P�;�8o@�L�%�j�bէ�}��ON����ܠ���il��8o�yHU	9�pf�f�`,UK�-JT���ji���� }i��s	�AH<o��������5ؚ�R+�X�����Hř�b��2!o��>1��n����cJ��8y����U�C&"	Z��Nѥ���#���P`�E�;߱�nq�V�U���3��V?�Q,�,�5�kj����g[�r.5PҔ�Xh���9;HPQ�^hՔ���F,��Xx1+<�!�T(�m�_4�&��b�� ����u���Z /�e*�SU���)L��Ǜ,C�TW�����:�gek?� 
{���v|o��l��-�^Fm\2�i�i5��.	չ:8(�u?���p3��+�\��sCd��dff-���<�~�k�ߔ�Ԭ���$.Ǉ�F�kz_$;�J�N��u ��Wh.��u�.,-T���'{�3���߸d(���,��> ��J�I(�2κy����X��&=��a�)��o�j�R�&C��朏�a�.;D5��
��#�ݖ|c{A�1.H� z}S냾NѼH	ݫb�}�}��>��R�>> �CW*�h����0V������P�y�|���XS�ݐ�K<���E�dB�YC���/��(������=�oBˢk(	���>պ�H#뿯g�t��#H]s� ���Xɜ��i��g$���Lc� �����(љrh+�'�b�-�F?�����o^J>�A�gq��h!,�]��Q��*�|�Z���K���->zτ����sqi�ii�^ȼ�����zBK�os���?c���ᬬRf]�57��.6��u��E�ء�n�]���Y�0��,�<o䮫���	��˘��C<F�,�,썊&_uxN
{c2uqIK[z'30�� >
����M&A�2@�<7*)B�s£\�#��@�{�Fd�u��8bF"�9��M�i�kQ}�ͬ��-�U,���>G�n�o�����N�6��C�1,�x&�8s���'K�&���y��1,g���uh�� ��'��������K��N�>�_��a��k3O����qW���Y��eO5�C�u�;�gNo���Z�ȱ(�_o2�w�Ѳd�3nX�o��1�5��-X���V)T��L�Y�_�LQvđM�Ǖ(�E�"�T�;�")�VX:�j٦��^�fZHQdD�=?��cH���V��Nl���,lt� P�Yt�]�!��Goo.�����䗕��`ֹ��'����W�C�k��)E�:'��F	{������1}���Z�&ӄ�O�z}���b�(L�]���+��l�Ͼ�;n�qeB�Bl�o�/_2lW���.�6Ht�����VphG��ȭϳ�2���� c�s����kB��ŠD�Q�p��˺�d�������q;���|����]|�=�9"��"2b���2�.�2����m�h�V�
�����aƂT��c	!���F�%H��� �j~n��&�����ғ�R#�h��G��^?7�ւr��?�`SpH��hP�uU�ee	ͪ!L�𫦦�K�#̝�`�L���zĀ���Ɛ`*T���6l��#Z������E��c8��0��yqtZ\^�f�ޒi��&�o�e�rPl��Ɵ��y������ o��/�-�B#�r��
&�j�:7n�Im�eg�G+��d�k�f�{	#i*��4W�1O	�ې."s�d����f��Y�	����~��}F�c�39��t�������l�B��^I=�LҊ3D9h��I	Z�oz��5f�[{zR9�l=0�>@/�uNs�Ķ�|S[\_�}X{ći�6�񕉑�0��3�/�I5U.AO$�S��2%������TQ_7k^��U�����1���T���$3$�ӥ���OZ=n���-u+a^t�l����mm����������o<\���֜�ݖ�s��+7烰����G@�s1��‶�TA��'=����fL+�%�L��Х�e���.�n��Py�Mq�r9MmM��3\털�N[;"�3e�#���T�!b��싹��t/~�Y�[[b�Q���Wn[$؉.�]W�+Yi�2^�T�[����ԎLp�3�8t�="�G���]}�卤)/J�i�Z��(oy�Pmb�;�#M��2�l�}�j���˨���lGݦ���^�I��O��J�cӽU�x�:	����n��ޠV�O]Nx8f^�pӇSeK'���X�O:=YR8ǁ	����݊H.��@��4lXc,*l���=?��<<4OT����	#e�2�^]�8ԿL��+�2ЭM��l�o��n�c�\��$��H"�:yzc$:�����QWb�կ�]$���v�֊
�$���~�߯�n�/
87#�N���EsB"��w�7�Ԓ�:�'R����n6؇�p ��������J����	ݵ�Pʉ��Fd�*��㼨#��_EH�0*`b%]F�$���G}L����Bg��P����I}_W^�N��@��"���~e���n
�ELQi��1���k��j^��}����06iˊ�͖5)�W�7��G�`ii������[�x.��/=�$+M�'�|VG���*z>��dt�ՁH�')[rA{�z�lq�A^�hZc��t�#~���4��[K�oLE,(M�}.·���4����:��!#�	!�_�m圾V��׈�����ӡ[6b�bv`a�r���t&j�Nɛ���`�[/��mL;a|F����j�&5dO��(]�R�$p�8`��O���	A��������l4r)��,��E�q�ֻ�bɣ�T�BM�W�@��.�^!>!^,�5������L�|�������R�hcLh�D܌:DЀͥ��J��QP|��\�o��4���.�z<x��ԗ��:;�G�#%��{����� �ެ�DŜ	���-�DAyfQ���&?���Գ�yg���Ck3���b���c,�;1N��'ü���f�w� ��q���\�]]��q�ʩB��y�5獫�3�߿X��Gu����_���p��k��/�:G�C�&������Kdg���N�X����]'n^8���G&�b���Z���V����(\B�|ŕ�Ё�D<Z�0d^Ga��������:����I%h�Slؐ�T,|���W�QQ�s��(ci����L)�Huw�^�Z��|?0������Ff��(C�@�F���ߢ���T�S�ݒfS⅏�dq��s��͛���Nɐ�^�H0�tܬ�g�<6��zmRǓ�Fvݏ�Cd��ߐs@	�J�?�򲂆�}�(姍\����Z���]]��E��(��U�2��ֿ.%�+q����."��yS&��tVWWK�Abs��Ҽ=^��(D=X�T����
S���R����^2��[+�9�a��nn�����e���z�Z.�_+��>]����N���(Y
�
E}�zQ�u�+ݯ�\aQ^2�lx��~�,�+���'*�*`�r���<bJ��m��Ѽ2Z�aB�U��%O
aѢ���numۚ�����Ӎ��`� 6�V��o����m��ii�Y���=EVKQI�B��E�3��"s2�R��/�����-!>� Mp೿�ԗנ����y����<�����4C����a�y�Ni/��M�.�z��۫�8��'��%�vJ�l7��=�;��"�呟wz��#��x>&7�[��]'
}>�6)�#X�$�@4|p�
�`1Ȝ���KVu�����}�3w���.�v�E���d�ܐ�����Z׹I����~��\Sp�&J� J����%�M���+��Ɠ޹�a���	��r��bi
b;�}X�TGY��ܙI��C�R����b�_�rPo�{UU��}��f]�w��&*j�!�%���գ���K���y�y�s�9���5!a�F� ����ngƤB+t͐r������R�ӳ��H��i�Ph�YVzX�����<��,����o<͍��5/�>�`䖹�`.M)�0��{��!S�K��O`R<���t��<�BY��=��Ta�O��.}��#g�qC�0ms\A*��Y��1���}t�^i17kڢy��`�H������^��#k�lQ歉I�����P'�	O���&-d�ڬu�HM:��W����`�N�ߗ�8l�L'���8C]���	��)Q;��TK�ңPGFF���f���B�6e��Åޢ�L ���y�2��ֆ��U��/:6�PhUK��r28���I����g���W{�Oޫi�5"*�#�c�2�����V-�y'#
�x�?���	h�7$ 7~^�)�m����~�>���E��ei��<���#v]`ȳ�RK���O�?���h�Ζ	�����d0n�������pE~�!"\��rmdl�]7{h-	�v�r�f���$>ux���颷ו�H������#�*���$'�Z�1_�<vaVU�o^,�}�[R��JQr�#�_�t$c��L�c05c�{���R��xֺ+7��,U���RS�:2�_���'�IΜE���:�c؄~�+����,qr>����
���у��T�[-c���&�n�P��Ļ��\�N!7�����;;��QZ�3�����mɦ�Dd��x;���?��bk
ǚw�c<-Ha���6�0-��ϟ��>����\�KQ)+�}�Tόv/�H����4j�q܌3��t���%��n.ٗ��З,�o���bt@��v|y���֞�@u{�FB�!ǻ7��U_ɑ|Y����,�[Sc�D��@���Q�OR��RL~�/�D���z��p�1�..5��A!-��V��Oe�gK-C��o
�����2p�"?�����Ʀ�����f#!(!��G.P�=S����.0�C�B�&�;l�hL�,&�hc?|��٩,+P6f��}��E+�-ji�|ɉ��`�g~7/|K����������{��Z9�T��ur��ec{%�*�u�@H��yv���7��9	����d\ۋ��0�W��M�4'R�q��H�2���#~�b����.؉�_��TȮ�W$Z;�W��6�^�F5�������L�G^�[�/Ȱ\�Q��G��Ť��O���Ҟ��
"�M�'������M���(��׮�I�ڌ'[(9�e�q�0����ol�;�T3-���7aܰn-3�4�n��X�P/���Z���o^톘#44C�p���N��,_|��Qz>�S�4���i�?�W�)%��8�yAʪ�?�ҧ�V�������8�m2�&JQ�e�	�����*��*X�ܮ�ϐ�M���y�ݩA�$�/�����g����S�
�CB=}��7�0����k��x��@����}�G�	@0ɺ�bU��epl�l*@���I\�d��OGb���Ʃ]�BC�ڭ`�N�;%�R���5���dmm�|�Jף&/'����ƒS�����ׯ_m�u[W��Ҵ���<���{���6j17���$�����v�����K�$A��;#RP��6�m��Epᷞ˓ՒP�צ�gP�,���,�8�><A��H&)7�������[FV��������3�ڕ��%gŧ������oQ�H�|��<�J9�����M	ZP��A��f�$r�˜����(1�W511��sC�'�����6{`xDH!�Dױ]l���F�*/a�e������wWo)�ia��dh�Cz�K����G���;���|�aRyl�)Z��dD�56��o�;������Q�v�}�K����ִ`��Qz�ȉ�2�I��^���^� �!����"V��_I� ��Z�����Sa�6�+���W��Boe���~�m"�݁ 2Y��W�GN(}O��t�����va/�\�x]�+��T䥌��y0����z�WC:ӬQ��K	{�)8}8l�h�`�l���R��졜(lTHJ��_i �q�	R ��������Y̰A�i�{��P��;[_YY�7�������Vx�v��@f�8)!�ǯ#`���虎�r"��4��N����p�&�)�J�-�-
�.�-9���;{|O1���/��lee�2���k�ݍ:&4%?�RQ�
ql��6\#0�aQh�'�<<<<�>��Q��ޣ�¡�Yv��Ȣ;��٘��P�����-�ͨȹ%�Ύq:����݂�=���1���m��A0��>o��Zz�XP���YҘ/��*��9��TN�1w.�c�d�E#��<��YN�a2:�F1>�Hw/�kJ�:#�:��~\�pĻ��^���c�06�q�H�#�?���ժhc����F�L8�k? Qk�̈���������P>k�K%������eJ,�0��5�&������7nl��{oQ�*�4i֟�$$z?�	E������h��d���"��F.�@1���ߝ4nw�Ĉ�ڱ�� %-}k��5�/{	n�wm\V����x-�Y���?NOMi���&%�����Xq/bP��x#��`�bN��\�p��h�6��"�^��p4��i EH�"�}؟-4t�m�Eפ!J��Ņ9 �!i�����i;�#M�>�[\0��8�^�x�G
�Y@�}�;�3ꆇ��X�ܽLp��N|T�u�g{��0k����a�]W�BVk��:ZtN�#�����:���*��A"�`???�}u�(sq�J&�Z9l��3_�����'5���Ӎ�_��$%C��)����2�uxq����%����2��Z�-*@ڽ���?U76BQZ�T�����6�1T��5�})�;8x`>���f���O��=6�Rz^��O�G�h�@�ґ!n��S�y�;��A.x�>E���Q�����8�9P?k�����Q���g�1-�a�i�&�)Y6����B4��%>�ǐ��s�*�J���j4xuQ��|vn^����'"Q�<���pF���w,��#��FN^~5��6��<����j���!��A���J����_²�❎����={L�-�Fm]���w�ЍVXC�z-��!�����dyyYZu�/�g(=q���D��=O�F��LK�n��;Ol8La���PZe��[p3�b4�OR6�֋����xZ�	a�v���d�՞��)d����3yR(���<�����t||��_V�GR�3�y�Y������P��**��3+�M���2��'~�寔�Փ����&:p��mq�X���.6W��5�R{8��1�t�,G<��D�Ē�����0O���?>����Tl޹��Ơ�F"Uܞ}L�徺���L��xXN��c�)*��gl��ba��36V�
�~}-�p�����ފZ#���
<��U�Ĳ��VWu���.2�G�|r��+���궼���ѱ#B�y�# O�JO�vƻ3w����*����8-��;�U�7a�rF;�<Z�+��F�\C���{���=�'%V��M+��.3J�1������������޿�������^��spp�����^y|��L`x[j�`�q��:�!a�l�[a�{�w�I�YwyU��aX�ݪ�|�����*��l�V���;���("�}m�.�^
�:�4�v��z�*���f����{e���o䭥`��k��Z�����d��#����g��������s@����x����i�Y&�07����`��h-z���X��c��#����R�1Q5����ۼ<Sx86=���n=啅KX&���6Ð=�}o<�{�"E�3,�4���*��*�+������[L�"��R�^ٖX��- �� *:6����#�����"~g��|JW�k�́��������J�@밐�)?�5�	4�,h	;���W�~��B�!|ck�0��p�D�o�R�'!2^�b���QL٬�_.��xЧ�MM��VZ@�o\���~��}�8���d���4i��Y��7�2�V)� �j#�K�u7LNC�5��ߐ��Hgljz��_CS�zm/_"<"�C3eR�)�G�����9`ؤ���b��?�FFF:664��[R�H�`��U�WA��_�1�j��;��ub�f�ؽ�S����A���T�f44�N4���q�2�_F�ʓ!N�������ٗE��E�^��������*���]}�� []�"�5`{���J��[O�ǧu���T%�mkr���yo�dŚ��w1���%��	����xtMqKI.��]��O����5qR��7[�v�/�j�^T��[t���S�z9}�P�����^~}:����)�pb��A�c{-S������VM�؆��<�Il��~�8�y9��6�=)�Ц݆�D))���Y�.{�4���Y�x�+�T7�oٮ�(���~�	�TR1$��a|������3�L8�ښ��G�Pe8){Tov+
�� #c�ܗA�B7j,mV�����멅-]o�p�����(ABDJ:RRZ�;�n?ߐ���u���]���W�R~	J�N���BEN�Xj�o��ʸ���J��}�d��qJ#���x�0j`{���L$�?������T����=���gX���&h9>������eo�?����\l�3ϭ�v ���V �ﷷ�<q�?%��^E��]�玜�H~ O���y��2�t��㣧B�Q\��b���w$��*02(/�uM]�i�7
�S��{�0��d(0�x�K��d&���z�ax�)��R:�%'�+��[\99�T~��������0	D7�=2�7b���'�M��me��|Ai�\��I6yv��oW�~�ƫV��^]y�Ⱥ2�Ay2��;�E���32Nmmm}�,�|�Kln���7k̪f5Utj�����R{���bן�;;;�ז���F\������{��z`��a��A� [�
�1��n�imJ���]�	�.t��v�:���Z,:BD��}��@(��@:���H
���d`�q�4..�~����uF*�=6�m�m�$B+�e�U�B[�^ݘ>���h��O�A�

C`�=�
���~�"�����Q�z������'�O���()��)8*��gg���տ�w�+��_@������!�8�ܩ���q��\�<�o�ΰV\������N*�55+�a�R�RY���ψ.MU|z�,m_/����p���I��T����|�px��!<cѣ��P��������N�UL���ΊF�u���=�cw�|B���_���?��=�VD�{�G9e�G?�'�E�D�������y�j�7GΞϱ�H��F��c_Xj�o���#c����.��X�(�f�R����`���YmBa௜�o[��������g=zb|���v�I�&�n�G
j��~��u���q��M4�[e׵�� Ml�p�
��E���&&.���l��i� ��a��}u��frr+�ʓ�#�o�|p������d=�Jn>\'�������r��pdG�OO`���\�CL�^_�<���/G~=*#�|���K1�������	CB���,����b����71y?��30�!o�-gZTXxH�d��S	tz�~�_���kh4(���w��6�ͮ��7dٖﰎn_h+�7����9Ӎv��-�i�:�*a 8�P�a�E�!�f������<�A�������`_�����<�i�MR4Ջ���i��ZZB�WB��$�;�x�����usE>�Edu֣ ���S [R��y����.�ޑk�D���lrP�0oڧ#1�l�=<ȶV VWK���z4�|~f��T%Az�}é@;4�i��k��b���*���{ޣ)��MD؄=9��Y>DF9֮n�0�|�'��8�M�'f��W`��}�0�JfU�aa�t9����ܚW���8�ԑ���$�G6��0𥁭��$�y^���67�@�;�x27d������Q*%0'Z�'.B? ��,8�����#�qn�����z�،���)Q�����1��`�[�"�����Ty% ����0S�������z����5�����'M�~D��?�����ð9c[ߘ9��\�-�^��&ҧ�F����<X拁Ȋ������[ZZ:�F� +�h�Ɲj����m�9-e�EY�S��=5�Lb���<����N���|���7N.��w��\Vv��"#�\��}�g�*�Upv���q�q\���~{�b�w�D�xÓ�ƃ4��c��[B����R�?�!�3l���"]z�ǿ����~"����PV���o�1�Im�w Jbl3��D��	����!V��(R����Hv�d���z����8�yтɡ�mHM��>LR_0k'hoonHQռ���o*urv���b���݁��glb��~���?&��ti�/ �pX%N�s�À���2�!�'u��H��)y[޸`a���l��|n�)�Wv�������:G''ρ��S(((�����GGG�u[L�g7@i]c��#{�4.?K����?`���X�������SE.`�[%b�[N��Y[;��^K[hM��"Bam:EF�e���A���������TW;�$0VOL(F.�X�4�3�s�%Ըx}}}X;o=+ �\��'v�%����}$ EÙ[ZVh��/��n6���U.@��Y��!�[� ��6<=���gDފ�"I;Ie��A��(2�HQIIKi~��`^�w�K�;c��nĺ�/�G���ቜh��J0 ����Ӓt ��B�OT�����G|7y
cj�Y>�������z-����2$��u�7�x��%'&_�����x��S8	A�ѐ ��f�m#]��g)���ˆ��>ã�w+�v��"�c��p�&Ѹp�I{U���ȩ���o�fo�5�Z�wS�>b yb��p�=�؎3���W�����L6hfxO���{��t� )n����*�I��fu�z��+�敏7G�Ξ��ÓKK��������S;ٌW�8�KT^����b����g=!�M��F*E��G��G��JJ��W��F��B~�/�ii=v`
���~^��$� ��Ňǉ��rfu<�3�^b�V>�	y�7_.�_�Օ�g|GDj��R�y	m���l�
IT_rN^�����á�!��a��xč�����o��*�A��!b�g�C2ay�w���x� ���E�P�,MN:�����H���..��74<���[�5�?���CS�C��x�%��}���n^����Ԏ/�`iZٔ�VSs>[�R)6�aNs�CT�#|m���7�
A�@�J����h¼8�����؟�y~�G�!-E�ښ�s�8;9EG�NN-66�(�j�
v�*p��S��nӪJ��L�ǹ�+�>	��,�J
B�hfP�V+�Qu0�y
q���m�|-t�����M1z��RC˯��)�6����"I``!"��,X��;����pV�/��;Yz=�%2{Uٺ��P+M/��ȟ	&��5.
���!��+!��z�W^��٠��CB�PSd�}�����6^n���xU�W��1e�Q�ƙs���ua
�`Y��7�Ԋt�Tܶ+w��5�/|p�dl��.��N������B5�ϠY� ~�M���(�z<�a�t��)��ϏqZ���	w�����HHu��I�J�q�`�+�q1�G^�1�D�]�[�bil*�>�d���!j�������p@�daf�	�:���aw�j���8г�޵�e�;=-�k"�x�l����w�F�˒��,�/�͛6"S8���������|�1�?�&,'GƇҹ�Y�-��,;��u���k>���җC�%ZRJ����#��� �foE�W��C�p�2�>.���,�����Vn�Fa�A���V�B :������޵{������(FY*���ѽ B�l^.��w s����2D���B��guXA�����KV׌���Ϣ���L^��	�,F�C`�`�puu�h�O��
!�/ \��I5hvII�&��ohs-4��噀+��'o0VI��U�v���oh}߱��3��E/Q��8���;�c�GG�D�XR�(���95G���c7�W��F.��ްP���$�E(�������i80y���Dck�c���-��+���&FP�ྒྷb�)A�����,�>%'�f�S�`��sڢ�o����̌.�C2��'~X�0�m~.M�9��(_��ϴ'�õ���G��l����ܦ*@����ӛ��g�:|�=�V�ux�J�T���F<2�;��厸����������9⣩�{\�жÇR����;d��.�j��g�׆~ݘ�6q�VZ\���k��,�G���e����:��|�=�y#�@^�ϟ/i�����`}��1z���$�ȑ����֌������D�nsMo�~�/�D�Cd�{�r��x��	��ӵ@�{ ���Z�{'?�ޞ|���͕ϲ3��\�&��J�Q���6z�ϷЊ!��8�ch_��I�~t]�81�<\`V�G̸/�h��O�v���4 a�n���8����RT
�8yU~�UZ�8>�#�/��R��p��j��y= �*F�"U8}��&���sC����V�7�>�����V���KD�!4l�벑-�I"z���Β.a|?�f�pp��>����T��u~q��Z[S�m�`z��O�7���y|~E�G����Iyppt�r�����Sr����tt+9��kSu��\����Je%GD3͵rB#y��w*v#>n�rz����R�!�\V��Ą�����p��o(خ+��v�W̜>E�5��￸������ٝ��yHeE)bbd�)*m�u�)U]�����FsbZ�~&q���������z��v��6<,�*�3j'�I8�5�孤8�`D�lM3;>�b#��9�i���R��5���|����r��18}4*�#V���*~� 22b�)�}�C��8~>����ܗ
r��߉	��c�U� �f�X���c:33�m�f6t��zv�8��Ԕ�������z�"�ju�~���NS�7m�(S������_m�-�uA�~�5[[;UUW�]�G6$�4
��=ģ�D�� JZ��u��m���R~.*���Q�KS�'p�gF`�`��Á���쬥K�v���+���;����u}%i�Aֽ&r��
[.�|%%�47t6ȓ�\k�����=�J���=�y�����<�/�����{�VYl{�_����R�ع`�ޛ�0��,��)�����*%e!@�V|�u�P�J��ü�Fs�g9���+;N^Ӡ�kƿ'ޯ|�{|a���h�����x4�a{�瑝��R2��Y����Q{���tj�!��H��a>Z55�[������B�<�m��Sɓ�F��L�Sr���kU�k�i�?�����^�܌t+�"���XB�
�ښ٘��&}��v�ƈ�,3$ L�4���/s
���}�f���d���7 � ���T�u��|OD�g+ !-'��I��4�Cf%�1� �:),���8�[��떊	�b�<e�����Dc��-!�
���A�禋-l��K��/��}�t�7�,+/���i�f��yriY�S���L�������pc֟����}|L�������v��f�J�"^��4�yC�R�ԥ9L�t��[�MMW��N1zP(�"�}DȾ�SPO\��upo���W��'*�k���"�NB�\�Pihh��Y��6��?�9�Ƞ#����暛������!Yi��7���q�cc;Bz��~Y-|F$�-V9��{���"?n]�z�����`6}��F���4���*��}~/
�5�1Jjg�M�_ug����q�"9"1H�"H�� ҍtww�H7H�H�]�904�]R���s��/��5/X�s���?�a�{�Ғ��Y�y��ll�&���-���d;��KJJ�'��-9KX��;B�t���/R�h�¨��D�o�89O�$��AC7�VV�gA"�0�%�h˕�1�ų��P��Uḿ��jl&hgk�z�--���4��grx2��9�y��-���!g��uv|����m8��*l�w���[�{#�9Q ��~ة N�L(��w��2,1�'����	д�[�ߨf��f�������)~*�<��A��:#��z�"���:5���*������@� �Y���6 �n%��ub%�ծ�	�A���ޑW+>r���9=�/���m���e�ÂP�㟦�����ч���z'D9@-����RN�@j�EEEo߾�a�Ҟ���JRw��@R8X�Pۦ旅��A��s1@�3�����'�����^kWF�o�U$4u=Ι!�����yv<����grDԛ[ej``�f<���f8��0ł�_/�d����DT`�C�Yb�s�/s�)H��FT9!�����X��A�ӎ`%.�� �5~���$���q�ؖ��� �[�o�[�7�QI/�;M�&���?WO��j��Jl444�i@6n }�����9����E�ÈGr��,Ps�� 7�����D�-f�V�L��k�yUL�탞��;��?<9���]����Q͆�g"��bɁ�<>�2<���$$�F�Dq0������3�=�E枼QȜ�VV>�vU=�:��!����b5W0kg��	�n���ݐ�0 L��z���
mϽ�F�:?�WopNG�r̾�����C�I�2����^M}oWN'�(mXp��4)����������b�G��w"Y��"��q��52\:�CSNe�U��|�� ��!'JI�pv�X�[J԰1.�A�'�w[[�Q,�=�����L��t=��6B��>��~W���~���w�E�KH�������R��_PC��b���JRR��	R%�T�%�������Q����X�$��a҈ z���� �JÙ��F����������~�����/|���j�E��s\j�*y��y�>��;,x�A�1��t�#���' u�/tr}��p�� �7�

C؀X�4�Q�6����˛Ų
�X`GE�ݩǬO߄��
��0�2���ˑ�tp��67�8<00PKp��������-��J�,����j�c�?@���JH�;"K:���Ͻ����ա�<����UuX���66�c�#}L��|n�0�@��p̫���I
�/�l^�pm��������.��r��o~�:r1OdRG�7&�����3YЧnzii�h�z�T�M���{||�C��gv-7�3�>��S__�Pi���ko|v�K�},���4e>�����	}vf�Ҥ���^U�%g��a��*؞@MYY����E�#*������Yd߯��\��x���Qa>BeGܫ��X��*��$T���O���;����đ�YD�n��Uޡ��
bR>�O-�n�J~�N�ۘ~�gEϐ�F�pBJ�'~�w'�~��漋u�a�B�l��g�`6ML78�0`�E�+-���n�|��3��*�ed0��^]S󜥼�$o0��V?G��p8��1��� ��B��z� �Tc�:ba��X����nE[�19��׍���޶�<:��$�ܓ
����JO�!(y�N�i�q��g�t��1hD؟[ t���0L�Ia�70�����3AA�+�G7��"��55�/z�* 0*���ǧ�ߴ����O������� ����MMWI���2�)t�y����^f
� ����_��^y�zR��}�a����qO���a"ME1��̴c
�!:��@���zAdZ!���ac��k���Ilz��7dV�4��	Y
�M�bw�� �6����1�"�~�h��4S2��cd�?�*؍��]NN�/�G�Տ��=��>,H�; HG���j���Rk��d�,@��lW2�H�[1��سui���C���ފ�ƚ�R�g�6))�#��KK���(zJ�f���S8,�����*����8�
L�_�p�=�M��N����{	�\�sT�w� EaV�g�n��t^z���kv�|B�myf�'���Y�(��ڇd�/;���=���C<~�������:M`ӫ�w㥞�sjՈ�M)Hw�r������7���{'<!��q���R���u;2�>���t@0{��d���2{{�A��t�#��x����l�˿9�H2�J铆UO-��0O=�u��0�Q^N�{�9}w�$�e�}�#��n�*����#�'�V�d�؀���Vp>���=�b-/eʻ6������շHr��N�ﳝ]C��ډ%ߓ!�L���8g[�gX&bȟ���Mn�>e}���c�5`�QR�
X8{�ˎe���v�Z���F�H�9=����ÞKcQv�
�l�7�^L@�^J�ͼ��nn��R,�������GK�=�eՙt�fg��mK���ˡ
���9ˈ�D-��ڼ�<�OK9O�!9+𕲲2��M�DJYaM힇����c\�ojh�5��\���� Zٱ��]L]���va0X�q^9�Q����~^,M)��	���R�;��
O�/(���jW�PX��q���^�"�: \��q��E\����j$�+:"��$�|_tM&���5�y|xM��[�|��
�*ӷ/Ǻ������Q���l�l>�?����50Th�z����(��/����^:B���5L�h��{�w���II;U���-��1oٌ�҃�N ����w��I��:�X���|��Q�`�"e���Լ�Ȇ(Ƭ �K|3�g�<C��~ݨ�\�睌�N���{��C�/2ѸX��t=����Kq�QA���r��c|���������>�8k
CϜ:�~�Z|-=W<�f�`��ʂ�۞������մ;
A�W��~,]{R���SF��~O�*S�h��H���A��&�[�C��"�0m���7��gvo����K�R�B=��sN��^�.��/ �C���&�7x7c����Yb@���"�g�Њq�ET�(�w��t�+��Z�cbb� ����SZ����,���AR������r�v*�A��=6e7�ˡ��1��7��Tlɕ ߄�;�s��f�����57k3��p:����^��
���텎��M�ߟ�A��ۭ�S쫚�t}�>�a��g�����;����������W���,)�'$��{�����#c�C6��3y!yl�ں~�]�R����
j��Fv��qΒ'-Q�w?o�H��J��������G�y�<�?���ǴJ͚Z�����n�&�=�_5�[&���m�T���9����A��-hF�'�j8�ӊ�𰬐Á����Ն��{�ڹ��������dh�&bKKK�I��矕Q�����} �S�yb� �aLí��iQV3X�qt�xAP{�01���%���dIYY�m�#
���?Q5�I�XCL�	Y
����z�~�m'�]��Kz{y0�ȯ �eB�h�B�L�쬣�#�ė����}�G0rMVV�J����-��Ͷ{7t\�]J>��b��P�����yw��o�{��2/lŀ�}X�����$�C6H�"��R���qcF�t����2��Y���9�ɳ��rI�޵���	�3����^Q\L�b�5#�qk�/��b4���ǧf���{�R�Q`��>���z�*E� �7�O~�*[E.Q�8ݴ��	@�-�ezvc�|8��n�1!x��C�Q
K����cz�h��\7d���L6��\E1�[����S2�?/�ƈM���BQ�<�I�������>`�^&���Ǻ�Z�����CĠn///K��s#���U�:���̴N��S��<�g����|U��yTY>L�e�Ԩ���Ia�S�/r�;�L'�����Ke��Q�lmn*2�k��S�����K�ܮ	�`���]d�]�_'�1<����W�r��>�,"l�S�m߈CU'a=LU����R�>�'�S��l�%�� ����"�@��sX� �v������λ���5eO\��I����t�t[����ˁ#K�?a���X����S8�����zfۣ��+66�g��$�+�8�J0�^��rM�I�!���!@H�2��7QP7E��� Ĉ���7�4����p=	��w�!ؑ��7�֞�+�W�Pqv�ϗ~�ο_3Q(���1~��amCqb��+��g���k��S�M�T��r(~��(��Mܹ��ov��Z{{�@D� ��'�%�ڿxܱ�V���{V��A�zݦ�5JEn񍅏թS�w�W	��K	=�pp��(h?�Zx6��Yk^}=�
�Fb�u�0
T'xtyi���b-z�ɛ���u&�����\�FR!�'`%[[ۦ)��F�۫�G]ϲ�Th'�Dy__����,T�j�����y?Q��ES�n��-���X�y���渴��ұ�z}gg���4D�-_��m��{��;)�0>�QΈ�ME�A��.��Yi�t��2����5??������Ȝ�UF~o��oQ���[1ÿ��b���E��x#�p��������^���nDn��ϡ�|���>~��KR戈��)k�ѧ+�j����x��N��nFvûk�+�	8��j����t�_�h�� ��A�`C?����:�C���߮li��+��|޹��ͼ�<��)�g�(�)Z���0-7��*XYX�;*�b�ME�͡��ԕ�}ƴ�]��Ȉ{�M��g9��1��	��fD�TMo )Yk������d���
�	����L���1�iԪ��Z���S����JG��ul5=?_ k8?m���3��:�ﱟ�vݲN�������il2��I {���� �^�4�A�n9����p�[�����2�2��?���Hn���QR��-��DǞ#ŕ9{ǔ��'��*�\+z�HOO�?L�74��߿����c>�,0u���s���	�`E�k�[i�kV9�!:ޓت�N(͐� ӫ�$���m���
������q����G��m�=��l���t��=����6$��oX+�������BU9��嬳�sş_����>7K �^0�K��-ڑ m�HL*A���\���{3�([���^�����ĳ 	{�%cV��-�?^��];H��Z����V0��mz�<��ɡh�J<�P�M�!wĺЦ�y1Y"���N���8���/xߊ���[����$� X&���F������4߉/���M[H�5�R~d&2u~>��H�6R��۴���O���G\��Y��)��lU��Q�"*����2��M%�>�n��ֈ���e�>M��sx��H��_k�Ǿ��3��E�+�("R�=�IY�I�s5������c��얖�gX����_\\�}2@h�~2�bI܍v�����w�"7�5���}�Fp��a㥇)�Z{d�c�P-�HY��5q��0�K��*��r(d�����SBb�q���G��0l�V��1��w�6ԍ'<^��Cg�&ҹη�YF���ҟ�9��l����^���7Ȓ 7RSS�G߽���_5G�)P��v�9����׬��}A���aE� �Vz~~��o�CmDi�<�oE�~�$E���
)Ĝ��
���X]fbf6��G��.K��XA��S���#ۿi�=������ˑ C�ת��^ئ�"���!���8��|�ݦ�q�Q��0&S���y4��X�#Yn��|��f6͠(U��Ԝx�h�^JT�[����uZ\������R��	2��:����_sA����6���j��yĒ�ū� �򞓀��]��1@�y#螝��
�K|ţ��DV����l$%��c��.��Leȟ0�5�����׳}��,�깥��`�|�I?�ETb����1��U�/Ԉ���E|�{�N|8��)�/���\+����@������r��d��D�Eu�2Q@j���?pP�ϡ�~	��]�yKXyEGՓ�.�99�V��_z���Ѵ}#�{Ƹ��F4RC]��g/#����sX��-+��?Ol��8�=���Ա�񣶎;� ?;^�I=L����>�L�JqX����ʐ�o�m�^ɯy����5���4�r�����bu�r��9����gĕ� ���x���1��T����k7�X<�ɌC��ߧF�U1�RA�p�{�b��zڗUAi��Ѹ���t�v����{��d���L�
�cg��t���g�Ȧ`,«���9�"���-[+���d����(SU@rC��a����H"M��������m�y�3����Џo��������z_����>v&"(��F�E�����{@a�+K�.0��䖤���Y2gf^���/:��v"|_}�zq�n9��
$���F��-�s�7���Y���iy�������ҭ����y��%[艊��y�r��_@|�s�z���<?�����|�=oVmM����(#�?��0>��d�e�</dm	�3��C�A{�ʵ�ck��q{�Ly����h�@!�d�A����LF>�$5>?^ԇr��rwG������e��q9vAN�X����j`�����u�fa�I�`�~�eC��j�����`���}���p����}���y��de@�63�Q5�55]M��D�' ��v��_,�ʊ���2�>*��nT̯�+�	���!�f�܄����m�e�f)�檥G�zB�$�Z̿t�Ϊ��8�Ͽ>-K�ILgr�^\G_#*�4	�%���2!-�����b���ӧ��Pyjcgݯ��h5T5�4�@�`1���o����|���:�Q�Ě娉�?����y̥���G�_̬��ڸ{t�a�d'�P�v~$O���cud��#O��&�������Y2��%�M�?��GR8��չt(.�	s���v��"����)��o�A3 �{�QCcj�WQ�sC��a:�^�~DG��E��*:�t���r��9J�U�@ۻ1
��g�di��I.�S���4�G�>�i�=?�d;�h����+\�������L��>��K�۽ea�"̼'�lX_�1y�.C�EP��F�ST{tO�	c5㘫��<�B��Rl_�݉����y��= �#3��*�7��B'�c��PZ��І+BEO�7t�.**�CD��!�3���7�ȃ*�}Ŏ"���"o��h��ϛ��?n2[A2��_H���&��jJ�A!��_�:|8"t�J��.��	�[�s��<���g�.X��Lx�컍���a�Kj{��90R���EM���#_�cN��Q�9@�Oc���sa��C[�V�p��<�r��=w���������~���ݬTT���
�4�1p_$&%��Y���A��ϔ���\2��H�ӟ�<�9TM���q런'�qQbM=��t1Xv/��x�n94	������ډE�z�\��7����KN��:ߖ��� 1B�)�I#�j��Ν��DDӷ}�⮢�ÎL`P��b����(��1�A����w��9���(��dh� �!s�Vu#3ga"t��>/�ʩ��U��vk�r�>�B���~[����i}�N���W$H2�jrR��S���~�O'����P��������Za���HSt7\���y���čM�LΔzؖ��.Op�H���%����S0%�y���l�w���#kN�:�j��il٨����Yj����	8� ��6ԍ�ϑ���D�_CW��r�L��ng��I4}�����Ou�?����k-"�d^�1��ˌ˃/��U�P"�
\�{0:6Q_�1�W<~���r������4�PHփ�huXy����rγ� r���T���6v�
 ����oA ��2�$��)��~�E���neA-Yp&T�(>����8}��b��B���zz2$�D5̾���KJ��(�@�����-&���cd)����&Ҹr�z+�U�V�po(�i�GfB㽤Mi�Ҫ�ŗ����mh7(���l,�yp�b����	y����'�ͽ�'�Q<��S�2-w8�Gd���m(�Z2�E���"@��-��v�!������LPQ�;1F���i�ױyk���g��ʩ�O؊��#���Ko.���9K�ʴ)����m���e�N#�\i����>M��~�I@D$?W��a���\=��������Ϣb�
~��5�z8S!*��yH���~yqG�?tn�d��A�eKl�A5Y8����fh�XSK8�D��=�C5Ͼx8��fx�*[E6��.O�eߦ���J(1+�]��&��i��F��;1��ׅ������� �&	6%?7އ�H���[�"GO�*'�έ��t����<�hv���ɩ���.g����v�Ã�L�_��i�yֳ��ݴ��`�kK����1�V��X��I���Zf�a�g7������e#A$����	�X�Tt��v��(|���+�7e ����2��t�:<���DF�����U�\�k�!I;��w�L�`���$p ��_śD{vl�Nj��؏��� e%��e[�{ �$[�1�WV�_T�V�(�K1��{�6x�:�6����#����d�nIʫ����e�k���ь��z'1�^�8h�x���	-��
*_���b��vZ���8+�����>P�Т�s��.���H�]<��� �������{n,����9�uM�l��KJQ��Bޣ`�j�^����F�Oq����2h
x�-�Aj^��)KcE�{�:o>���A?u

�h�/�*))�Y���I���J�(��8�%�0��>O�>;c�m��A�mU��b�َ��y�iN&�}�e,��[����!��(�����L�B����p(�����\oڢ�k�2LU���t�NǸ-�rF�<"�HC##Z�0v�_Pi�-�CnQ��r�А�y��BUEl���� �+����vy�fX 畹�1)����}z�*K�~5��r��������G�aX�=��Aˉ"�a�؞C�삦�&c��K]=���NbD��m¨BIX���𻚪�ġ����������:��L���S���G��|�I+��>^mU�	eU��{<����.e�0�&E�uNԎ��n7��i�.ōԯ�"��4��z���$����������hdR�Z�����}�w;S���A"qTМ->e-F`����Ox�!���jO`�M���5ߖ��r�Q���5��f˙r���%��?�����k�hAS��{F/?�������1��߿��խ��%k�;���F�W�J�Qת��j9��I+z�y*D\ ��-��>���wȽw�nPo�#��lI�~���7G��gZ�!L��hC0�څ�>gXn	"
: �ina��\�1��>��t��	�dQ�eS�s����J�2&&��˛�ʇ�V/�STV�"����?R�H�=<B��֬�1Q�xQd�>�_��8�����c�p��D"�}�¿�L�N�~�G|d"�7�_ ��{��謂��TL2�r.���=v!�U�a��NN���n����mZ�jZ�޶�#B�q+t��b�z�	�r����k>g�*#�>�Uʡ��wt���G:2����04Y׽b�P����6CLp��㭍v�Q�KK���Q���~�O�=K�J���o���N���^ߔ��iS�>�5y.9	��NݷO��ᚱ��4���������DoY>͌G����ѓ0D��쀲����Ok._��{�)*�-�����s�!KPU��#��dY�bl�*0���,�Pm�~򓬳ʗn�w���	`��C5ߣ�?�'ۙ:��Z
r=�EXt�c8B�c�.G�.Xb�0#|	��Y��H��r��d��壢A�澮�-C��x,��]�	%�tfE'�{��,����bml�����g��祗�z����Е����R>p	��Qr��155�/�����tH݃�3Rz78(66��&f�]����̦�E�pE���{�0d��8��2o�c�?��(Xƫn�=�D]��F��n�V^�|�
K.�	���ga'�/�r�[�V[�-"e����iôk�Qd�������>�ol̙����F� ��k����Btb6f}��u-�*9��&�:79�K��l�jC������0���&Omb~c�Z�Hwr/�T���5\z�� }z*�q��/��<e�(	��mfg����?����<��»)�-j𭸸8�$�V��{t��e��={
,?�{�U��bu`��ťMT�Qe���=:�s�z��R�=�퍰U���ARm�ye�Tu�6�q5��?CkY|�/#������Y(��x�:�R�����v���f�T�('7ɦ��oN�&�z�������'��& ¨�J�y���o����'꯯LD ��7��ji�2��%u=*>f�v���<R����;���ZW�ċ�t�����C��#H�Sz��湗#��x4�Td����ڀ*�y�F/V ��/�����^2��Ҥ(hY�?���Y��b�lC��:!���M։LV�m��" f��݀j��{ۻ�ʻ%�m �w���E�G�,
Y*%�Dt�ښ�W�Zw�)�S�q|��Z�},�ĵ��~S�_ǥ��3o��G�d]�\��U�|��us�ݖ�X��ô��K/D� �"��J{��I����`�RG�x�|X�nmm�,ƴ|�H����5lY�-�8a�c^s����.��S��^w�UĖ5)h��K�n������[)�;��v���sd[ �]( 2��ӷ§��S�(�x�W��@P�{z�W�$����T��p׸���2�'��_xxJ��vA�s��)*$B3����llĽb�	�h��̂mA� S�,^U�Ǝ7��������v�t,����(<��Ƃ���ʓ���ǽ���6�0����pzz�G�-�	�Y+3��#����4/�.Z�.�YBD��@��B�����L5z�
.	�H���xȤ�_�2z�sMVl��뒇�&1fȚ�!���6aG��*t��ҧ��f�.+WA�5�#�r�6����l2�q�����;>��Q]le�60�Y;��`b'eW1,�� ;ȏB��FP��=E�rY��Y�MB���o���aQ���}qY�S;ˉ��N`̓˃�O�g.xȋ�Eˋ^�����}��p�﯐��L><��Ԣ�Ã����|xFs�������5ȖT|6e�B�6+>�xo�q�E�:�"�V����peQ}R{��ɐ9Y��FbN/�V��nɓ}�P���w_��M�]Y�f��Z����g�[��H�H�Χ��42e��5-�G��T]Ϥ�������SQ9�<lR�BR��ZS���p��.�qYC9����nK��H�g p�H�������z����`��&YxP�b�5x��gV���u��^���G*%{�	�$4��*��ǩ����U+cHm�L����#~	��	C�E�ل4"H�d#���=��pw�/C��1O��5Ϝ�u}��n�{�])�*_[箫�>>W�� >�r�[z�����Q�g��Í�U܇3�b(7W vƭ^��3�ߣ9Y�ßɵ����=�xo�L�MָH�� G�����5�F��,�P�����S�Ҥo5�y���GJtt�6��s�~�3%%1��g��{�[��7]	�=��9�s�] ���O��� r�vh�}��I]��=v��$SJ˵��+8�����Qi�叹������)S潇)��Kn�O}��S�@��xvv�&j�ψ���|�lͥ;�;�<�F�u���LZ�0�L*��'��Ώ;Ŋ9��W�,�[���9���{QQ�Cl�}E�	W!fk/���z��j��hX%����LM����;�r�+W��ڠ7s��^_'ŭ���T�LD\���?�� �d�l5��C<|,����߬�Jm�GLdv|�d�kP|p��EEJE
?���{M�4)D����G�u_c}��#g����#c��k��ۇM���Ǥ�jDz&�Y�Bp�Ԓ��_��H!i<R+ �K�Sd]&�����zX9��<5"~�]4�r5�p��S�<"�N�2��s�t~ZS�.���<�2L������<Qx�H*����b�i@SU��`�P���>�k�l ���5���ⴌ�;upc���~�D�nh6\��kz��g���wD#=����t~^�&��Qj�_@�5�PF��#Gg]nlA��v�*��f�0H�g���ʹc�{i>����GSD�m�J*�*�r3j2J���;	%�ք� �O;񛁏m����c⢹`e�S	�&���ۻ��oK���t��nG3,.������Ĉ�X\��V�RҊ� ����{摤��
	��؈�eD�c��wS#�ieo33<<'���������=)���;L&��T���4�,}�4"f��R�b�!ĺ�-zEN�UA2Q<�� �nȥ��XzA��^n�q�Gc�H'�������� ,>�{~t_�4��ߧ8�#�Xs�;��h��r�����B�*��W�?�p�k&#[[�7'A��u��?S�T��n&�P�LX)t�1Bqx>�<�`q��$��p�}��VPЏ����;֑*n�f��/�%�����VH"U��+���/���h�r�����\6�m��iv.�'ls벞�>�$t�bGs�ċ���Ede�_lR{FQI��u�suյӝ�:c?�?<2B,G�#F�W}X���.��z;ի�>���&Q��ޣt�p1k��k>&�Ev�|�Aя��G�LQk�k��,�铊�u�$��@��>X-j�;�IY���Y��U�����B�tu���������/��?��U���Dvww>������y�3��<�"G�lm%���6��?: ����a�"Q�GA�*��Ѝ������:�P���(�qC���I��Z<=�-�ǉ} 3{��0�د�%��)��q�\���I�<�c�A{���%����>>���O�2�"��6�����l����8� �r����lH1%\)a!��e��л|�܁��Uu���aQ������H��%%���/9e�{S�VF4��r���ބ3��O%w���{��t�({zΒr�Ŀyܭ��m�*�'��7G��HM�O��z�m�X�B <�p��F*rs����\K\^�1�����k���OHL�?�L�y5�)4��c��C������ؤ7��z�/(��".������{9�+��6������c��50��"� 礒�/11��Pb���a`X��`@�.��b�~��D��q��PK   �<�Xp>r�  �  /   images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.png��PNG

   IHDR   d   1   ,�   	pHYs  .#  .#x�?v  �IDATx��|{�dWy��޾�~NO�L�L���<w�v���$#a�mDJC�P1��!N��ʉ���RvL���*Ɗ�`L��Y���Xi%����~?�{���}���힝׮fK�5)��ݾs�=���}�;�������O\��ͦ�o��&X�z]�д,��ʊ\|�WW�ihȍ���f?�y�Ѵ�a�t�6wձ��Ӥ7���}��5F��֩�ٕ�e�k5���0�4�U��|��;���|��ݨ5Lk�g�����\7�k�wBZ�K^����60eT�@���àۅ���fs{�R����é9�o���-�	o0�b>_ �j�, աNT�E�X�����V�����b�PD����h4갚M�<^�s[h^���c�~�jQ��՛�6���C�4Jyд�HLr��N�vw �÷���Z<_~���YM�K�	���)�v;͡��GWu��A�,��'hhfGnkT݁�_{���{�é�/D_�$6�f�r�X��O.\����+��!Ē��AAHoȏr�!T)��r:F�"�ȗ�Dm%Oɵ��W�3Ff����H�͢G~+�$n7<��=r��Yt%�omA����AdWV::������(
0�Qd����P�5��9?���1LNNbhh�TJ)caac��p�d�\>/�m����33�������A�]�ő��ҙg0v�8�����٩֞�d0 k`_c��X\ZB(�a�����ѣ8/s���*Bd��[����~�a�5�r��w-Lk�jqY���y8�=������}�r�C&�����I��N��jRM^״�M>�ԍg����(?X�	��X��	�¢�auy�,�а$u�#'�D�Úb���&t,כ�K]�\�f]�o���!%�7�-ܲd���O`�T=d*1�t8��A�yz�aS7Zo�{xO`I�wI����J���M �ǲ�w�u�	�(Ε�+�G0q��:a\�b��=�����cM~u�.�Wם�����(=-�(=,ck���H(�Ǣ�!����%Otw�+�S�)WED�X���E��R��S_�oL��	�h�Q#W����Hw�쒱���_"@�Zǲ�@Ƕ����Ւ�D:G��p,����#A@�4
Eda!��"��k��qJ̮򙴙�6��g!�+�:|��e�_�Z�)�隅��7��H�\�HG���.����~/���MIT�5�㽘ns�dG�"���
Uge�>�`9�����;�_NB("�]��$�/ͣ�;�� ��ea�Ӊn:`t��?�+�a#� �y��:���T������.�`w}8���� L]*��BT��^GY�n�(�J"�I&̺L�lH�ti�/�Pgy\�w�B�A/2�\���܆R��+��h*u�CC!>]*#�b]�u� �&J1�>+�?&<���%�9�]$�.D�C�n*=��Um¥GEĮ)��ǿ4Bd�Sɬ�X���"���ґRr� �VQ5Bm^4u�b�Ʌ<La�卢m�5�\zt%�A�[K)+����ҥ�B�k�糪, ݬ�QS�g䠔P5������S�H��Z�"�oʪ�69��]�r
�F`r�T�"\��#��(
���� 6"�ź��Y!�\���cT���-"*�O�HwXʐ�!T�9��B,�H6�b<7/�r���]��˹$���ɪ'�ůu�����k��R��w!�K�VW@b�ȑ7� 7ʈvxQ�6�zj�+��b�}[ܽ������BiM�%Y<�m	�P��v�ŏ{�eۨ�~�]�������7�C^�#�Mnl)b��.�����<r�q^>��f�,ȭ+1U��wMY#/�N�|.C"�%��-���K����1d������0ot��#9���=E4�\���LY��7�Z5[�SS�Bqz��l9P�Gm���s��(����^Dؔ.��P��G��"�2�gfWq~=�L���;-6�u�5ҏ�>��Q�k"��D�h"�SĒ��K��|#����dr��b�H4�%ѭ�K���(b"�'��-!N/�����|�{�_,X��"�\.;D��h��p�T�A���qE��tZ &|{�Ĵ�3�6����H�IM��fڢÒ�'E�5ſ��_��\��	c0��B��>(��/��U+-?����D��Y*"Iٖ�E��pA�����*Wip��Ҏ�2Y()C�����R9�m�p���"�0��*"+�J�J=����l�Cd����]���b�|QL@q�j&����+�p��f:���,E�,�b��17��/އ����΢�t(1�]�ؽK��hÃ��N�ΐP�[�5Zh$���j'կ�J�>���t�R�`�7�i�?ԫ�֒��h�i�z���l)u:}��ᑖ�k5��ۧ���C�ug��KMkY���Y�W�R�"?���U<1�Al�L�80s�
�h�Z"uGD��NQȤn�{�/��b�~"�H��|��e[�+���
�!ѣA�\���D��.ie]�¥P��8���Q�RH2���;i��)�V�{{n�������"\�.��B�N���C��bn-�����('b��|�4�+\�oD�}�!�~���2��v�R��!T�y��N_X���FS�Qr��2DDquC*�$����p�ًaKqP�P��2��UAC�ԪR��Q��]>����Fw+e���0�CN�3���];�p�Dφ\���؀\�����0K���$�?��$R�m���Y��h����ex�������w�Ƹ�>���Fb��E&�.0`}�Q���{����������|E(�D�X�Xҡ��Ԅr���sgyI�w�E��gr���ƺnᶁN���1�:�8���Ȥ���8���yg5W@SD�߸Z�փ�P&�Y����$��iM��'�)�ծ�!C������m��CMGQ����:)�˵ֺ{�%�-��s���xj&g;}�(D-���'���.�wee�1��ư�ɪP��Ӌ�5	�Y�B'�P�ni�T���4�e���q̊����&>���_�G��uEB��o�#:V���cZ�coC9�#�!�,��3�Ю�ZADR4��ٲ=W��i���7{GGF�$�/-��4�J��L�yPG�笋�,�v!��!��V j\�p�GS�9:tY�+*��̨�-�t|��wQ�����ĕ"1�:��)
�n/����0��_����=Jw��k�wcp�%
ZEz9W"�q�h0���~�ד8���tFE�a��b����8[�G^(9��{h���ͤe��H��Nn�"f��fE������;fz��=A��r����ZΥ��ٻ]d\W�o!��@"1��X{��Xz���_?�B�TU���ۏ���B�CH	
c���jc�����s&�EMĘ������;;x���um���\Q&j�x�j]��5Ok��ɺ�P������T���&y���{@D�p�6�vw�60��Gw�妎'��P�+xO����ps�I�D�q!���@�܏�?}�P����ٛ�c�&U�ײ-0!�r͂��|fWLr��"i�Kٱ�.J�p����c�i-5���%�uu$�5T�oˠ��H����Z���y�a����
��K���r"��f/��	ȶ"����_�"����R��-T�4������J����/a��3�'��s�����sO鲥�����Ṅ��=�n^e����B"H�D�AK�&z���^UO����"?=�Ӊ��2J�+h��=�D$��H�����u��{�@7ַ�j��g!%o�3�j�f+(�"0];2-�.����8�_��_�ן@����)��!���٭�%�^�ήؖ��3�!�b
c	?�s艉�0��3��(�D=N:j8�яb����cڏ�~*��'��t ��`��h�o�nLtca3�D��,B����I6`uD�ٰPsy�����Eyg�TCI��)qdoL����&F�!��+�w��l��ld���GQU��~�u�\8�l�w�s�i�t�|f5�G^\���k�����3p�8�?�t�h���V��� ���T9
�$d�+G=dk;y���k��فB��V�3j���johT�-k�R�P۸V˄"u��K���?8��ׯ��V�t�զ=�J�ڈ�\N1{˰�G{�Ss+����x%@�{ؘ��RP5���QR��f�f�g5�E�x�62�\ �r��������N!�3R*�j{�~%V�U�zl���w�������%��'��3��Af�t6�̨|�JD�K�q�C���yԅ�F�r=�v��2_�b��k�xS�0HX��Ⰵ����c����RNcL���x�ٗ񫷾�x��s�G����-�".�9��A����<4ػ�*����"\���Ԣ�lq׸l7�ہ�߇�D{=���C��^�TɁ�BH]fq{��w��W�XJ:���k%����5뚋-4�8L!�:�~�����x�,��I�����p|H���_�����b���݉}�[
O�.�t�T�,��WIps�J�!��x=�B�ob[��j���1����&��f/�-�Ft3&�!�nx�`�fY&4��u���ģ,�9~J=�v�f��'^��>p7�ϹY|�k����|����8��;nƽ_~�r�8�K����p�/�ŲP/s�j"��N��%#\��D����xV�8n10�]�!�{�px�������e�n��-��>��m;D�̕-��ב�_{��B�ܩ��_��������o��ď��z�Gg��g2C�p#�]z�B��i�NzA�S��R��D���r��$U�v@���]Iؼ]�W/V��;�콰��b�rx!�_͛��fْ	'���,�������?����?~��ދ�gV�Ȣ���K_���v<��ϫ���~�x�sxaa����#	�[M�	̹�Wn4�)����Na9�)�[-�R�PW��S�s����ѦL�V)R�Y���Ĳ�ƀ��;l��j>4s�̟na���ȓ/�)A���.��K�
1g���R��G;����_S��4-.&Q��>h�������ž��>��*�O")������Q4}����%WV+��6BFGG���>���U�R�v�p�L�z���Tc� �ɪ�+��`23�#`|���M�w�x<�+�P�=�kT�T��)S=��F�SO�,H8=��R|�@���Q���9(�n�޹E��xw�2}��B��c���B��$�����zJ�8Pdu���`%w�Z�1����@�eǌ��ۨ4�D�k�����wu�pa
���na��
�=:N����yL�����{'�VR!)��N`�[@��%=�ɍ���=�Y��'�vּ$�䍩�dm{ϝ
����P����f�w��XIe��q1�W:y��G�����6��M��tv]v��Xˉ�<��J,ߘ���>��8.>
�|��_=�WX�D��~'�ٯ~�H�|���xdjf��>Ni��:LQ^w[�Xv۽�gD�������'�l �^�}��JK��6s�9ж׏�8���,E{�5r'���~���uյ&�guwv�:�p\\<��c�j`u�E<�O��N���6�ʶL�����-<����S}�puA�?�'����W�X�=DH۟Tl�j�۩ ��]��@�L�ǽ�\�������m��I}�q�cv�U��C�N2{P��$N�N����;�<U��4p����[7���(�Q]C����alb�Z}�}l�F���au@��	�D���S�[h�Evg��X�k;^�^h���V���g�-��l�5���<o��3�e�>b�,vZE������C��+����7���9s�i봕�%
��B8UG".��P���JU��fg͖x!P��*Ң���ZU��#��"��Ib�����e�E�im ���X�u�p9�9z��c"��
��ф�:cC�D�`GH�!x��f$��iJ�ch��b��m)hM��Ʒ~�[>4+>�3s+eC���}j�-��$��u����Xm���1������ut��^�BY����7~7�����{���+����9@��9Ãe#�O��?��֖pPC(Ɖ�x^Cѷ�7�;�%\��i�l��:�H�sH���::@��0�G���Pg1��b���BŚB<�M ���c����`��˧_PQ\"�ͥ�9����_�
8�o�)�k��?�Q?��3�U�\2�4�,�x�u�����s�>t�B�erPv"���:yD��{Q��DlY.��ݨ4�0B�B��ya��0�=xy�������BIwb��B.G��h�x�R���G�\Q�W���nLt�{���Xr���S���ʨ��J�0��y�I)~��� 
b��Eɦq�/���g�j��2���Y�C����s�!ļ��,ƺT�J8�}.r�UǓR.r.$"k��;X�xW3�
w?�<��������8�=��Zωǿ!��K���Mv����� kn�d���g��Z&L�����$4� �?�a�6�ؠ��,S#/�V��z����Xb���i��>��#X�[E�j���E���\�����1��Ry��|��re|~�k���L=�`�k� �{Q�)v�2�a�X8�tY�/���@P�s��5�)8�K.>��yq���fϟ���)�(�|���3�#��x��C~+� *�]9{�,z{{7�B�V0,z��#��5ܘD����׿��:1�(�n�XvY�-eZ65���7E��=�Μ�	⚁�|C>~���~Y���$�g�U�~lȽ?:�B0o9׫g�&�v�n� �����
�צ4$H��v_�i��H0�؄Lq}�!Y{�F����9�N7e:V�ί;�wM��*�y}2Nv����d�E�땺��R�����`#z?����
�-?=��d�x�r�umy�_]} ��'7;�����o�F�[��Kr������l#�`0�B����pH9K5��z��133���qL�o\X��)�1��߯"	bũo����9gRI�~��ȅ{୉�|����p��������a�$򻾾����H���e�����o���j��K����4"wߏtt .���a��2����oJ�7�g~[���)�_G�Mw!;J�~E���Z��wO��$a�O�8�t�9r2�jY���K�o�5"ױ7~�N(��1w��v��0��h\��@�1��C �DL�����[�E��:�N�(u=�a1��� ���f�e����(�&n��*��qՎ���G�J����N4�.�W&2���8Rސꓙ�������/q����R/sxk'J�n�$�1Gd������/ɵ.�{��F1���*�\��%�����u�\"����lQG��	�:�0�ힵ���j����rw����i���s��#�8��wn�~�Ĵv��m�s�:M��םb���M�o�8J����n�p�Q���:j�i�*�    IEND�B`�PK   �<�X��g)�
  �
  /   images/c1fb8ae3-abb7-4800-a199-c8a1e0562abd.png�
!��PNG

   IHDR   d   B   �s   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  
kIDATx��\�k���߻��d�dK�jA4F�H\BK��N?p[���/�C�P(n�R�?Ч�ҧ��o�@����UR�QS0�cl�.�lY�W���jwgz~�=������������;s�~��9�s�LBD�O�<�D�B�0#�R)�L&E�\��j�*����$bϞ=b�޽?��o�YLNNv���#dvvV,..�l6{ƶ���,�;*��!L
�{t|�ɓ'o���v���#d߾}��ݻ �;��n��������W�92H��I�z��h7"G�Ç�����HR^V�h���e?Iȫt~���Gt�#�l� �aQ�>�����C��m6�����F?�jK�Eİ�~�O�^����/؏���m��\.W&���������!���bbb�P>�o�V�#D���������
gΜ333�T*}�:��'��h�u��3���=I���b��	D��X,b���v!�o�p��
>pR���={&8Б�G�8u����ܿ��D��d)�N���3�������;�������"GM[1�] ��1��$ #.;�|�����z����N�:ձ�G��+W�xvg�1�T�P�����uk꣏���?�޸q�#m�!Q�sB��	�2D�uP�7a����;�B���MY��۷E�!�<��!��aw^y�uw��!��:>�!�t���'�����ѥ�·��"�Dx��dv����y�cc��4.=�����vD�t(��[YY���L:$ ����d��w���&����(��P[4g~��='d���.ҹW��&�v >YU�&�رc"N����0��r�:�P��ᡡ��r�cI"J�&vtx=ச���?9��[u��r�DMOOSL� cy �H�S͝0
�F����ˁ�V'����>H�#�0Hm�I$(��. �	��ras j��J�!���_��x0�u%5�OJ�*"0!���h���������d�C'.-/c��*O�m�ȧN�C$�.��:�UҖlo���˷b��ϋ�J�a�	�H�(��!��m^�0����͂���P�\I��!0!��8#T��`��ُ�2�F@����יt��,����BH�������>̕4��k�@�jnb����ٞ�(��5���`�7
�)!L4�
��2�'�G���SL 0!<;	�Ӹ�L�I���	�t�2Sf�~eɝ�a��`uez󃖄@l��4��4! :�7��,��U�&�B����4��.B�d�I�m����u����*�ج�;o��@�����J��.�v@�=��>h��@+�v�����κ�iG�:.!~e��< ��?M�t��ۅB[��݃��&o��|>��:jbB]uBM����9��J��!rX�"š��;�{����G��6U144$����V1�׮]���T�g	Q��TWu���ctl__�$!��q�������c/^������!6�����t��9}	�"��t��gGVΓ�;$%����~R}������{cjjꗃ��� �7M�����oY��3�.�:nCԭ��N�w��Mˉ������$=��e�))�f�I��`��X�G��g"�W�.]�300�aGgY~����_Y��� ǹ��s���]�X^��xNrT�K��xK�V�U���1~�lB�y~�h��Ż���;`�k\7�Ћ�Pw���z;�M���8-T�JKH3R��dB�`9-Bt��mZiK�XH���u��#=he����K~�/�-�D�W./���4�W$;>�m�����x�r@R5�|n���!����!��U����9�V�??�mC�H��u��W��Z�F˄�$��i���v��V;�����*�<���cx��6&��sq���"F�P��':�`?��OB�#BxB 8��<[Ӳ!��� OL�#�-�	���dI�+�I��ȟ��6ꬲ�V+��2	Yu�/Gk���5�!�kE�C�:�WiYe�yΕ6��D6��m�0G����=�>��C(���5ǳ�Q	Q��F]U���!->Hû�ePG㍫?Y��5;��S	e��T櫵r��)�#B��$�S�����E+���)���-is��CTP�Z��~�����6|ޟI�*"	��B_��7)��ׯN�<�/����9�8j�!�mB�0��Fj�-L�Q��8z�lI!vw�w�f`qH����fg��ŭr�r�5 �~��Y1���������+u \k����u�a2!��N�:�\�{�m�N)�D<�X®�˗/�x���m%>�QZ*�ga"{�&�JHPpI

+�Lf�}�K����و ]!!rX�$���Q3ݽ���9����SHR�I��%�7Kk��d�jB�3!�&��u��&�p�~�\i��E;�ʌL��l�I������#5C��l�oT
��m\;�]�����׌j1M��BB,� �
��8n��{���!�n&��Hㄔ�ٯݲ7^v�Tn�qJJf��,�?	��{6M�]��u3NȾ�����<!j5���%���p�-�M��m�	+�z�R�,��	I���<dD ĉ���P�\+���:�nW���t	1�.�T�R9�n�B}	q���|������۵bص*�
���7K�X=v}��P	�?l��v�l��k0xO�n�����Wㆰ�v    IEND�B`�PK   ��X��&¿ � /   images/c209dbaa-bae3-4d96-a84f-55b6458b16bc.jpg��wP�Q�/��b�
�(��"]��N����6z3T	Uz��CX(RRB���f����{ggvv��ݻsg�x2��s�gN�O9��<9�8���R�TPQ T?�s<��
��˗�����z��5Z��44��n2�1rܺs��;�}!N.�{l���"b�8�R�De�D�D�����U��W��0����ο�ROSO_��\`���@u�A���7RS�g�o����Kԗ�\�FC{p�����.RS_���'�o�5�}񧗙_^��`�x�|����h�7��+�w�hXo�����_@PHJZF��#9eU5uM-cS3�ss;{G'g������@����Q�1I�)�i�2��E�%�e�5�u��M�-�ttvu���ō�OLN�/,.�WV��wv����)GT��T�{�?�a���¥K/]��<T������}�ˌO���`�x{���3��5���o�W�C4�<R�;��?��z�ߕ���yΧ �/R�=a ��#�������?����?����?����?����?����?����?���`6T��UF1&��"�a�s#���l��I�jl26�;��I�Bk����H�%����r(�.���i)�@���'�l�S����H]8�L�c(�'Q����\]١y������G��9�2�;��vM�[@҄�#qP�N�Qғ��i����y���K���݅�����j�����G,e�W1J�u CU��k�7\���4��I������7�P��ו��P��[��x;�E$��:�Vɧ��VVF$��������?-��*{�]8���@w~$�[�D���,]��(F��)��O؝ՍQUrLW�;�l�S?�;��ha������������ڍ�����J`��!�b����.N=�c��������y^���.��l�� ?���E�b�S����}�� ���iP�V��=�4��w�XՏ
ek��N�����w���BB.��˕f���N���e�Z�n	�I]ɳ[-�`nΣ�O��8���].f���7��i�����֙�i�?�x<�����L�%�-�=3O��.vsu8����m_,fD3M��T�,��QI3ݟs�rΏ������zM��5��Y�'1�M���H��v�o,˸�a��,F�cƶ�y�̗�fj=����#����3&N{��>ڱ�+:�N�;c�1U��/������?��k��t�,w��J5I޴X�WgT�	��|uh]_�1�C�T�����>k��3|Ik�S��:��^��L���~[h�u����>��*���@ø�ݸ)M�n�.s�ȕI����\[4d�*!�C��a�1�0�m�;�Z-�:K�; ͝�����N�������>a������3�<�_Z�ZbQl�h��𨨲
d�0
�06�f����R�X
����&\�VUeаGN�9IŖi��ܪމ��P!�4]�|��ũ��Q�}���?p�\�a�RĤn.�h���X�Y�'�P�g��Jk��s��v8.Jp��]��^P���T2�f���l6���X����7�M\b�?v�TąL]�}48,X��~���Mb��X���;�uz�������:-{xL���`ϖ�O:j�0K8�;w������z�V��Tu�i{v?˓��U0V�/�����j�J�v78���0��:���.zQ~���l9XW����V��ƻ4)�n�q����� #i�i��d�?>��7�~\S�=5���`�ݻ{V�t`TIV�n�\l�8u�j|�|Ε�k���~�Hc��n!��f�d�N�7�XD���iwQ�.��`�����u�Fʾ��?�����2�[j\�f��m�T���^�r��W�(b��ے�Lr_֭ؗ*p؋ �Rps�m��\Eeg�� 4��sl�F�L[j2U�7��z��d+��t��#��?vvF�<QS�fǶ)`_����A�_[���+��U6�o�މS�mh�U�k@��@�$vr�u��0}%�|X]��)�I>����󰽫�s>d�2�8n�q'��/�6I�]�$���zH����K�nW/~!���}��"�0��U�#��xM��������e_���g#����H�e>/W�'Z�u%�3NY�
�n�Ry=��S�03�0;�狸_Tj.E_/!O�9t�-,�g��n��������ƀ�ǂ�?��	�9Na~����,a�V{�La+�/�+������m�D*��/��&�,8Yjv������v��-+���,C�;]9�P�VD-��GZ��p�/�r����x��^���l1�jm7��}<宐��K��?���nwBY�j�mUX��"���Ӥ�!�i��&���d}����O��f�u�����
�Xt�}�T����N���A��$˒K��7�(S���`����� H+�ژ�t�J��6���e4cb<Q����_���Z"HP 9?/��K�)��8�F�p�����7b{��V���2���sG�^�B����T� �4X7�u� Lh'���W�,m���}r�"��_?���#Bm�b�d�zSš�·�@��S77��|�O�ѵ1��F3a�V���_CĨ'�|��L�LS�]�%V��m��Z���n&���U
�9�4j<^u�)���{���ΖyZ[ʅeQ�֧r�����`���������>���,0�@m���g�?�5V6g,��Z�����j�ǙH�<���{z�r�۰OHo{�d��M5�w�O��XQ
�c�a���/�~ސ#Z��<\^op-�l�p[�!rn�Dypy.�爔PY<3o��ҿ�_��$Z�p4�(���W�s$|gx�1���&>c)�{�doo{�S�V�ag��[���:L_��/�֖%3/����|��ح�EKډ��sO���'�_�;F��!�p��:�~F�ݘH)&�A��+]������� ��9���5��Ҿ7 �YpL���س��$Q~�q'B�gn<��]%�$= IJe�w��b���=�e�PO�6��It #����}��;�����e��ʕBC��j"c�K�4B_�>�A=(o���ǲػ���\���nqN�1��,��j�o�Z��>��n$=p��z+e�DX�[{��r�?s��3���D��n3�����z�"���H����:�N�j�%�i6ʦ���QI�ʯ��N}+
�e��#~̝/�Y\�����3�h���_Oz�6������%]Tq�d�M����5C���k2���[�/)�< �?�Ѓ�	f�Î���wXk_����/p�P2y(^����(�s��*�PĔ�1L
T�����r.�՞�'k.���wΗS����9jd&/�D�BF(Hf�Y�?ԥ��x0�e���.�j��cfF�~}웼�6�S��O��u���Ѱ�����	ݳ�mN�ѣ�)1/�^mζ�?�ᰘ��5s�%�&�!)��e��9`�/��ʲ�A�������01Ha�K��C�g��\�6%����7Y8�EaǢU�·��K׬r��-;�]s���T��swJ�	�eW���r���k�R�	Pc��$�C�+W���qڈ�{vΠ��Y�G��7G�����Ne�AtY�ð�n��� �ʡ���E�p;��~��k�?�(f�4�X��)����Y��f�]�?%�|�ONۿo@�ҫ�'5���^���3�|�1��Kp	l(e��󞭨�Ww`u��O$u2&�Wx�v�������m���:��Us�V���(>�3 �����\�j O�G�k��K��죵�M|��3�����`,H��}� E�VPx�%�;��	�)��5��6����l{���">�� �+>�w�,2։�ۍ\3U�����b4�=Ve��0��+�~ub��`&��sc��K�z������_�����Ǫ#_56^�=�x�*o��D�j^����QUGu�.�A��L�w_G#Zb���6�3� �;��8,ݹd}��0���me�m�/����&U,�,?��0f6�wY��q��do�׿��� )�CY�u���w����-���u0:��$�*^� ��~�˰#����g����`�A�{�~E��'����\�"�A�I?�Ѿ������D7�B�Z�����t�:T���}��[��/-�H	��Ċ �?,$�VW�GcMF_�"�D��~��9S�	.?O�+��L+��\X�g�9���FR��+�0� �����$�����ο�ju�J/X}l���(VX�0[�[! ��S��.c�d8�[fkJL��tl(�۪{M"g�J�����okaa�{��?�}v Ђ��~��k>>el�'��ǳO�D��b��ʘ4�c�R�b=�f�|�M�&�w���<a��Ӭ�y�X�2��
P\���;`�F��p�����	s�3��Q3�{`�M�\�a�Q]C�$�{�b����������v����2�CRe��B������o������q�L���x�a�i˘X�_�@J|'�Jo��x�Lg��]��.ut==�y�	P�{��_�-�}�pJ,V]}���k=Q��)��c�}���q!�0��j����XRx��%Ҡ1K�L`Y5p�c�n�WN�M������x7����m��Q��>�[�o;��9�3�e!�t�?��TCʡ���a1�~�W�v��iϘ�/���s�&W��\���F���'`��ni�:`,�z�0�r#ڝ�����Dd�C�Dl�l|�^�zĚR�8CVC�f��Y�ٶ+�O)-}�����h\�a�����B�,u���Y1òG��m��#��̘;�Wȏ'��r$`�n���g�/��ϥ��o�<1ˇ�{�c�8	�tc� �48gEc�`  Bbs�|;ԢяI�]�������ds�����=���%WFu����#�Tՠ3f������
?���Q�fF=3���E���id:��L�D48��d����#4eU~n�SO�/<~��'��5��	��'q|kl׫�.�/\�;�n�G+]����el��^{w���4}q\�O}hrf���Q�؛k��j�����x�$�s ���jW%Qf��E���W������9@���mltO1��]�ݲS�Y��&���چQmS��a���ɩ����rʄ�>`��ɲd-o8��	�x�=b+(d9p�A��8"O��y#zY�xv{I��yCn�n���8�.Ξf�#w�l0Ҧ�t�ū���E�D�|7��u&o�J�,��t���w��Fߗ	�#��db:��w�:�y�v������fN���}ӹ�J�,�_RϦ���)nF���ܥB�k��3IVWwC]�����oZ�|���� i&i'��2�r��7�A'C�ۂ�6矄�����0lvy�*�94=@+���,���'+��5ǿH�Z�xU0�e�M)<.~�%�w�P�V���XI�0{��[ݬ�}"T�c�|2t�����ʔr"�6q5���٨�=���{e�DN�-��A�+�����-�V�̣�c�]+|�yQ<�嚑JU3;����1ɝ�9A�u�T�����7��\�ULlS�Ӫ' �L�����#�x^�J�HH�;�>~e�̌3��;Wo��;j���(j�/}��.	?�\�hQ�$[&z�S�9��<�*�jVa�"�c{�3՗Gb�Y�G��tz��×��8%�6<��>��;A(o�ј�����ZWk-SW�	�A���E���D�G3���)�x�B
���q�ّ�*I�fIУ����Z��yӥGHۄ�y�f��_�c������.��6��y(�-���E��X����س.
ޤZ�_�
����"��g�c�D�YMl8<�H��~u�x���]�-_ �s�i���_�@�>Ɲ�<$yE��Z������;ûC}�U��xZRް���<�Yνy�}�ɸ�z�)�eNok�ֺ�/�!�$����|��p@�M��;�e���\�{і:-���z�}X��ҔhToRe�w�(�� TV�*�^kD��yO�8J�!]��ٰ�p�G��P�������iPO���#�Â��\��� �Cv�r��T����& 
-_��V!��KE41K����~]��}���'��$x4i�[�t�y��g��!�&,�!�U�t"�,b�=��S�m�Q�
�)��KwG��1h	��	��b�.��b��c�l�c���4��g@;��<կg"bS�,vcz���+�uv����8�X.� lj�/�;�woP�	���y�-���g.����L��Zx4��y�ϺBg䲠�j>��FK��V[E8���h�Ϗ��$Y���~ڄ��|w��� ���x�j��ȇJ�*����F9l!3Z��kV@�d������i<��k�L�[�C=��%g&�� w[Я����`]���
� �҆j�_Ly�ifoV!R�(�c>U[��[hv� "A~���zًA:;��gk����*W!��|a�&sNׇߐI�_�������/�U��[8b��qY�쥺��c�[���A��X������?�z���%xph�"2Q9s�w�>�rZ�����W�6T����R�Or�ؔ������t�z��l��,���y�p�n(�e�o��������
�Y<֘H��������T�8-�cU'6}s�,� U��[1+ǣ�zl	S��'�@d���Z�~��������_)��������F`/m��ќu@�f*�^�EJ7�'�J�s������0�K�]q�[.hM��Zd]�V7�����G�@8��>����T��V�a�����yʹo�����宥�"���叾nO�P���b��>�Um�"���7'��n��b�Om�c47�M�oLk�͞����V*:��[ĭ��_�V�]����hW����oe��ں?TGN�6��g\#�閙�Xҋq�@�[(�[�>�G��2�ѱ���Zu��yy�7IXE,~��#yT�I��1�l���2�����!�7�GW��1�d�wJ�/p�\1b��wUb��j}��-��\�� N�"d6�H�x�X�h�#��D�Ů[���O>v�T}�8f��E�����["�?�-f'�67p���Qȗ�bi��W��o�hd��|T0k~s���u�d�6��T�@��3e����P�d��/�u�h.o)׈  ̄��=����씭�F8��Y)�^�^�hB�!����!�YB� ���z<޷�����P�� ٓK�R��Pw��yj�����#�+���7��ݬ�~��A�Tm�6�@�{q�|�x4�ݓ�v���oD��,�$&��t�IrC�w��h�����}/^:�0F&��B>�J�s�qu�,r��t���}����h�w���p)�Y��V]�u�f8���i��kN�l-�����S�m����� !�n�)�j�g[t��s@�������%�����ƗrW{�(�7��#��ڇ�3ՙ��6���ۋۿ�+b�%`a�DӴ�啱�s�(W�#�Ukt�v�gB�����;J�,+~���p:���s7�-�L�r���Kn�7�)�[{ 6�*���I�}�<x����תe��c���J�ж �J�0�d�����<�YF�$�����pX�C�0���F<�DĦq�#���F{�T�u��!$'�=1�u����Å�/M9�ˏ��#��RϘ��=c���R9;�OVh�ݡ�:��%� ۽A��D-Qfu:x�B;�.[��/i��R����v�%����L+y~�<,Q!�,$��'e�w[��|�b&˵����:c�8ԏҼR[tJ�7m����I��6���icR����?������hx��&�ϼ��'��$��n��:�7{�ts���M�<-����g,��Ba����{9�+tF;'\�ŷm����I� Na;�/���59�(��i��Y�[� 6ٲ273Aq��%�O��	b�"
֑%�$� �����Ҡ(��Y��jš��d?�gB�_@oHR}�p�dе��`VR��+30d
�U����Ƣ$\�i�4U���=�_��;�J�����ȇn8��bbO��5�,�mbZ�?���V�?�<�t��8�9o��-��	�m��D`�c�/�+H�t��0����<��/Ǝ�j��_*���9?*��CۓK��H�q�Z2a՛��+�;>�������~%BfJ噴�r���5g"<����d,��.�yb�V���jG�5���M�����cḏ�gUA`�<(ģھy�_�d,tf����*��H��U��u��̨�u^��W������ �M��-Oѝ�։ɺqUS瀢��������ꇿvX'J��k8�%����ǽ�H��)W�I������\��Px�1t��k�u�b5j`�� ��t��]�D����!�W6~ń����S��zjF� �B�'ȭ���B�"=~�/A�5�o�Xv�y΃�[f���J�z�.�.r7������p�z���C�Z�q���o�����[�A��E�����k��(s�R)ͤA���⳿�G>]�ſÉ������t7Ю���[��¾;�tū?�"�7�����Q�IW�	�ҺY�Mn�gɺ'�c�zYnǋ�խ�˂�bS��n\�(tT��4q3b]��HV �:Y�k`�4��s,[Ȱ��@r����5O�Է�!�����򗃻i�55�|�/�z�T�nbE}N�#Gx�컌d�[�󚘊D�4"3�kr�rK�@4�{����K�z9� 	���/���S�nMX�Ac�(��K��~��r'���沎-x���t�V��J���f�cF�Rp���K���hb/��������1�>���Y��iJ���c/#��Ki��D��g:��H��i���*ۄ��Wl���,�**8��K1N����t��Y�d=�km�D��V�|&f\n�h.��[�9y樸�>��*�j� �#��k��v�g���д�BGȜ+��%Vh��:d2�V�C�o r>�Cj�	0�gN����z@�x�jJs��V,VLZSƇCJ#����V w~���'�a��SE����eL�$�؋++U�3Lᾮ7��>�8�#��@���u�,���}.p<G��Pİ�|���f��l#{]��:������R�)z�%
�1V��w�<NE�^�iˌd�v>�N���9���c�:�+�YoM��	�J7���U���u�<n�h�p������d�������H�F���OW#H��Wq��YR۽o�A�I_�gP9�6��V����@X��﷐�g����5R���h�˫��V�P�Jm�d.�!%�S"R@l=ʊ+���0EhT����h'J^����"$H�x�fM��<GEbmF�GT�>�Յ�˕ֲ@:S��t�K���JD���}�'#��Aqa�أt˻��FX�]�5.wU=ۦ.c*4������q�t��
]UG�'���ϲ6q7%.f����"�(���컛�cfg|�[D��^�n3�F�K�H��O��p��B�`�:�~^}ҥ�ca��
w��1"l����&���׍���P���ճ��xQTV�����P���:S��bu7?�"�7���LK*��MM�&�̶��+F�`��o������#>e�����K��_�Z����P�=a�I�4�g �O�P0��y<�S��z;�e���+�"���N�-�.���Z�e�&�˛L� �����k�=���]~㞶��Z���s~�)*h~���1,i��ھK�0 ��y�7_r�uߟL���;0Ca�WmoGF���;�.�̪B\տ��bt����`O��7,*
�/.R�n���;�U�Y����W���Y�ȯ�D-ú	����5�n��
����=�m����1����N���r��q��5��!5��;o፦�z��a�J����Ğ�R�1����	��e@��U1���f��	t�@.����G���)��>Bo���|*����?SZ�o��%�l��!�~]�:K����6b�FF��ksP�)�rK'�1�gr�����pf��8Q���~�1w:ox](oO�(0б�6��Ћ ��;�`k��
Μ�S�MP��TL(:�؁���Kڰ]�ɏ'm?�_}Gv�/�(S7YoE�����>d?������m	��f�2W2�B�70�l���k~�O�n�S�m�p��('B�yR8+j��p���(�&�;eʶ��x]�o�
Q�z���v1;�kT�z�L�(Ґ���k�̓����[�gݦǃ�^E$8��&o6N�]�s������22,�*I_�5���A�Z�T���A��MH�B���g$Bm=+���=�5�{4Y?.��0��e��J�����5����[w�R��QZ%B���S��53�F��ԧ�#�Cӝ���̧��[���7��U�O���I�����9��Ms�J�vA��^n�d?�k�*Ƚ-J���ڏ��T<��'�߹�g�٤��^/%Y�tr�o�hM�m���8f���Z��'{��Me<�ß�_Z�ހ����	������dH\�'e�����L �Хz�����P�ہm �2Z$9в�'z��1X�ϧ:5�VZ���d"i���1�U��h;������k*+>��oO瞔�<�~�jX�������b����+�LE�'=o�Mz�wu�Q3���cYq۷�_� ��4�:n�s
{=��4�'c[��j�r`�[��o�4����hFYB����?b朰	
qOT_�y�.ӷ*1���n�ˈ�?���U�C��@�ť*x>��׳�:ا�ͮ�T�r�x�L����~��t3,}�}*8���v����R(�\a�q�}����rs�����-*VI�-�+���-t��H觎p��/�u�5�-�#�&���%���Ǻ?��%vA�n�w��i��O���Z��4�j�ү��j8��t�����W��p�q�9��ˬ�r�W�kI�ڒ"^��ؚ^���6�'��DGt�k9��y��O�^U�����E]��!��#`���ٞt�\,���I�׷�(�~9La�0�m�q���ܫ&SG/�?ք)�'g�9r� +{B���p��Ȃ�y����z����y�k����u�y\��R|l��j�H7�w���4�dN�y���W+h�����B�в�{���GNnN/�c@��30����'d��Q����E��L�=�'e� f��;�9��b���J֮�q� � �u�k&����E�q2lE�-i��	eѶT�{[���׫S�-��^�b��v~V��ꍯB8w�ɒ?.�ǣ��
�}��L?i�A�sA�2�><�z���
��&��������u��]EQUa������+[!���C��_�1�~	���4Ⱥ-W�+���&/SlI���ǅ�8�֑ ��X�������t��~�,
U�������h���y`�;鱵�;?�ItV];]�*2�ժ/n��L�p�3l%�=�����yC���^��}�Y�ڝ�ŤwK~�B�9H���?l0�YV�Tmm�?�B#ϛΆ�\�1��,26X�������iV�����J���M<���+C�m�G�{8���yd�f����#G�q�pm��E�GZhC�(��[���f%���:�D�\Ө_���d�/��Ktǘ�~Xx�3I� ����[l�:� 1}z�Z�9��.�
"H]�����ٹ>��K-Y�eb���Y�&�'���eR{b���ެt �����)tɖJ�T��?+xd���Џ~���ؼ9R^��e
7����\#��SO�&��a	2�P^`Vr�rC�"����-�(t;hf���ddk���
Li��r��n�3kK�rhk���,b�]��5v�
�]�<N����i�h]����B�Q<��Ǟ�C����ӵj="����`��g^[+l�@�!"`c�JuN�b�;g}S7�xnv��4�I�i�3iX���}T=�Q͢U����>$��>&��9�������b�`u�7��:�y�6�)6q��F���"�&������xT�ʊ��z�P�W�������7"U��D����[4R�Tz�����~�o�=����Ъވ�QY�c�v�#��h��(����t�v�%
����uO_�Z-������JL�z=�S`���(�t���qV� �"��Su�h�I�>{���:�fo�*��k��X&I;����b��$z��;��lj��/G��X�q0�ĳ_x���w4jN]Gѧ\���p�P���n�|�'���l#�@����X·��⣄�D��m%r<#Z�s��72KW%z���W�8����!uF�:����8]Z+F�W.�řq��|��+2� �F��/u/�ב8����ҮP��Ous�RF垊 �v���S��4�޹d�ՑaTC.l%�����e���X�Խ��z��/`jd�DM��c9���B��*u]ڙ���7�DWV����{��C(Т���/I�$ᵫ�a��q�߽�02߈�h[&���rubMp�m���7�ar�7����#?LV�����.^'(ݐ��������c��� � sj`��ED4�Q�{��d�>��2�6ΖL��d�)�������
�L�UU^�5��_�G����;�]*:�.���z�l5��$J�B�� �ճ�a�-F2���Kmt�l��%o�g��j��-�I�1f��H�q�0tK� T�-�g��g�$��������C@v�Ȁ���߉�,>pa��h�u1����]�p�e�߳λ֘Gi�{�olU
�qQ�}�(�-� �푗?�8ѹ�lFѥ���j���a��B��ύn�䲢�m&�,�H
�\kZ�����wcD/�e�n���zx���jj1�/��{t1Q��ʯ�,��˾���7բ���{������k��%;a�q�Mo3H*P�ï
��R���Sho��XܘH�~(3-�l��4Cm߬ �zphLr���_K���Y�to3֝��L�弯�^<D����
���k)��))����8>r��DE)1;Vت���_-�Z}I�A.),�'����	]�¶�6q�� 46�P]�cL�����z4w{?�O��ޡ�d�S�3Қ@����L	å)��̉�~�k�O�}D>b��O�杈���&.�"t��8��kpgk���A�婀�L�Ი2��,��gA�۾�ZIW��&���ܥ���L��o��.�Za݆�.�@�>7�93�[�Zٛ�7����H�}q{���ygܘ�m��n.e�����~o����B�{����)����"�f��R�8BY�������RR�],̶�����b�j���-H1&���d?��QƐ�k�9k�L�E�ؾ��	}�!G��}����s�j�0�}��a����+g�B�?�Vob^�w���5T
`�ֿ�F��_\�ϣm�������
W�]#7Q�]G��!��"~�WCS ���݄x�;�2���cg���R���(Yw�F��>g�]<i���z�!�})DH��d�:�Fv���h3WpW�2��ٿz�$v�@K�k��[�Pg[�<kߕO��?��ئ�k���"psh �/Mkܼ]��5Q�CǶ��A�Y���q],��]u&M�3'�T:4��f��t�k���W�{�Iz ����	���z,�?nke�_��cdJf(F�e�VҴY��ɛײ�����ݲ�>Fԝ�a�Q�ǥ���#�y�$�|����j�ַ��vo� z��4�g��1|��ު	�iܥ�	,o}����.���mvs�2:�]2�[�ع�94��,��7�lA�o��nwm��n3�cI�$���z.Q8�:45̏1 ����w��5N�v��! rKD�'<��a���ufƼچu�*��.�f�h]bzN���"Yw��>?��~{�e]M�o��ah�X&����ˡ���BO�q=�4:i�籚���z)���fz{��	V\N�E�^�G�*�f&;�wp�ٰ�b��{ǚ���e0�AB����0���;�.�^�\]�+�E.PYU'���E�pQ�s���U�9mI,�������9%�y��@�]
��_=����'G�f��v�d�R��.P7��L���� Y�#m�uz���4W҆��5��3l�mn���ղ�����4[��7M�g�j-ȤQe�����],��qo�����#m0��{�����&(c�RR��u��[}��u�U�]�/P��8,�SW��+��7�]�r4Q�dXh}{ۘ��'*Zi���ۧx�+]84����$*�ح;gXbj����6^?J�񔼐�
�A�\�} �ϥ���V�M ��wbH��D�U?���sT���Q�)_v�$fҤ;m+@�o�WOd��@� ;���m��&����&�XVZ�=�W�?L�~=g�_�>�a�n2����ё�K�z�7���d���GA֤��'VhC1VU��^��%/𻥮=���; �M���+�1��c�;���5#K���(�?=�n�Ï�.���O��і���a	Ҕ�y�4|���X���o��?���XH�n�Sׇ���ZC,�E�N���үģbM헵���N"9�ҍ��|�Sf/=˝��BQ���/����p����8`{��4�/lGeVo�|-�ⲳ��ň��a<�B�|�|���v3�1����� ���q�ޮ)�V���O]����n��hs߰�1����W>��a����h!ˏ-��r����i�Jr�n��$�c��a���oK�џ��a5!���-�k�)(�U�w�7�� ���!
�~jz�!��X���&}�R ���W���f�wl�g((-b��}G�6{��kY�
��r�p�P�=��8N��M��<�%�R	�� M}2(n�)d�-���|綥4 }%�S��ǭ�Ưgg-ϱC�F=݄2�)�����Lb޳2���+tgX�"�YZ�ל�֛���O�t`�m���t�@OA�Ⴃ�z��\S+)���U{��!O�L]�U繢�-~��=��z[��q�l�������'4i-�:�L���U�,b�֗W���o�͜MXB��3N�>�Y��zz����,�!��-G�;�wR"�nB��m�7���2��UY޴���X����F[j�!Zf���V1����yk'=O{s�3��fe?��[�3[И�_z�(�?�.�>F1�&��\��MQ�F�$*�v�E̿X����qQ���j�f���j��̀�_����I9�����c�f���Oޙ:�������X��kp7��l��xo>�k�������lWͫFpS�����%�Β[ط>��uG-���6q���˜e�"aca-.l��Uj�m��N�C �2Ŏ^��ne�����<��e&��%��MZ� ����e�+��Bu�U�]�ǿ�5e�s�O��j�e��D�}��DF���Fۗ^L0W\��uk�g&�o��(aǣ�!'m)7��@�ϗ�fO��rN�.ȇ�"]�>xHU��)�\Rgf�%?����3��ƃ9C�v���ŧ�5c�-��&[3}�v���۷�i�:0&�7����te�5�MO�)%i��B�^����(J"�J@g�?c*�Vq���ǳ>{uU -�k1���n���.�t^+G�����|�Kl&��5����iUY��$��8�2�5r������=�=��L^���yo�g��[��t�}fr�t�y�H9x��Dm%,wZ��H:��E4���j������]nmߜ���;���`��ۉ�]|Z��Dy�'C��h`�*Ƨ"���0>�o�{���(��t�l������z��4~,9 q�zBg�� ,@?��c>W���˧j�Q�(ݿs�#�	]\UN��f�k1���d������wIũL�9�q��kHc���D�2'��F[��o�i�ӽ=Cw1�� �g2�t�=l���V��zI�5�J���U��Bj��Zl���<Q������$��ڭ�&d����]$�Y|d��i9����{O��|���h3n�[��mD�XL�?�ήb��K[ܹ��\����f�62I�
tFEcVX*W��)��)�]���#{�ț�_)�H�V���:��=�<��'ʺ����J�s�w�C(|[j��QH�P@���ƑS=#�T�LͅJѢ��ewR��������A�n�lo����N��Go�������^0�W��z�M�j�B��7�&G�Uܪy�:'�~]�����8��i�"0^��fT�'2��C�-�<*�-��oت/�@O�G,`�~i6�f�9�l�X6fi����zӖ��+@=qX�[8���D��HE�.N����tJ����m�m2�C)�4z&i57{,F�_8;�&���OLPDT���F������f0J6F3,���;�$ƀJ�@b�Hw��}}������o�s��\����s]�Y����p	G�L��/f��.�
��fS렇�Z���"vB�4�{?s� ���y��ڦl����|O��MH��9�m�/��u_$��դ~�jz팫}�P�p^�0y��OР��~�4���
KA�/�E=�������1�m��)����ؽ2��D�KShI�,'��!�a��[�gw!�ɽ�a?�&>�^�����!���8�n�Pab!v4�����C�6�j���gh}k�E�1o�8��+���g�nb�h�¦)(��-<��!7$��+�Jed~��|���-���#[l\}�һ$�<�j�,����ծ�w�������>�9|\��^ ><o�H}vPC��ω��Ck�]C�'���-�7����q>�V�AO
\��NR��ݾ��C �5��Ƕf��b���s�w��5�\��4��DDև�]u�i?C�����⪶8�@���ނ?�=|PЃ��*�#�̩خ&��1lѽ�}�9��YXi�.m�$R|Ү�}��C\m��s���sjO�BT��=A$3�
(�ǶDo���v6���}�ي	��P���s�޷i�Ƹ$(���9��um����]*�m��7~8C���Q���$X
~^����a��J�1���é�+��=s]>v/��T�����vT�Tǵ�����d�ʐ��e�*&�'5K����{n�y�L���-o��'It3!��Զ4;.?��U���%���k��I�4�.�O�ѭ������k�>O��r�\Z=2?�0�t����H� ��b�jJ	�zOkG�!�o�w2
�M��:��+��Qw��k�+�c)����;�׼�o8��vL^��
� �ߓ\��>/� �R���)�'�R�4�UI��K�,cΨ��
�*�1_�{��`X7�.�
yl��]���s�?(����W�s	���������	��o�3���^�
�	V|��2q�O�f#L�9U�|���YjTkY#�;Y�#X�)Is��!��VT�i�D�_0���ә�C:�g�$��3�r���<7�?`��35�Q9|X���Y�p��卡�i{��&���)#e��G�[$>��a����,�`��i���>�~���X�
06���n3 �$�c��^K-�T4lP���>p!����,��:8V�N'��y�{�Y�� 7���팛����Od�"R +��IN0�ȭ�%2����^�S��WٷW����Z�l�|���i�Ϣݻ�����Qn��J2|d=��V�&�RD��N?�#4���r�Wc��($���%�	�s���<��y�z����bK)�-[�K� ��V�7P��M�OY��>��zjn����&تܽӨ���x��<[����9l�T�$�ԛ'�rb	���h��ZcI�b���:�}��������)&�	L��������v�)L�>\U�Ȑb�����E�]XA�-���<3��ÇK�f g�6�(�Ȏ���T\�J��B=�X�!��Q2
�.��_*�^��s�}\y�a��#"�E�5��� �P��O��Z�� ��V�Ѧ鞎36Eh�)׬xwW�udbY_I�`F���sJ�@Ն^�py>�>�<(�>�r�gќy�(h!�+Mk4,�i�=��s����V�q>�c��nâj�v�S���c���,񡫚G'%����2��oE�m%sO"#�_¦�0oT���;��uC%�J>��N��f�WOT"��<���i����RJQ\�M"f�\��+�v>:�"q�W�;5�*��em�o&D�{�y��L�`Ɵ�/���i2�����ٻ���j��J)-.��N�פ{�t�N"�,i�^3x��$�:���o��gf�!�/[Dv���>� �\{T����fu樨S|�E2�V�?&�lu�v�'�|���&���{+�Nn<'4�
u-F6����L
�88d��ʥ|fL��f��|M�zI,R:�e6羏�O+�Ve������T��?��dT'��W���-�|q��Y�j��,h���EQ/K����CA�O��,��f�A?l#��f���f{=�5зq�(D�G�|\O��6@*)]X�ɓ���1�3ykJ������!�O/��Y���'���گm%���UP�����V��:Q[V���,�!S5i3�C�O/����ZD��$���FM�����$�<�i�U@�S{A��7;��\�¢8�t������!R(��z��t������N���W�?{X{$�e�f���v͞�4�1h)ў�Y!����%�W��lLA^V�ҋz�\\F;�<I�o1[`Qӿ�d��4�@���v���ȝe.��4�m�=��?M��t�6֏Xx���D�[��Q��|x�+�˗a���hf��E�8G���X�s�
G��s��(S ��g� �U�� ���{�4Ѧ��Gu=�R*d��EͿ>/��,�����ڞ���W2i�+��J]�1��{�����`Z���K���q���#,��"G��B�X����f�9�&���iH����R:��m!��m�'�4N�'�^n,Nae�g!��W���IC~�l�E�����"Ru_����:bD������q,f�: m��M	�jǫ��X5U:��_�|���唓�^�����l��v���Y�\&��%Z��
�u��[�k�t�$Zdl�P5e�^����L����_O�(�|C��q櫿���*O�����=�_Ս<誩;�/��~�o;�<�=cx�$rn������^�ɗ�,H�b�L]U}E_��ݘ�MCo	=vG	9��j���[�-˃����g��n�!
�됡*����-�:��`Tp���5��U0���oǹR���ĩ�WS��J���yg�R�#�֥� �#�c-�
���1:��E.:��G| m�Rk�W�oI���Wy/��㷾����F�lb��f&f���h!<���f�|�2H�ч頏!��l�9�2@����̏/sM�p#+0��~�q����������
��$Yڨ��;H��_np��~�T;#*�S�EN��{
�M�ҡ��U����ˬL(�_��L�&>0�ӚY�f�:A��W��\��4hz�9>f���FDKX��K����}�� �U�U���gK�t�po��N%6L�㷯��(��뫋9��{0�^��W�g�ٶ|W{5k�i�[|K|��i����1��})�ڐdV1�ힴ���m�5|���Z6�S͢�����N���@!}�fX�g%X����{x}����P����+,�>�R$�,ӭ��p#�mQ�@���]��ݶ׵;�7����̥ٶ��'k���_�%K�ԯj��^.#!��9&*��/� ��"�t~MÓV��$���#��̚k�D�5qnR�XS�bXq����<�:�Ф���Ʃ���z}j/��KxC)�Ց�����{�45f����S	Bۉ���5�_�L����>x
z����編o1�����%������k�?s��Ĳhb��Bn�n���L�=���g���Y�'�s�}�#x�J7÷:�[���3>͢w�~>+��mp���"8`�B�z�a��j��ۏԚ;����v���i��Pa=�P�9^�֕�����'x��B���j��ɛ�*`ڑ(;Cf�:Z�>��`��l��Y�.ހ33��X�'��4��kB��NB6._�~�H�1ps��ՙ���-�z�{_z�WN��j'C�6?*Ab�'&X�1�)��-бO�@t�W��4S�����FB�L����Bp��z��YS٠�N�at�W-�M�g�S�`Jb<S�c0~��$��%k3���BIV���{������������Z\�mƷ�h�e���6���!Ĳ���~�2�uO�a��ˮ��/k�]� H�$Q׶��V<�ՉQ��.�>+�-���d�e�kK�����u�L��^�1*��3��it�7�Sj�����c~��~�nщť��5Y����Ht����[l���A&w����N�oOH���]���rE�e�=n��!����k�b��:�Qu�S2"���M�aD|�CD�3�i�|o�}d$	rYdþ�N�#-s,egn$S5�vAJcQ���9U�a~���{����3R���J��Þ����o���k �Ϛ�'�yq�5@�#=�6��>9,?�$�1�Z�xW�^u�o�F>u�ur�N��;��%��mP���T�z�S�{;3?�]11/}�]��2h�<V�\kP��9e�6fj(�����	*q_���L�F�e��	���Wge9��\�Xz�dw+��2��V�*V�HF@�NINqD(Ҏz٠��t�:�mb���5�FG[v��i�G~����JX�/Z��]�a��x�][e9/���@'��ZX�EXʓ��v �Ԫ����NCH��J m����6!̻s�~! ����c0I_���/8T-��E6-y��[ff&�룦��l���	"*�*.{rR�
��!�\�~H��Gn�PK�_pdI/.�K�uA�\4�+�j�<f�{�7��
�u��M�Q��5������Ȕ�m�P��!U,C�$"������~Y������i��j�e�F�*$Z�;W
B5�� �d�/�1��Y��1�)D�2-��/���Pw�����Γ�.2r0��Iq�(C�T��|�7��r��+����7h�:�ڲD���QhCֶ���5���i=U#� ����Y�ə��2�&[��r�~�W��	Z�4���۹�	�7c6f5�vϕ�m���_.Ngaɏ���8	�#�i�-}��~1b�:���]4�7�����[��<x�r+�â!�=A��&��_�y�]�
?b'��K8�F�)?�]~��rt]|�ָ�>0�v��M�o=a{X%�ٝEF����m���aÚ|��s1qt�ۉbFw^M��`h�6��{20�Y��=q���yv�_�Am���n-�I���jO��/Nv%6d�T#�%��w%�i0J����/���8K��l`�DX
 ���JCǤ��u��Y�[h�*�a�M�,j�@��g���x]�k��ą8I5c��������K[���1��!��*P�I�S�[���4�Ub���z�;�c�t��p=��j�cr������D��#�.f1(���t:�Bm�rst�?�����]��`6��T��� ����6�6Kͷ˵"g�m�WfJ�({�g�^���I��x�����2��a��y��ˍS|��ɤ��?�I�g#���X4]ۻe?b��D6;�����2�s�1����S���3w
̷��XS+�C�Ф��_��ƥ-�	s_�+ȉ$������=/����^�Zdp}�l������:qJ���xP�]��,�ۯV���=���,�a�,�#HS��(h�x��$�Љy����P�2f5��q�������:~>N}��r��y/��Q寞����$�l�:V�.��l��%�3
p=���M\mp(��P�>����Y?"��*݄�*�X���珫`��Yd��:+(��.��m��ɾrk�](D"�b#��{gOzpN�?bW��ފ��`�6q`��-
�Q��(���t����5�m�`� ���ū��loѩW J�����t-���='t(����!ifjX�_�8rG�|���Mή�o��pHl4vg'7��
�u�4Jh�u\fw��՞D��{�j)/�xW��[#1��+���N���Qǈo8���������/�ă��y��/��j�9��xx�N�����fZS�H��"��V�|�%��+0s�Y����Αɷ����I|�(�8=+�c�z$m&�R涪�3_��u��Q����a$dׁ��Y�P�U������a
Qj-�h��}�� Sz�k���{-~����{=-���z ������@�/C�Oq㹫���Ѓ�k�Q�9qMR���x�T�3�=g 6��?��11*f�X$�eǟ�$��y��ѵ����S�=j�-���pZ��HR6M���3v��V����Q�����k�:�� �{=A�/���;T�47�P����*���򐭱_�n�d���� ��Ƅ��;fƠ�KZ!��aI��0�Bd Osnʳ��`��Ik]z���#�����L�N��!琤���Z��� %(�(����� %�Ÿ����e ��b�M�muWc��`ba���)��<=¹t4ڎNe�"�Q��n�>F��DD�E8�+xߎ���zڳfb1�[ݽP���z'!����Y�p�;9�U,�m~�R*:�b�>4m����Q�v?�s�5��*6���T-ɢ�Ee���et*�u��4r�x ��\�'�[���܍ �=O:Ɂ�L��IU�bH�6\�)S�T�58�ּ�Y�P57� �����z�?2��r��	�����bA5�_M5�:`��q
�W !~fM�X�n�Lg�9�^�s�N?0�Y�
���kp5)Z�5f����WS��n�di>��*�}~6�E�#HJ�azַK�Y���K��3�Ť�t�M�r��ƟB�v��D���Y��������ɟ�Ҩ���x����>(��a�r��+�-�Va����W�F�=��N[��~��6���3��"��q.�}L��?`:��:�^M\��W/�Uc1:�!����IG���5�͐x�,�ª��)�3�;Ʀ�%���j��Kܸ����*�8xr��	03?t����^=��QF=�'�����v���hN"U1�/�B�$"<��B{���~�Q�5.v�s��PZ�o���JV���\�.wg%������T����.'�N;����[�o� `$�w��]#ZQ���tq�1�)ED.�!��*�����J�����ɓb�����T��{�YL�h���ؿ3�uNe�j�-
,�Uj!"�p�Xibx����'�_VB��D�m�i�;gS����y�<���t��䯩���{�4�:�	I�q#����߂9�z�P��F$�Qې�d���
K�Ug̿����*�R��ݻǍ��cϻ��o�2S��Ҭm��\�f�B;گ����<����~�b]�b�f[u}˨TZ_�T���pMA
�D��p�/\��d�zh��.T|]"�����A2�x��zK7�/�Xv ��>���(9�Ug
�G,A+��>��v`ݖ0�=f�ɑ��-�&�wYY`.�=ΐM���V1"��3�Ru�DѸ��0��i7��]��RE�Dv�����<��r�W���BK�gME$����&^���H]�;t��s
�li�� �f#	jB����%D�M��۴;�2��1��wN[ ����0ep�':{ø3q7��,�TU:3�7TK7��-WO�!�ٮ]���DW����Q���1ÍsH�/����`�Z�%7�����b)B��Uz���އ���o7� ������t�x$��̆���E����>Y���ʹ�e�.����s<�GQǬ3o*���*�Ĳ�_�u�ۡ~w"���[��qw��V���������5g�Dn>�|������0<`'�s���Z�>�7����j�����M��e����..M΢����K��=�ք�{fī]��~鄕R�����~�aVFu��E�����K�Y)��1���_�{$�;�=	��?��|mT6����9�����4�9��m���5��5y��/q�E��ꝚH�+ �W�ɬ��bwHv���|[��Zm�u��#� Y�zm�|������q��s��\m��׋�ؗ����koHue���m����oGר�K�>�/���0�XL��_�R�	$�T5'A�x]����5wG1GHX�I���/T�L/r�3��1L�{�Գ܅q�[D�>4��}%%q�а8~倇�ϣ��n)mV��Q5�)���膮��kt�i�ڇ="�>a�� �b��GF�?gH����4k��S�<Bq��W�e�����Mb;5�V*�Sk����_cٯ z�.�����z��Krⷦ7��
n��<�8M�����nK�2M�����.U+7�j�m������Q
ߢio��U�=U�LS9���x��7�Y<`��",6�	ꉷ�-pe�Lx(������	[�����@��?�L�*�3#е;n�4����z7��uX^l��>�?x���x=�a�x���0����&}���3yܵ���%|la�{�j2ň����:��&Ow�yURz��:����Ƞ��Ӿ�p���z@�Iꢱ�.�bw���>�������ͭ>�.G`�V�f��4ٕMa�mG'�^��ɏm���ei���O�J����/"�����s���k�
g�ƾ�E��MX��X�Ջ�#[�t�������4��5I�buV�!+�7����8)WD�cj�w(T<��j��S�j�w���r���}7C���_�x�|��E>���m�G��:��DI�S�ߤ��h����Ʌ��N隑�<��
���B�l���<���.���x��[x�K9ץ)����"FP��]�4tAu���I.7f�.m� �C���PV���FX6d�D�P��ָ	"�n����x:Xc$��+l:���%Ҽ�rX��b��F
�B���S3,��!3ڊ�x��~���Xp�P�U�K�Ii�א�ul�@ FXa(������Fn�f�sL�yM��� �QR8}���\V=�����{dK�gzV�}L�#�����nܯF��I˞���x��߫�O�@��n��^�@����$8��E7\+4��'r���6�Q���y�K��C�?|t�����Ww��*P�T��w~dmS֜�a��c՞3�{�Uo0-��.��1�ͱL�i���wc�
���V8��cȹ�f^�>��m�9�i����+'�E�<��2��򕀋��[�ⶃ4����}G���:��ѥ7v�4�u������� ���³�ݖ�J�'h�ӰW�1�Yg��?"�S���=^=C��*zF��9�0���e}���Y��\��B�ۖ��9㪦���s���؃��/��g��i�=1
N�N8'�6˝#��g_���e܄x�aYz��%��� !��?�BPxO��f�b��Ĩ~��[��=���|���zv��]���C�ŵ��wMe}��� �I�׺��K��`�#�Das���ѯ�����AI	\��m��U<�n�a���H+v�	F�g��!a�F<(�����6�i�gÊ�ߎbza�SoM��%kF�i�N�ʂ�4W� �r��ܼ��(\ſ�����S�b�.8��]\g�*f�a	�
�����߀ �E%G�y�����f������b����>���BHl%Jz,�kzI�Cƌ�+@y^����r��SP�	>��h}�}�j�B���@��n�~!)�t��q�a�4`H�؜��E�I]�|�^1��txߊ"�U��=�o��7(�C�X-��Ԫ��������,ED����m�{)����&����w~�*$݇�k�A­Mg6�]�?`
�1(�%S#C�i�&�(ȘD!S��|����a���|�
��s�A8I'�,�k|α5HP�йw8| �L�Z�F��|Խ�v�NX���lwW�D���};�D7,r���@0�Ҽ86��y�4�y;r��{@E5/6]^_�dA�(�fe��&�9�~���[p�y����[z���ueMEw� ��-�v�JӓM����[�	�Z��~l@�[ZP�O9��]����F���6K��M�[�����4@W+�I͍��ۦ5���ڂƈ�˔��d.3���6��G�VMyFť��%��N!"{��	ΥK#�c%�ѩ��WI�P>���Hg�ǀ��=�XLzgߍ-�	t��:<?�U{ڷ�thS�|��%?���5<&W	����Տ���|��𿋥-�1#Rz�g�w*lL���F)�K�;�[��|׹��T��y�λ��:U�C�OA�"�
D��sv�4�2K���湉S=D�8c5��.�o�ҒI���p���Q�� y�\^�r�s�T�9��s�,���IA>�F�iH1��58�f����M��� Q�ڪ�v��u>�(�]Tk�]i#X�_�cӢ[����&a�m,A�RQvU���h�Y��:e�:N�$�+��	k;{jbOq@�[]D��.�޹�+@��m���UΧ�P�WYs�Gt윟����S�h���]�^b`x^m�G���n��p���!��T��Ѡ��`;��.�}��uoZ���]�U ��Н��`���ڇ4ot�%L�;;5��N�5}Eg?Mkv�<}�YLE^^6K2h�&[�ۗᤄG����0�s�(�z���ԣ��~�t�nsM��[X'����#ѓ��Z�U�"��F�������P/N��f�NH�ў�8�uj7��*�ځbo�qv���D�Y	1��!2��� ��Y_�֘�e��K�A�Ȅ��+��S����%�K���%��󎑱q)
Y��gLU�{��]�.�r�����A"{bZn���K�ʴN�u�Y _g@5t�J?i!����ӄ�R�޽q�r_����"0�1	P��Ӆ���8L��:MZ1>����&@1� w;��:��GX�l؊�[]d��]ʊ6y豆�����K�X�jaH!�\7_Z;V~l��aB�wL��XSH�j�(�[yr�HI�[�/{�r��T�Z�Y����o�61m�"���N�����B�$ӿ��؂Z%n��v>Ao �N}6�jwN�}��rFi��^�4ϩj��:�p�/�#:�/I���Ħ��5�IRv/�>�7��:d(m��JF���YH�?5N���6��3 �+�ˉ��\L��@��W֤Z�h���I��p���(�q7ǔi�eQ#t�E./���^��)��8IL�q+���h��� ̾�DZ[�2�ף����v[�㏫oꕓ5M����{�4��h�l`饯Y��G�vG��E�~�4p����'ٯa1t�����ʂ�)��(+y�����ᗅ��o�mDW[w�����1[T��K����@����R�{4��yߝ��_u��g�K�+�𤟠����Zs}x�jR<4���6<1M�J�xg_��_t��{GD�=������qA��f�"�U���T��2\��gh�Q�m���>��������Bk,��a���y��:6� U������Ğ���m�{����Es���7a��d{�ۿ	�n#�����`��L����p�1ծ�!d��P�Fb�g,�*rꈚӷhC��^o���y��j�f5�6m&ŗ����>�2�7�6�')oh�T~�b���R�r�^�GF��1`�ˏAܚ���k�_�l5=��O�s������|L��$ V�(d@�A���j4���+@����ҹ�z���/M��iY��'L���?w���i���lLX2�It���9�?����Щ�RP�d�M�(mB'?�>��y�O�-���0�Z�~A!Z��?��_6m��xK��5����E���sO4y�
)���^np����Q�k�j؝�'D3�$ڗ��2h,)�UP��S��k�n2�3z����]A���.��Y���r��|�Y��5������	�������jzǰ�!�6[.Eu���w���kIy��IG#�V����8�~��+��`�*a�W��\�^'���\g�������l�iw�ָa��٤�Զ�x��`��\�8�QѨ��{�	 $�X��#pe��$<y��8\���C5�3UR���2,E�؍+@h���ٳ�E�ƾ@�q�ɾ0R�Ļ�u(�r}E�L�����ċ-�`s�!��Ah���|R��D�0JV�L�>T�ՙ��TV�Bu�^	#b�/"�4MUl��[c.��R���A't��?&vě��Ӗ|�?⮓�2�w�젨"5PHg>#�%M)�?��,��T{A�}C�����8 �Ln�M���ڱ�1�a��N:t#�@�o���͛�5��������Y{^�в���p;٠f�i���hfwrÛ�d6t��Nw�w�ҕ�e���W�����5s��T�o�|u}*�5σφX7�K�-�5g�_"��h6a_c.wǝwW���P����t�Jj��p���f���4wV�s6]���Yg{zh�}�ϵ�b�C?J�-�:��dDG�ER
R/p~2�AW*W����[��˔/�d��傯蹢��!�EHu���曭07o����1�z�ϟA��HM��wQ��+cb���x�YȦYl��]���ߞqpʭ�DW	��H�Os���h��~�7<�|�j,�gE^Y"�U������������n��jhJ��5MkuKXM�R��d5c��5������+_롙�?��[�BPzVbɒc2si��/:�Be�c.���3IH9)q}�6馳V�\�@$�+���Y�tq���5��c]j,bo?k��\$"�ἰ|�,��y�Ep��mE�/���}���?Y.Ώ�~��].���--���br�4R1��x\��`qj�VZ�&<?wպ��R���0n�#v���f5��:���l�a�RSzw��|��+�Ԟ5��nI�<)��i�}^W�h�.��EP+I�3��M"��&ث���a���(A��n��I,��+a5��Y����)#���Td9�����:�����nƌe�@VNٙ^90+p�A��<����mR	�%�4�Ň��+�[	N�1���j�ω���t�ϱ�����75����!
��M��f��ٍG;4�zq����FA�oo�TZ$&^^�"�#���.u�c
e����"[�����7�W�������;��SSĂ8u,�>,�#(L�UuǷ`��|���3��?�nR�\��ɜ�;�m�4�צ��:��GX$.���$K�A��Mz�)��q�o	�?*�1�p���j!��\B�m��b��|�,t+r3�4(M����>S����}�-��O�$AgHK��Ճ<xı	O�ֿ}�O/
bW��
�>�SM\�\㷠�ofq�� 87��8��Y���س���4��м���%�{���`+A������L�)�4� 
��4r��<,S�����%_�� S�Jǜк�-��|�G`n���h�nm��Ut/�z��/<4�t�e�{a#�^��ҽ��>�λ�BC:�u�ǵ_�m	��*Q�,��HG �He��~Z���n�uFQcw;!BnH�Ts�%�����!N�,,��l���j��OA�1�r�ʄw��40�ny	0��=C��������&蠚� ���h�]i@�^�-�liI���m*��?�|�p4�y��kT ��u���壣�iO9����T}��{&Y�w����~n���b�f�{�lpdN��<��W='���}Ӡ�r�?{S��LU�0�h�x�{�q}��@.�k?^wK*)˙��QA4b������� <l`��x6��%���y����}�D&�8�m�<?�@�}.nk�L�ƪ
�"��Ia��n�{e������{F���ѓ�j��m}%��p�^����j����8���Bt��|��0�?V�5�gY�����xk���a`2}�;�6Inˣ).{~��l̦���#��������<�,Ѻ)~��_���LD��I+�r��#�"�
76^�����F��jPV���Q�D��T��p.1�<g��i�$Wi��B��G�#�����)��1V$��P�R��6)U�8��
�*=�#v�K1�PV�|[B���ѺhO��]�O0�*fr�3t'f������m�����3�{�R�!wS�Mg�{�Il�k�e�tsͤqh�ripI�7�xV��r��-U�t�����½��̱��>օoj%�����B|7M�a~��cA)8?��Ѿ���/ ~jZ�t�EB�aQϝ{��ˀ�M�>у����"�(S*bv�=nW�H�״��j�AЙ�f5�0��
��*��X���Hd�:�?���mb2=)�M�Y�.0�[��-��+�1����~!��΄�6��I���2�s�����Ϙ�]�LF�_���N�5�O��J:=���$��4Z]����+bkV	��ӱ�7�2����= r7�;1�:ټ&�}��G��%b�p;��D@�q����T2a���nI����Ml�)�ӴŚ���7[L�#{�?�������|���䳠�����e��f�*�eۊ�� �[�0g���yV%�u$��3��9ȍ�2M�����^|�Q��u� ��K�������sJIm_׀�~����!F�ݚ-�W��������ևz�o�+N���v�N�pj���Gq�����������Ы-T��L3[ɛ�Hf�]��F�:Iy	s�����̶��I�:�ˎ���h�����5wПg>d7�	�1�z-X=�+%X���m�,R�r�I�8	��*C3q<��M�s�,�D�>��o�_ϯI>�XFj�k�4��]�y��ZSY��x8;Oӗz��җ���\��I�k�sM�Vk�&�9�EX��׌��Y�Q��Q��p���ܯ؉/��ɲ������A�������Kn������2�_?N����haq�K����[(�Ϛ���3^�*[ž'!�n�
omzK���d��-5|�Y�sT���56+sY�h���4p�z��L_�<�TC-m��x�'��L�z�&�r��zS=�.�?�|.���V�t��F� F�ܯ 4�-T���ȧ�Ĉ
�I��P������ȟ'8~s���~�,�s��fϼ\����������>5_Z�yN�]Be7�*�{�+]\Ce=�����2�Ƿa�6�>-,H+$7�@g���M=��ҬQQ������D��6��v�J��iwT�� ��^��
�q�X屐y��q��/	����=���$1�3XS���T��=%�u�D�=s��k���g����o������kl$��r�R��	��`�����q>V�����Z�ڠ�(q
{|ц~�y- ����P�_^E�u�i��Ey��t(��=�D�S�5�O�j}Q�׼�,|�}��a��|2��l����N�j��,ql^-��9S*����`���?n�A:�nd��]����-��\$���U�BN,7���1�S�5��G]1#3#����[�/�����ح�}�i�GlS�t6yT!~H	z�#�IK�����:���<4g|r����F-��v��n�HH�P����~���Z��Њ~��w��1��wX��T��MV�kr�=��{��"�(�u�I�/��,E'k�DT��eʭ��y�� eώs�P�9F����;�������E�P�p�Q
�%�@�,�n�=��������"7�4�c�m��U|;��=N>�9�q������>�Ǚ6�����bק��%�@�{��Y�Y}.JRc��.��O���v\�H�?�R��wϐ�1�E�E�m�s���&ICb�s�Xܭ/��>i8.�4a�/L�7�v/�f�٩�D*�Pj>IaMe*�͗�苯Ϳ��pҊ� ��IڱL�4Ԭ�㔝o�B� ��2�1��݋u4��A~K3�����ޱ�X�zLl^+�(�H���űѽR~b~�7��l˯��'=���.e��+�U)���82��ĩi�����4���?��6;b`�BYYqς ���"A��c���~U���:��R	ߒ*L�lv�'?Kc ;�XLX��,"Wb�b��ږ�w�.Onin.r��6~f�w85��e.�5-A�;�G/���j���=�z�x"���e[7d�Ga��' h���Oi�w>� (�F�Wv:�"��|�Y&�&����-�v�����O��U�(���'���:|k X*Y(���~_*����ΛW��MA>|c�N2Ծ��Na,�'*����F��]?E��L�V����ي+;���U��@�C`�~�h���&򒒷s�� �T�_��DF�L�A.p�6�m��M�/��dF����j�)	�/Z&��#�1�a���B���3�Er}6e�|�r�Xl8���-�0���9R�bw�~-�0c�$yIL���w���bR�%ɶR3ݐA29���H[��~wΩ���EXw�_=:1�j��7��ޚ�);̑4
����b,�iߓ����T���<��i�� XI_��r/�W�j��Fp�r���S3#��9)2������pO�B?}fk!r>�gT%��y<v,'2l�$7O�SP�iA4�?���?�8���j�����%�U�Ź��T�;(4e�������>E�seS�V|�v��#���z�����ժR�F�J�5�V�R{�M[��$��Q�ڛ�M�P{�xլ�6;[�����?x��?<o�v;���u���~ݮ�zJ��3gX?;�ܟc�Q�Z�`�b������WJ5j�.�����	�[�̽�'��VI�����ؾ!���&���j�� �����?�1�.��c�"�xV�s���*��T�x���C�*�E;q�H�z�TK={~�ی�^l�XI�-Y259��hNm�o���/j�3k�X��r��8��;M��y�g�=�A��y��z��vfD��3ןn¯�M���Cf�WT�祦}E��]��N�{�?�?�s/��5:��@�Bk���Z�*y!c��d�i�%��1
m��QBּ0Q�7&]��|�_�����n}��S���|�˙x�C�2()�
ھ�͜�5��},n�E:I��_�ﾭ?���3�툀���/���{��㉞��Բ��lf�QR�ګ�kc��H<���94g��'Y����E�(���^n�3���:JX���W��:��=��l)R�����OdI�)��.�v���?Ͱ�o�����|���"�ϵ=p���2����2ie���t�K³�}�.͌�����?Y�2x��W��.'���_$=Z_b�� M�3��l�k)Y���W��1.�I��dʾ��D���	V�?���l炙
���%-j����q�� O��?]|Ag���V�� �0�җ�	/�r�k =Vo���f�}n���jq4b��H��%Q�(����֔�dߠ&����ǩ����O��
g� ���Q�����ֽ��i�U���6��S:�ņ�H�tV�+��=5���<x+G#��*��إH�TڎqO�=MiԾ�B���?���J�Q���-��a5�ӯ��LԚc�3Y������r*QF�!^��-d���-`W���&��3�jWg�̋ڷ2��	��#[�%���V=��Y^$��V2i'�v	m;F���1	� �Jስ��z���;2]+�Y$I7�|���p*�yD�sݙ�0Ifpji]DD��^��gdHF'���,�+'�+�\��@��4w���19�=~� ����2]�TG�F�F�����[�J�%�í�ni���M��w-ۼ2-(͛�t�d�p	���:%����n+ZO��B���D]	���ܩ�J�V����m�-�<�4Oƺa�9K�ץ�AY
�:��[���J�HЦ ��0���2� �'3�K/�����F��$�L�ҭ��}������(���˺{is��=z��uܿ�J���20�"�T�|�o!��|*J>�b�2-G�i���=�B��ԏ�	V���Hc���Q����7cI�$	�xv��`�}���WH��ʜ.�6���4P���g�H���A���4�$�BH)xx�� p;0��i�'d���z��%�f�M5�.B}�� d�|_ޱX~����/�r/�����2���,�����WG'�d_�����H���)��o�����Rc"�z�Q��H=ߴ:�n[=� �wBn�����ƴW��~�r�=1���23�]L#!�'���o�����7���_��[d��M�!���	���ޯ������,N4�N���;T:�?��GS:�N����gE ��zX����U�5>%�6�Hy[��;B��,nϦ%�ψ�������.'�ED
�<��O]�۝+�G�.ms�8�8�]|����H�Z�A�c��1�=��Gt��ʧG������sHs��M2�_��RSԩ���,l)�0n:5#�/���o�.����8�a�e�kp뫔_��9h���nOt�vn�W�ݺʞ� Hb�&��?��a;�FM��~_��.2q�%�<�O�a�"Pt�^��ԃ�2�wn����(�C�}�zV�����p�v��:OYm�\��ܒ&�:o�fh�6ȼ?����XKå� xv���0��
���$�**�ݙ�� ��o���t�r�JD��w�r�)�F��k���f�/Dx�7�U��{x�g�b�5�㡠�g�W�/��eʣ�G}D˱ p9�w"�UN"���ϳrZ@E�{��$��_�,�������j�:k����g��3ߠ!Qڭyұo��T"cl�D�k_=���%,��{�K&4p{�l;�^�Hm��x�3.9!����~bj~�S������-k1�ݚ`v�K�Ø�M�T 󆃠KΘ�\R�C�b�@l7��!�����CC�!V�V�ж'�:���ӥ�u)�2�'B�����?b�o5/0�<O�'��@΁���H���
�T�3d��qi�E���?
p��*VG�L�zh料\B|� ���� �߅7�`�m[�y�T��<�^�2wre��&��<ͼ��X�DgNv|/�"���c<��������A���!l���8�0�,6hbg��5@�u6dBw������m��X�h���;}5��ZTT��m�24����a�4���<+�ՠO3~��Z�3)��~��ݓԋ��<@R[��#;�Đ�~T}GHq-�#Mt��4���c���Tf��(|�4��va�����d��H/T����?Y�k ���QKM�>#�HJ�C��s+����婵:Y�W��4�'0(п�N��9�� w{�Sv�N*�0/*p���8������GkIV*8\%��F���ó~�IY�C���"��q�2�U��?��Tv��w5����l�U'j��X*0kT�[d����u���>j�dg3rlQ�k{��5���|����7E��Ş���X��i��O����l����ѳ�-�po��:������:&T�v5��Bk8c��)3��n�����^
�O6z�-Q����3*�%^��/�٪e�1�;�V~�M� ���%��+�U���㫱	����6Ɲ�H��GEO��*�p�n�_���W�/(�|���\-ةB�r�3�P�����Pd�c��\�_�7�A��r�NK �S���Q�B��zm�^o:-b�����)�� ��3�g?�����U��������ȴ��f����m ����� �7ea�ŸQd��|V��|�J&�]Q��m~y�t�T��<4Y�Yu��^{�k ��0�Pe�
s�WΥ�L�n̻[��?԰�<��|�i=�Oh��.S8�ʃ���Ylݷ �`ˋ{3�
澏E�?4Q���'r ��j�v �b�g� �F��G��$��,�-6����
5Fy��}�7�.��է&{ew���am����*�i�)���W� S�w��{_���m嵦V$�DM�t؁1��Y�w�+�K�
1���`�kW���>�֊�gL}���4�|S�S�*�*�#��[V�(Zs�J�ԣ�[�=�3�Sg��jS3T�	0���{�x)�YqF Sm)��S;�8����u��5�����#{#�qT
Ia:���%�i�������Ȳ�OY�at�:�tf^+�p+�����a������7k��f���m�77����w.^���E�
3e��F/�y�f;��Z2��"��|�-^nB����<k���������^��E����������l���~�7_-z�^Lޡ��h�q��E�%�J��,�<^�~3F��M�۽xr|/�X! �55n��1'\�|�C��Q����R�2�팴>B�������'\��#s��g�R?��8���_��-3�6�;$��K��k�<�&����:���5-�12��°�:3T<�� ����	�sѥ�I�i���'
�V*��=l_���<ZlN�*~���������gW�S��G��k%s���-630�{���h2|���q�ߊ���������_N��e��G����7;�Eo ~�:�KP�$Ī �U�u_g JK,��[��n����z\,/�R�)�3�H���w�dXM�|X� 6���+6�xȜ{���:�l{���������2<�FW�� ��5`ZW��ʒ8���4�~;73�N��l�@��vT^�m����������s�h6������O$:?�-<�L�=�1m���cdU-��n>ӥ��V5b�8�}x��3���PE�ć}�n�����,SS�����ݮ���q�!�$�SQ�_�Bq0�>�rR;�A�t$ï�]�iV��7�c��Jյ��&�4iB�߸�?*��4wq4���%��t���g��0�ՏG�-�+)6�w�g~�~���b��ԦM۫ϸ�V��.��ʪ��"�$�������r������¯�E���Q�t��,7N|��w����`��oY��iI�E���~��gJ�r���Ze}��g'���Y����sLc�W�E�𭯨Ðf�V��ɹ���C��d�#O���Vs�q������D@�#�{��h��=y��G��(ʥ`*�6�޵���NOé�:�g��p����z	˂wr����2��m1A�"�}���	X�g���մiz?�S��)n�|����A��}d�O�儾�*�qK�;�,�c䪺y
��TK��+eϙ���A�g�k@4�F��xbF,��L���\d#E��������j����S�[@9�-hڶ�j�0jM�D��<-�&�d�dqX�}���o\�q�8����0�Lq�����{a�w�K��x�K~��ɍ'��T��I0/�Q��a�����B���#YK��C0���"�-��F�Xs�	���0��:��]�(4���KV���{_H�2�w��������/��l�ʩR�@�Rp�錓�-�-ԙ�%ϗ ���ު{>�����?Z͓��z���K�u.~M���I�ӥ��xe�Lʜ�QE�����UƈU9�@�tc������g`7?��H�?�::lNr����&��z�����\o�`]b��Q�Ւ͒M�g$�Q�T�Um�0�A�w:�KꞫKj=�+9^�
���:F#���d�����:�{[#Em���;8���TR�QD�eG�:b������_U<��
8%��j�����\�b}6o�ȜVz�����ϔ�������L�.�ݼ�3m��y��h씂��
�2�÷�B�0�|%�ދxv��Ǫ^f�-�~�����5��Z��Km�ݰ1'��{��$�ވ�P�=��^m��]��E�c~(��K�[È��}ز���L��/ ���3�ٵ�1Y���*,�qA[(�G�MX��̏��<+�VK"����e����<�/=��{�����~�W��(��&���;)>�/��7}x��$o�x[+�8q��=:5(p�ٍ�]��B2J� p-���F���6�4x�A%�+�L�-(�#N�H�e�;�����9��X|n���nx?�ړ���Z����j��&Sf��
'4�qt�I>�p�����S�x�c�˕%�{K��}�S�?c��1_���/�9�M ˰�\ʺr%�=:��{?&%��o��[�7��!�_�(�n�Ѷ�W�%(_��y��w�6�IkY�wu��D'DҍP�Evɪ���� 9_�~l_��D-](u�&ɑ~~��v�<HO��W�#N����6���CbR���Z��u�o���6��R����Cy�qf.�Wg@�M�#�8��Rsb%*N��w�"Aؠ���|����D�L��I��3W�<��鮵�5zcU�T(8i���VK��d����]Tw+�o�<]5ٰ:�V��.�6���WS��^�UdN�_!�.������;b�i�hX���I���d�Z,�>Mg��*�.q�P�ף��CP���o����W1��I24!� ?�K�K'-X�k�&��J9^(rI�z����Q!����v�GI�n�!�l�g��ӶXs�X�^D��@}>�O~������s�&���n%b��ցۊ ��gM��Q����*�3�x���F�Z��PW�!4�pT�=tj�7�Y��Yx㸛�t�,�`���%�&�r5.��`�ʟ��2V���M<���6��LXַ�M\�Ǳ���k%]��eQZw�P?�m�����wq��مI���p�a�d��u��k�3�]���P�7�J�M l���C�Іe���DΞ���1>�ϼ\��Z�Dپ����h5I}^e�|��GvrճXd�>����c�ӥ��?���	��C1�D���Q���6]�����4����߀n�|�ۛ�����G���^�\TʥD�*z�T��:��j�
#�M�T�e��R�H�z0��yב�&pM/�#��@���8)�}�� �������o��ӿ@�<S�7��W}0�)~f��+h�W�d���|��[U{\�����nM�
#��Z֠;䨑z�GW�n`��h�,�P$�f�-tD@�{���e5�\`�ό�t�_���c�Tc��w{t$���cSN��霗����.o�����6��ȵD&��xgw�d�nߊ��Ol��X��sn^n)ڠA&=��Y����q��B4�[��������T�	w�g��b��.S���2<�P5ܒM#���⑑��k���I�ۼx��-�w1�q{'�VY#��[/�^��x�|����~Vn&�P�
O��d�Sr�p��SI�0��75%��r�+�"�Wڨ1�u6'��A/��@�j�����b��Ɍ�>}�'���Y�˹�`���ԉy���*S�"Nד�*zJ^7c\�[��~�褙�A��G��kf�_is�r�p'zTh�ڈ�{Q�T_5O� j�SK��A��
�J���gW�;�V��'Z�2a��N1��|E��Y�0��� E�ɼ߱K�z�w�xcB��WZŚ���y�J۾�a}����ι#�Pp�?F�S�[m^2�լt!@�})����]�<�� ���(��iSYgP�TnXVe�6��#T�+r9���<��)�i0�Ԓ��n^�7�I���Sń%�������]4~�@j��1�R�������Ϡ�g�	TA��۷I2�#M��=�"+Z�0�3����x��H����"�#����?e'As4Z���[A@v��
��}�������i-5��*���zk}�%���k@Z0�|{�R���ڙ){�u��镠�>U�_�<t�N�ѹ������\�ݯ��m�?<)�I&�Μ�ff	��;��?=n��^�ͬ�,�ߟ��RT�tWȌS�'�+�Ѭ�_�vx_��4u��H��/���'Zu���=V�rs����ޟ|s!��{s�a5�cȅ�NSRo 	�\]
{{�֠����D��[
H��������L���ZO?sv;s_�v��"6�̓I��9�ӷl��7�q���C0�FC6:� ���N�]CL>iɫG��}ur�u�we����U�	xfNC\��aU�܅�I������Z��P��k�Vk�S^��b){A��NJ߮v����{���5��,�e�g� ��8��t���I�~a3�35C���Xq�Z��˃���c�_8:h���5�`�jhU�s�F̑ b������ݫ�dZ�:�����j�>҉��ݪ�����b�#{�л��������%�)�[8#W�;]��h��=����j8}����y��LQ��Y��2yܳ����J��򚘟�
K�Ő&���BLA�5@���~���@�.�0j�� �I��qC=]�"��sÑ�{o��{~᭮Ҹ�����ur��(�`�.�]�@��ĈʾŒ��z+�Ib��7��.�#	з������ћg׆���x��x�}'�9�ǲ�FQ�T�#��}R��5���A`�#����N�K���::y���v�i|�dl&X�8�h�A�oq-p�ʥy����x��F�X�e��l��~|�?�{��_���_"l�[f­����8�����}JDY(%�x��Qkѱ��Z'/S����?sfOq�Nqe�ѥqU�����i�<�2/�D}�4o�q���nj�ɚn�6��U�TpXE���ס��WH;�_�Z��X��xC>17��j�c��t��eXW���O�f���`>�f�M�Pd�����W�F�N���q�O��ŊPB�����yM��3���C�wSE4+ �*�z���ui�ˎ0����#}9���*0ŃF�_��*v��^����L�S��t~�K���.20��?(�m��rk�)7W�DӲ��i�e�W�~�'��*"��k�J��B�Ͷ��ܡ����n�o�O	�@;j9��'��w9����$~��`���!an��GE�6�H�Y_�	ׅ���
w)�`9�XՇ0�]z����|�DaǕ�5��q�	[-���ak�!WYda�sq�"�������$g�ר���6p�	�v#��Y��%���٧f����
���94S_� ��q� ��'��?z�]���-sY�X\����,���e�0�/a����	n�a��W|�i�G��6���[�d�Q���T9�7T��A�\����h�T�����W]�t'�ޑ��-�7�gg��!�4
>���-�:2�H�d�pmu�������zI�h%�t����b]}`]?W9AP�����,���Ds��q�q��}+iS�ӐũH��c�4�V���b�tr���ی�R��to��\=��:.0��ޭ��fz�uT�뗧�5�#G����9q;������/�Z�G!Lt}{�F6Y�Ҧ��f`qOľr�k*��S8>����&�?|o5�(v���br�v�B�d��e.鶺���*B�9���7\2����Y��5�Y.�{޾s�V��m7��5�ؚK��൅���8�S��ͮ�����'�g� Ƶ{���_<��D��`�u��eA�v��6z���f����)���X?���q߄���o%nyw�G�/���v�D�rb�=�E�������7�/Fd�؁+o4��?K�vm�?S��v8��|3��ÚqN
+
�:�[���Ya�vsհ��{���>�w��uR�Q���؄�m�����$ݠ�(-N�щ���pEyڟ�� �0����f�dE�?��:$�c=�w�?� "�SdN��t�~�1LT��"���A�����~M��������>h���3��GO���"�z��(��6��+z��4��|��ɐk ��`����Rrh�C
�!^\����Y�^CҀ���3��v��)-vҹi�D��->Q��Cg�9����k���kz�T��+_O�9 �����x
Q�֥��s�&M�K�����ސ}���B�`M�:�x��|j5]�w���"����)S4:��5i�5���)�b�}��� ��\��J+k�-ֿG��Ŷ�`���i3��e��X�cZ�{f7G���M��E:��\�cǩt�2�>�Y�Cs.B?���Bk�N{���)��{y*�,�n ����f��흸[�&�om�2J!���p�<��Q�p���pAg�I��q�u�H����q��X��T��&:P�+��]�P�뷾W0��i�da���&�q!W��5k�&��1胎�cG�:\ؚ��2e�l�r����X�ӡC��%����R���S��v��B�"K���:����G9S8����q��ֹx�y���M��a��x^�9�ڗ��q�`1��iZ<������Y���!F
u�Ak���7�]��z�(pb��U�s[C��鍑�W�x��	�'��e/$����o��|��%��#a�'��3/���K���`8Ë��pllA��@
��5{z�N��Mzi�����-���rݷv��PXّ���|�s� (�t��ӊh�pSLB{S.ú¯O�_������[��A��G]@-UCr/K`\D�]bC2q��.���E����Wn�:��;�`'�4��u�8�l�������ا/� �o;�&D��P�WN�X7�8T16�#r�GD,?b��O_�����U�P4���(�V���8�dq�] �}zr	
U1�b9�b��� 'm�5.8�`"Kq���u�f�0q2)����3�7�3~�F��p{��\jX�E�9(�����E��@k��Ix�J߸o�oI,�p1͒�Y��Oy��UU���O��cqt�=/ݰ�`�:	�#���sd�0 S#T��O<ɴ+��X>����Sf'9.� �{k�!�|�o+��T��Zo2=X%�r^�{w'�$�~i��R�\�>��\�����$:�ɲ(�/��)���s�,>Gg�n���;�0:H.���>�����m¡�>Ub���8iR�}$�?\��a�Y f�^��&,h$t"�(��d� �PXGB:�<������h̲�FZu�I�-d��q�r�A��ɢ��3M��l�}�x��u��D�FÑU�q濄oQ�hf��.#ZO����="�Zz��G��E͛��-�m[��@� �=��!k�D�c�����mb�vg6�2ND����_�qU���Շpf�_���ɳ4x�,����&�L�k�h�Aj����B\k&�>�2/�a�I}��Rr=�sc7��|��ng"2�썆KD-�����ߌF�o�/��
c=�lW�hpQ��(�\
���mE�b�M?�Ku(����2H��>vx�X8�g!������Cq�D���]֙|e���\C��fccD��o��Zed�g���<�w�H����2P��k����c+�M5�p�kC/�/�؁�`��w�jh�y}�L�#����T�y��K�+;�7F��@�`�c�i�\��xx	�+�nS9Ї:N��V��'����4��EF�Tm#ί�Ù�<���y�R�"�LG�p�Ȍ0K(��)�~��T�.�*x�m�.���˒��[(J�l�Y�;��u��9hWaPSXz�ʼ�����a)�g��@�]���+���T&�L�j�Y5��"��h1hK.��1��Gk:������k@�kk������{~�F���/�_R_(�>K^��7�Ts__�?�}5��J�S�"�Q�챚�u`\,�9w#������ۜ�'�� ��2�^<S�,0{ ?q��u�u���V��B���j/u�%,7�(k��y�+��{�+M&v�d�&gA�ov[t�� �l�Gк
��[P��a�������r����R�\@���x�������J^�ea�Ϟ_��Sy���l�T����e!F�_�լ.�i�\��W'~I��Y����g�O(uwA�I,�v0 �p˞��੥� �:��������!��tW����pߩ�4�N�x6��#����6^���L�7{�䔋Z���<-���&m _�-nL�ૅN*X��s��}����=���0����0e�}Z��!w5�	6��%����#e���׾M�9r�+��|/�N���}��=ݛ_�wO\ȟ�6,�J��i~3���Цc���c+��D4`X�8�>�zZר,кM�0���k	�Ӵ��DTW�/��{�-��HI��)��f�|��׍i����B�Ξ�Xk�znԧ��@�G��x��hM�F�F笔�U1��35?,�`F�|!���EM������*��a���@Ֆ�M��z�� /�E"�ݲ᜕�6	㐿g�dwcsK�a(H������×�--Ѥf��r�W�;vA�X��o�?y#ps�*]�R�ֺ�g|��5�߇q�-^**&�!�t�E��e�

�03�r�/��agK\<����"x���|���3��#ƽi��r��D�P5d�W�!f/���]����s�|��-��X�j�@Ճ]Cr��N��=��"@t�x��.vP��mocK�p�����o	mzݸ�x��a���k�&$��6�.3H��	��&��_{��5���jo�m��F�W$��Ol�.�p�LN�r��U���#`|38_�Ś}tEշ�I,����Y0d"�Gc�x���I�]�3��(��,.�����Y�X����5�?^����;�8��qR��!(����o~u῭��ؒ�d'y� �HY9w�u0�t������:��������XH��͝V��͗��aS<��×K�rfQ.QRh��2x����[l���.��e�]�V[:B�K�KBͨ
V�~@��.����̽��2[h{r|6�F�ǯ 8s���#��yL���8��F���w��5D�7�	e�P?��o�x��V���2&���u��wU��F�p��{4�c��]�#\s�����]1<n���%�x%�4]�A:#H��T�.�~�㧣�J,�	U����5`�@�%�$�������+hG�C:ѳCb/{*�F}���}�M/�Gx���#������07~��E�ͮ�j�r=�q��d�ϕ���AM�M�L������:h��k��|%\�>�y4��jŇ��5d_�i�|�$=�������?�|+�E���QEȭ�N��aզ��HGU��{��|��5�Ȫ�e��tۀK3�n$��t&_���zE��U���%�w!}	����ǚ+WU�(߹��@C��)n���m���t&�K-�3�,���Q�%U����p�`��c�˻\�)��ߺ��RA�P��U�e�(,��|ipH�~���S	�pj�|-f��)�}���%/�Q<��PqY���6�^B��a�S$/3#��n�-~�fFM�w���Z%�\�z�`�r�)���N�7��,��:2���r�y�u���%7>D�?"G�hla�oP=�˶]�����`I��@H�
EaX�2�>�1��0�XBD�T���3�I�L ��ȋ��$8���0edh�lՑ�y�Y�$lPr���^�M%��xb�8�\9���f�h�ȥx5�e%u����o�q�A�m���̷���y��'�%�*���Mww�YY]���!�<�U].'>6F�%�m�id�z���&5�@Ё�Jp~C�\����V(�EwQ!�fؼ�!3�[��z�����B��dJ����>�U;2u�#���Y��D����ͤkHx�lș��5�L%��Q�˲���+�j�;���e���
��(����<�&��3|k�7fN��W5�Z�ەx�>^���^K��-qL��u!h���ՏRp�(���ob��w�%E�>&��ޱma��A?K��r�/�jFy�Υy�\L?ìX0V����o���|7^,@FUq��4�Wc�����.G�,�n��ut�����'�uUF���zA{x�=@��T�;�a>�¾o��`W�����B)�t���$����]�o�\���B�K��Ѭ�ICbkt+��9��3w4�$�=j�Çs}�������g~���{�N�v��	�|�u�4����.�}��Q��4 �W5��l	%*��dk�Q��@�����`#�9��r�m٫
O�\�����+��F%��2k�n0̌Lr�V�n>�%Sz:>v#�;�RL��F0���ZKJ��Xw�AD�cGn��r�J����W�o���=ځ|cL�~_|f. �C;�����g-�W��z��Jï�*"��e��~M� �d,+L�����Sy��G�T��Ŋ��3�{�w�H�*��SN�Bo�<���~�G�e�1Q]hvS�œs�z�D��,��e�YT2�6/ρ~S��� ���y�6*�����o�n��u��SV�qש�L���Z�d�?�4Ǽ���}�g�Q�p��P�n2���F�&�n�=<X�]�҂�����>JE��-�M���kg:O�J�O3o��1��왼[ɪ�������rw���]���{#GAx�Mg���(4O�,�<|�����8�Xg�͑�'��P���Gn�A��Q7+��bA��Gr���������"� U1�m�7�W�3yLG�)8?�!��Κ�au�z����E�� �b�o���JƱӉ*��ߚ�?������q�;��R� �'�d�?��;�}X�[{���(���dt��W����#?�[������Vm�#)�����������Tc5;c3N��V;o��j@��C�U���k��C<AO�|@�Л2�g����Nꅻ#�+y&Rqܓt���m��,|�jYi�&��ǫ��� H��3~��x�\�mN�d�D��ۨJ�Ր7���E�բp�(M��/\O�uj�/1kn�� ��Ь��{�	�b�Zz$�z�*?C���Z��K=W��`�H�Cۦ��t�#kE�E�ܚY>�N��<�����F�I����r�[����Y=��qp����.�hJ(o:��2�d��@��@[�A�=�֏�&��BJ��a�Y-�lS�cdl��3��Y@����v�O.�8[n�^���az\�I������$�.;��(�K�s�u\i]���F`��<�0��N��&,ro�j;=��d�k��]Y���yB?4�|�q�	��zʸ1���vu̺�ڋے�c�A~����y��!N�}[I\ɸD�� u�9Tx�)��X{��yU%� �6�n���Y�9rs�|����n*[�Q%�?P��a��I>ܖ��q3>/��L��&��p3�t����uV��O�T��B���F��!�b��N�*T�}B I��?�䈰�Ԇ���U�WG|4.�U�ȓJ1@��qFR L���e���%o�ڥ��EW�4�L�����$��"�:�u��J�D67!f�G����6����e5��~�����@C-����1}��a����Bs������25-y@D�@�:�g�H��Ĳ��VT�.�2X0�a`�<��v.�ఋ>SҊ¼f���X;2lĴb;�[a�#�n��*����F�z��0[0i�MF��6ם���O5�r�D&�0�k ���{S�oy��x����n�*��c+m4����j14+k&��WV�TVP�7ɥl�J,Lys!�H�Jw|�0�1 �3�Yb�<Ca�.ʈ�H�eڒ~���x0b��p0������.y�M+������`n���m��������;&�f�J�26S������,(�A&�?�SA�+�6	��ָL�Xceѭ/\(b������<�*
��?�`Q�$��B;|�[3�Ilg�}��6V �
����TV����H3��B�f��~V��
9ٓ{���#�F��:��M�/���:��˽
a�=�9���� q�#h�b��w�>��7\�!W�<eb�KQa���y�	��=�]@�G��5d�6$Ĭ��<y_x��X�zn��@I0�R��>ad��q���1��K|���!vX�<¥%���#��{��VJ?OL��k~@,"Wk/�&f�x{�J����#jG�}Y��3�,/��RG���5�EZǶ޷�����B�κ_"�n�[���!�yU&�R�Ӆ>����%(yj���Rf,�	���0,Ɋ$c@�6�?f���1�'` 򯣌\e�wU�Ê0G�7�a6����J���?�1�z�N�|�n�k��"���[��0�u��K��W�uӬ���7:���A�_܎���r�)1����{�P�;�Uk@�ǡPiG��A��8`�y����5�~:dp�ʳ�d��<� .�0υ�\sP���w�&�eIQ�=���X/�K�.f��k��ƪ���2�O>� ��NҞ�j���������\�x���"�r�jKb\r��n�s�����/
X�3�MV)���E{����RI�����-�k#����6�7w~�n��wN�`^���j��{̛To�k�{=`�^�Ќ#!?I�[������y�q����"�36��touKr�2���S�r��g(��u�J�,V�@�[~� ��s7砲�W�*���A{g��H;s��j��<��D8�S]��ބ�+��'J\j�E��S\���Z9Sig�1>2ι��eY�.߿�>����RK�Kτ�
�7H͕�v1�>0pz �YMK�����K�0|�Y�ע�E�	�����I'�f׀��#/c&���s��B�0{��f�jw�8U {��a�iri�YX�̭�N��j��|z������^��iY�?����?�;�*_��cȗ��� �BL�rr��qs7t@g�$1qG��d��g'v<��HB�T���J��=��䊌����U�䇪�hazq2?�4���j�0��mbE��4��H=s��:��I�~t1�v��b��g�m���捈�� � ���X����Z���s�r�m+����G7���ydL7�ʑm�tq���J��tA���|+�|Y���<O�O���ӷ<9��G�3���U��b�5 x�(��)U����q�m���+ 9���o(j�~�Pz�Ӧ��m}��~��D��8�R�>u#|��Z��0�����2G�|�ʇ%4e�S�|�Bn���.�����_���?ZADP@@�J�DZ:&!҃��i�RC�;ǀJ
���1p�;�����^��_�9��v]���p���)�šFZA֞��e=mB@T(�^�u�,�y��'�I�M��a���4�!��o�Ɩl��;�s����I��H�P̔�R��8�Hp��:�z��u��3yyq��z�*�����߉>Ѝk&�[�YDӟK�|2=\��(>�1\YGB��Z��8��f�RW�u<[&p��pR�oS5�S�3��z2�p�@��,��]ڤ2�|C��Z�.�3Y#�6v�~0�<��i0�X��]J�{|��ѭKtşc��B��d�G/�h)�p%�Q���JT8(�#�����t�'M?mv�u/���? X�#S8����I��j�lʣ�Pi�~@�a�l�Y&�F��vm(�@�q3B�M>��硆�����l�]:T���-A!5��ܔ�J������we�ҟ�H�{�7��v����`�DSޅYe���YT��ҙ�p� �װB�x���
��D�^R�܆�@��ۧ"@�&|� 塂���in��ho��/0���"��Aĥu�����-����k �W�������Ɏ��Rj(�����>r:Y�`�_M�hQW�R�yk���Y����\���{�$��<�"R����K�����5 ��z�;��Y<%�������@��k@���pl@ڐ�RTmA�T���Q3G"�1����;��m�%��9��Ri ��m�q��	�0H$�ȼ�h�J� .�F��PSW�V���� ��{S��o	x��r/�쥕�Ds�U/�x��<��+��$vZ�&��Y.�|��'�o.�7G�:��� �Ȳ��Ug~29z%��Syd��lˮ�n�*�4��3��,:��F�\½e�ȓ�}���p`س�Eݸbs��p S]<�ǥÔ�6ȖՉ�cZ0��'�������Q��;��|��c�H�g	��WH멽qd�����;�I�k6B����B�.A�V���;iX���G������|�'�L7��Cb�,�w�!_����e�U�a[F�y��if���]��V��!���
M�;����0wν�g��	B�c,2:��V��w,y��˥t��y��y�En5�����D!��?��t����,?,�r7�k����x-:LO�wů���L˞O���ͨj97lp���o�4���XPa?Y���D$LQ�ڷ`b,9��G�|H᫚�?����~f��&!P�!�$v��h&��	�j�[7�i�w\�}ZQ�����[���cx8�}��c��}��5����eYM�3�[�1�7ye���X�D�\5�	�~�;���*F�aO/�!	1�*�4�>0�����s�;"u�ϓ!^�G8���%o��t��_�'�9
�q�i�ZD���]U��\�/x�6n��I���������w�	�E��X̺[�7���;*8,�%h�?�,!K��r_	Ld��_��ܽ۽3ʥ�F��f��]�Y��*+�;����`�#��*	}=����E�35y���{J��|i�������\7ڵz��.�r,7M��Ǳ�f(F$�_��ӯ�� �!��[�kz�v۔K{���)�w���in�@a��q�浖�_I�[�ß���I��{�Z��m깋�ebS�ʷ�5����K2��bS)�ڇ���2�+���\����]t�`,������j�����u>��y�y�G[M��@���M1m/B��i9-���$I	��$�˰�;��:�zs�Pa4���33����π��O�őa(��6t�K������v�[[W��=�#��@>���Ҝ��8����c��������$Ya��>�*�ve���t$��45u6��&+n�b%��:� 5=} ]��0o6�S�\�</;zoh���pV���@��Z��rRaW�N$���N�}G������Tpp�+${�O�� !N��!<K��v���&��.�{'ݬf����A��T���&�S��5�\IۼE��4��ٚn��H��ƮS�Y[_�[�n�" ���z諺Ƀ[�e�����eq����˰���� z�F��k�@�n>������m��_N��7�,{'�[�����"P�cA	�p��{g��'��4��k�O�9����y�i�w@a������ݵˡݭ��"��k@��3׽E��&�{3���	}��#�*er��[�ޠ��R� **��IC�R/�� /����9�G�ȧ����Ș�qd�ʨ₮��E�����%o��A�M�����ĉ��h���Ʒ>������|��oc?&�JuqG��_K�?2\�u��c��+xL㭣܊�W6���h��%�H�3=�<;�Z�|�<���O	(��j��R|��b�`w�����ޫ/&}�1Y�|��U?�eә�H�i��*�$37ęp�r��T�=h����c�3r��;���A��yroQv�qc��E�M�&�ȹ��k@脉���]p<�ѧ�i�aTbD)���j���0�ߝ�JR�=h�WP��|��̪z��91���S%~Փ.ض���n\���G������G6?�)F�]�]u#��y��Ϲ��پeW�mF�TO��>B�,�S��</W�OL,��<pS9⡵��"�x9J����1�+�#d�`�砱�՘��Z��D�F��jjhg��ud�{ЎY{\�]l��{.y�q���-�J�8]�Ho�_���g���?�ԁ��/���UI܆ߥ��5�m�7��͍�/�ߍ[�{�=�������;p6���t3�K�����`.h�_.�1,|�Z�;Ա�!J!�i.z�{��ŵ�O� �H��OHM^Er͛L ƣ@��8���WS��$*��t������^~�����e���i�0�f����QZ�}�
��_%h˄R��K�:,t�a;��!��i:
`� �h�c[����p�� �-�M������k{�5�f�<n�I��0���~<�ز�G����Q�����ڀ���l>L�1��\�B�;�A���7�E��<*w#I�dѰ;����_	�K�0����|Bd��/Q��0�\.W�Qi��D./ �vO���`i���,�c����ů܏��������n�ZL�-I��r`)D� ��B��-}U4�E~cYSZ�L�[׌��7��}XIAH?a�g@�1�����\��(�$�^U�v����p��K^E��\.��F[od�?��ܶ��Γ#��+�����M���=�O�T��n̍g�����Y�	ܶ���'����Ĭ���Nh�Ν��t��XY8��*�� ���qW{'�M^�m�!��'y�٬��y����+μ��p�&�aُ�Ʀ�\�'���
�iW�d��g[8N�q�o�<ߠ�^a�D���"�b��	#��EŔS�xi��'��TS.'��� ��Aq��.7fߟ51Z��_���j���f�}���d�U>ZV�?nJ���Z)��:���|Y&d�=8�2������G	���r�5��H�zN�j�r��v�&W�Z-8�A�?���>w�p}d+�bRu˥t�!S��H�NCq�����KQ�չ�gL��o�z��D҄$��'5��Ci��.�_����n��&&����>�>,.!��J�ޑ;����B*�'�c�����Χ��`Yή̸ZJ�
o�D�ǂ�7m��W�VD��ׂR?�B4��"�O�ԫ/��3�Zm�H�%��8��Bnvű��2vz��em�˿���z��,��ĉ>��D����qXm���, �;��s�_Ӟ��Hb�,�#�M��گ:*ބ�Z���mI�1�
��O��ݹ5$�h�Al��F4�n�/��=����E
B���'�@��v0���;2�yX���{SS�/J�!����{�0?�Vx�f��J��(�?62,�ڡr�n��ƿ�4֯$<|eį�Z؆:�i�]}E� G��/����##�*I;2x��y����Z��P��LR����������$߹k�ߓ�L(�o��Z���([I�����Pmq���̄m8uX�(pbvXVJ^�<`�e�ڬ��ީ����Z���9�$,6�j<��>�i�P>���CdvI�.��N�e �_�0�ύS/�h~���n��t]q���oT�rL&;�-� U�l��JF�|<� �����^$��殷(4��j4���D��|G�R�&�ݒ ���geFxb�ĸT�=8�s�W�ʦ��r��.Ĵa�4J=���S��70�!�Q���'�>����p�!!'��l{S�,���˦���s�A@��H~Ǘ�z���_�y4��-Ǝ��O�f�i5M�8Ei��Z�|���}�Iɷ\�n�Zfc&��
C�Q�F��r�N����g���n?iZ�%�T]ܻبu=/d+ �ʟ�������R;�ni�ADL}}K"�d��W���{�������z�9y%q���W�/G��<=@��^�?��(�-0�8�~w��ɏ�yiM�O�����١�maBBA~��!��w$��/Zk����S�wY���=4��������h:�Ҩ'eMi�G�KT��j�ɹ|\�+�3��ԯ�B��e"� 0���%qG����1��#q�l�9볷F����,�We�$��$v�,K=��_����nc(�����!^��E�þWm�+jq3�ďN3%I�W<��Q滁ڗK�����1�$!6m�j�ߜ��9�E|�2��'oy��u��[�h��S�F�m�o�=��ŀ~���_��{!���_<��\��]�?L��)R�v��KK����T>2���7]�)݂5�^�\N3�Q8�z��t�s��5�^UZ�w`&"'�J�%��7�1��&@&1��
�i|�y5��G��T���댐�~H*��h�� 2��R���@��.կ��W����m�l�?��s�9-�4��Zn>)i���]�����Ͳ�˧�/g����j�n��_i��IM"4p#�>���1hZ/z����i�ҫ|�o�Y�]�o��;��KSMzh������5��<�'�|e��s��J4�a>�R�nL���<�l�����}�Ĭu����z�m4@���B�:�*7K"�n�T������Ŷe�����uR�6�(�����,	Ǧ��*�>̕Њs���\vq�_�2�n�-#�m��"6��u|,{�t��&�Ӡl`Ps����䚡G�f����;i@�n�^*`�o��|��9�˔�׈�L��Y�K��ߚw��VR��׆"=�$=���9�V��+\x���3�w��9��#���~ ��Q��5r�n\�O��Q-�$�1�B��R��Q���X~(Y0L��� k�Q�Ø������R���?�{��E�J<G��Ĳ;?Y�ł�(=�#"b��?�q��#�D.w3�t����L��JsB����wN��/�����T��,_�����f~�� w%��}�=�p����5�d<�GŶ�״���!��~.�=����+��^�k§WFle7�+�$�D�5�M#�2x����:�4@���6�:YSޫ%�����u{���g>���6�#�w���L�S��������v�1o:���*oR�%�m�ҹ�/��8:Sy��]x�|d��C7���璘8T��x��{�T�ggx]�nt=�`�5H����%Z�\��}��z�<z�Y�Q��T���>����Y�B�/r��m��a�]�^v�."ף] �~���@�Y�_�᛺�P �N�`aթ�"��-���n�9�T�[���hw5�Z��K��O�ĸBO.�fFϜB$����^����禗�S$g�_j��'��Q���A��{{�;�U��8
���	��Ι�����#w���qK�pb�|�i�y�*Yx�� t��J�$����H+$[�=�@{]TI%������R��WG����/�;x.:T<�����h��@bY��;[ˑa����3��ou�Z,v<�xn,H��ir���鱞B���Wu���ɪZ�f�ٹ���a%�-�Σ	�8�1��{�;]l8O�[~C���(� �N�'��R::De��\�Lܧ������ߥ=�_�lff�5�����N�&�~e�?|g��B������:��bM1���Wm��A8�#��X�� ����a=R>��P'�Y�%��oP6�[2��s�tW�᥊�&4����Y�wø"�98����lu�dr���L��wǖ����Kŭ�|X-��r�һK:��9�-v�V�5]6@����ZǉLe5��A�O� �����V�އ�E�r���.�@��ޑ�a0hT��� 93�/��qkc�EaPØ�/���>�F��^��Yɠ��J����)k���E�`��Ps����{Э�ݢ�(ΊU1GО�k]��1-�e��1۬�`�A4��o��=�w̂	�9�A+��#v��w�w�H1��h����MR�~iCN�D��Y�,�����d���<�UJ�J�>n�#PO�s���Y�̆���`�7z�,�Pگ�4��!��&}�/>����}P<,qh|s�ۆT���q ��-��#Mnk�K��$����\�g�ж����X��ݸ�\�ԍ|��#{�@�kՖ�{s�ӡ��'��H�ȋ��A!3��Zv�����nAQޯ���wt;YSE	�����O���jE������NV�JDͥu��.p���E�� ��<��A�J�_j��'a��F�̩��k̹�F�^�_s�R\Y�~Z��Fb� �ÿ�'�H�����V��?�dOĤO�1��$ ;��/PFl�B�N����G]a���i��G)U�<��\Ԇ������CO��G��g��Ϗ$np��JC!8�t��g������ǃ~�
��n�fx���X����gݺ�»���9������A�oJ�#��,�p�=����͙U�2r@���pּۧ��<��yͧI3�� �@=�N�?f\��!w�b�ǫ>$c��ZR�S�G�y�X���y��Ø�E(�S���{��i�/���������5�l�G�&�y#�2���֛͎eϾ�k��V��*�ݗ�m���v�\���ywBH���K�|qgҳ=��4/�|�ʲ�_҆v�D^� t�G699��c7UD����R��4Zu�pھ׀0g.'�J������KǴ���[�m4���#]A'��C�*�/eC��OK"52׀��|��3W-Ƞ`Ğ��e�fG9�����������������g�!N�Ú�A�J�]'���<�z���Rh�>�O&�{�P���c���
��Í78i��+T@9��4G�zUB���l���3�pb�M^�h~�4�/u>�_��;/E�:L���Y�½"�����7]�`���el��"dN�=��b��\ښ�%�ȿh��x
+_)�ײ훤{�@2%��;�"���'�Xg"��� ��e�'/�N��k{I��7��99�\ʣ�枂��l�^pF�$�`�9������,���ov'��/�&H���@�'+�,�6ZH�I�_�UP�r#M�,�3����&�J�rCf&�T��me��j��;a$@��3�Bt��v���C9�Pz�>!��|����)v�h��ؿ��^�~74/h�˓�&K	N./�%��9�8��j�zB�w��Ѩ�	Y��s"�k���ewB��M ko �u�R�/�����e�m0�<f%��O��˥�N�v��*=�c�%�v�zůX����M��+
s�wZ��]���*�*��_]�׀��Jßo=��jDM��3C�@!���A�L�A�^\LJ��N�C�5���M��[����X5w��r��5t���[}!$��qXk*�G��{�w���7xRZ�2��¾�EeICW}���EԴ�:��7w�_3��ؕ��~H��y~"�&��	�b=O希�N�8�TJ|�G��)|j^�3��I_q�����8\��<i��]���Q��ċ�cf�$'-|���{Q�����n
R�&Ψ��<���v!M�w��q(-����ۗz|��3���W�?Oj�����Q8�,'ޅ�GW���M=�3�A�����G/_=���&�h�wgJ��k	�t���Q�Ŕ���)�o�?Fg#/0�ڲZ����9��U'�B����؅�IF�$�Mʪ'X2���U@4�\��c@:T�E�?�>{�n!Z���X+�4uq+p��b��mQ#���-u�B��6ݺ�"t��Q�M����/'�xa��;��+ˏk@��3��^�(X�k�|���7��S��H���t/��\&�4�3GqnxwMi��Ta�L��ya�Ը/�܈-�> �(o�-�N9	�`�i��2&��2�G~�s��XLI�_IN,6*��n8v��g�C/x�S��{w����R2���R���M����S�[��T���*�`bMܘ`z�s��t,dkYV�aߣ�����J��#� �:n})L�q�7,vF,��l��Ag_7d���i���m�������9�y��+�:ɣ�P�����_����L�F?�1޼1ނh��z1'��xmTCx���c�B�ֺӎ���hSRP��k@�֬�'̼BW� �u����o��z.eyk��y�|���3�1�r��:�&t�ؼZ��c�[�-p	�j(���]���UC��|A���N����.�@��T'��"]�� �s���e��nȜ��Q�]��`�Ի%����̏����[GܻU瓯�0�IVxS��V��oӋ1X������I��\���.�!�$���F6��8���ҭ]��xV{�g��Y�c���GC�3sD�q�B���M� ��	|3_�ǌgY�:YO����f�B���ሊ4ğ�-��m�����~�R�Q�;��I7�%�����Q|`I�z�lb��I�w���"G�O�}ڮK@��W�.�3)xy��g��!�l
�r|쪟Q�d3�$��D9���R�V��T�a�,��R�&%��V�bt�Gw��>��O�`�@KU>O�b��Ṳ:��7���m�V�e�.s�J`�xY��*�����J�D��`���O�;H��MI����ts�c���,u�k����f/��Kl�6��U*�vx���Ϟk��e��T���⽣����k�F򥿁*���I�L�����v�(,`�O髖3}ȧ���k�������b��w���vd=�������<�"P30��٤�W����'��*�]��py����;3
m��]���_�O=��q[�m������١��]�Aw�<k��N�.�Zg�Q?CVY�0��$u����n��śIx ��Ej�)A��p�~)P�]�|B�"l���tYcϫ�GsB�=��:My�@����,��&~Ts�z>`�U#�J�n�� P�3n�ݒ_MR�?A�~���e~�)�6&\�	>}\_tV��(i۞8�b��'��?��_��!�S�ߜS�=���fXSҫ23�6��{os�F��[<�j͂��|Ȩ�b�g�,6�i3`K���ԡ��5��la��V���� ��~m���A�q��o!����z��Z�e��n.�O�՟U��|h�Eͅ{��H��V�cO�L0	���n��b���WL�c=��[I��Z�޾h'x�-c/J�Zn��;�<Yˑ��	T�[����U�ϧ����g�W�y]�������ؚ�E�}-��Lae�6PX���)�,�pq�-�6p�G��tQ����҈&ݗi��$�߂%�V>[8������B*����-D|��_�.;���d����~RG�����sZ�ye��*��1^Ŏ��͠=P�jj��@��zu����Dѻ���{��������Q�A@�W�m���E�4)�	�����s)���,�n�b��~�������Μ�5`���I);��^|<i5.U�,b�C6{~��X��Ta�1@
¥���,J���k�n����vE�����ƿ��~�{����5Z���7y,�u:,%��5^+�w���4
��{R�.ק��-��K}=��|\I#�D���5�i�V�?VU/�4U�ZEU��D0���Uڡ�B~��F�hk����ݏ���P�8V�u���t�S��K�`Tk~����L�%b����օCUW�?GZ��Nߤ7���Ũ���O���)�P�G��w�ѧ���|�\Y!S��6�-��m��3w�r��o�*���׫n{Un�)d�מ�W4�X���W9>�"q�T������`�V�\�蓬������Z�l=eʖ��r�w�qd�OJ�>��,}w��2��(�W��N�Ce<��Uz��#/���Y�eb��z�Rt/�|Wj�?�#ݫ;��;;� ��
��k ���M ��ӟ��)~ʭ#�2u��$	@F���?��-#�/������a$
 _�6��Ϗ���E+�>����J��;Ww����A1v����q'��{]=5��~��R�6�=2�9�ˣ�Ų�Zy��k��xE,2���$ձSPm�Q�|���[�-\���u1�Ƹ�ֽV��5 �y�l/���R�l��5��PʑЎ�klt����@�_x�m+�4
���gDy����5��	B��|���:��+��c�c%�FӶ�c�/�J������l5�n��A�%u�8��=^����E�vįE�bx�����-5R[���C���
xyZX��%L)s�=�)1�,Lg�^H�pe��n���L���_W=���J&������ܓ��ϕ�w%Б.�a�U����_	�-~�U#��@�4����A3e�@�� ���^��,���#y7���fjGH�!V��R|0���.��g�FN?2��i�w�U���ȍr�1�k��]���ڴe�FBn}�]E6�N5z��mB�tԸ�B�4�&��Xor���r"p��*-5L�_uS�𺓅���#�L>ts2���%m�>rbM���8Lu����烜�(_9�\�aa�p��ULQ��a�W�F3�ʓ���<Ļ�ҘI?G����A��.��i�0ժ��m�j�nd8�b�l��.}�wM�ߓ{���vdor��vBC�p�CqyAZd��=��%v���0&�~��!TE��e����[�7���9�<�j�
0������K��k�P��VU���iN����n�eE����yn�
��r�e��-(���Q��|��ֈ�2�+xr�zX�s�?��2K����N���Kڎ��N��1�J�(�@�� �[ӆ�D���_Y<�ZW^5 Z�η�{���3�DU���9�WE������c�_�������a+��-��:aȚN���H�5�]ShF%X�A!�n���~�w�����N$��R"(�L_ԇU����r�fx*.>��Ԛ'�l(;����њkU�]C؜��X����3��_YHqq�3��5�JU?���_��0�� c�M�|U�vV���a]�\T��2��K�BR7�)�]K�h��`���_�5�+j�E�^ܞ�W�a�C�|�Ak0��}9�)�]�R�+;�d�������j�F�]���H�3����P�]95���J�/(�f�W�C]����94�d�C��*� {=��n
&� w��ם�`�� K 5����sɛ\��ؽ��`D�����]�&쿥<��#Jc�N&��e�IJq��'&5jx�1� R����h���Cb[�.A5�����U�uI��J��u����C;�t��9}�������Z�њ,P�/��,����7"�>�㳚E��M:s�fO�hU�b�x���Ч^w��9^d���ފT���K����X�`D9��)�p�<)�z54٠�l�a��G�)u�@r�h�V=���iʬf�v?Ѣ4J�WOh��u(�����[m��o���n��.k��5p_4<�2����$xO�F���;�١|��Tg�~Auъ�{-4�O���{�Ib��"5q��Z�A�Zk��cK�תE��3Om;�Z�1�]=^�}V�9,��e��Tg+#:Z-��bR!�o˖Ą�M��шz"[~/I������X4��*[(P�p�����m���܏�Gt��O�]�z��pŊ��ޜ�s)�ϯe�憭� H��8ł.	-˕:q�`��7
�E��G�ߐ���ܷ�����eb��q�7��R��Iۃ+3U�Km��l���$i0�s?�L|Y���cQh�+j���L�$�F ���]��毒�h!էs|���W���(cn��u�>�����:3.[9�6�|�
ǃMqװ-�ޜ��LPE���Ė%F_E͙�gm&G�nS�K�8Uc��;=8��/����~<��2y}�+���P�lpꃶ�Qs��9sڋ+�nAi�ඡ�[�jw����o�\�bU�=��3�(��ʹ��F����� I�p�����M���x��������IM"L�
^ÎR�1"z!Q��d�bU�;�����k
��L��r�-Zm���j_N��\FNwڛ	/]��nx��Z�f�����<���[�46~*{���c1a�1p�6i ګn����q����7+�%������r��M�jK������ `ԕ�0�U�����A��M�h�c������^�@��7p��}C�'Ve]��;*����a�T�M@���n(wBe�d��r��;�H�]��j�53=�k�u��3���^��n8���+A�>�,&����h���I*O2�_�>�Q%���.c]�����;0��t&NB����و���+tX�CWy.�q-��>!ZB��/w����%R���7�\��K1)񵘶�H6�y`����o����2sD�v
B5�]!��%�p����*�t/�-|@���b'�O��*=��2n��U�JV+{�AbH��/WE١��vV_��n�0�y006�y�h��������s>�>g6����li����I�x�p�����0O���n��������$�cm�		�v{�	0�(I����/Q�b���+<����P��v��3�����l�Oa����>��c�H� b��pn��B
�T�<��wA� mF��'�m��6�Z���l�h��Ho^*�fu���y(���e�O�Mu�P���&|����kec�etˈ���f\����Rk�C��y�=ԋ}��ζ�P�
X9����\����̄�'\&K���%6CL!���j�+r�A�2��{u��A����ϘntS���y:��.�R;U���Vy�,��Q�s,�^�FU�DPۅ�7z�~���b�O�⩒J�Z�o?u%h.�ܙ*�2$
x��`���IL{�m-�L��i<���;tA���TL�_r'��h���Y>�N��-���lW�gS�a��6��4���di�YE�cX
ڑ�I|Ɍ*&
3�-HF`�fs��������/��O����,3�,?�̶�r�o���I����[���M	�3�*�4����2V��?� ֚�O7U�ťS.���Mp���׀θ��|���;�S�7,�K�o=&��D%�R�}��Z�r ��<bsJ��@M{����a�C�;[QU'JZ-�4Ѡ��2�e3��W��K_�G��vD��R��g<����}m7�.k�oǒ̽Q��4��<��]R��RO��$Ǫ��
���G���~�\O"oR�[_�p�L�?����vf�ʊ@�rQߔv���V,����a��b���4}�/���<?����m�`����I�~;�׍qBK~�+�6��.��7Qqނ�o0��$�<���0�DN]K�|:�S�i_g��{����޷M	l�{m�5�zx�VG[\ބ�Ύ��_�JT�p��,"h#�s�[:�pL�O���ΡA <e� ����	L�/�9nccdw�\�8�̻����ms{j�\�����_LIJ4ѬZ���a)S�bE��ӫ!�;mO�E�0z�j"�S��tx�kۇ�1c6?�)�TD�Z�v�9g!�Z�]��0z �gi��
]<`��>Ê?�ɽ1G��@�wZ�Ɏk�OW���j��^��W�LW�oqڮCb��V����y��xsq,�+b�S��m���mg#�iR4����fY����� ����/�,����U/,��A'[��V���b�A��I�"ꕔ��2?^zu�Ջv�4;��ٔ2(M�d#"M�j�H����opi�E?jra0�y�X��԰_��oG����I3ڰ�՝�>&��0��������l�����X-'z�������W�AR7��s�$4DF*�������
���r����O��5�`,�|��a07K#�O/��8d9>E&8*���w��2��?}�_���o�yu޵����mL���/Mɉ����I"�7��~>������w�J�/
���>����#���=KX��FOH�_���@��a`�����z��9���T�N����KK*lj�Ҡ���M�_��K�=q�,������[
��n;m�EZ��_t����w�N5��j-���+Z�E�C	im�� ����-c�����
.�;?�Y���A�<%B:�y�Gy�٫�@����N��j[�:��Pj�\֖���=�_��/I��#�ش���5��J�oe�0��W���i�+���T*˙�-���Q�&�3^��U���[.����<h^HP��.R�Y�H��
�wJU17v>�~kRk�{1�Z��E܍?�38+��!�u�]�:X^��UGd��'ﮐ|I���+�1q5j��_��4�tyo�+��F�cލ����)�n�5�"�t�F�	M����1"���H��Nn�MgQi����<��M�1H/�t�|��'��;i
tG�,_���0����.�����A`�?��k|[6��v���q@(&���d�����3,}V�zl��U[�xW�%��bn������������}�)�����cWCH�Y��z�M���?�R>�i�sټcC�~�I�� ���9��F	�mڸ�H���=��_�t1~�_Ł ���4��H� \��YO���>������͗���>3��T�L	�� 8QD�榡
��GU�����>s�5�i|8�����m�{��k�Sd\B������Q����l��y���c��F3E��c4j$�����݊�׀/GZ�4хSi�y�%#Rl�A
����L�*�C,˾���5����}�iR��z�<�P�9��g�oa�nِ���l&��Z�՗�`���@f~�G��o�sdJ>�x�N���t�M�k ����.�ٜ�۹ <h��]x�N]�k䳉`fe���G	P���,�I	V�]�L�M�NQ�{���<����çE�[e=-U�B;�MQ��e��ŝ	@��T��r{״Ǧ�Q��U��LOY�޾<�K�D}��'����;]J����%�pB��;��ܽ�(�"6�d��2��-/�c��Õ��J�0��-���h�l/9~Us�=���W��.�d4�j���*&k�i��k�s v���DEQ9��x棅o�r��6��5��7��}����LB��v�"�$W�W�~H��rb��`}�h�h�.��^��Zg0� �������v�+Mr�{�;9�r�!&��E}Iv��yq)�w���L�tx?��{��W[��+�������xd�����\�O� x�ՙ��R�'*�tg>���n��C���2Dm�W٪�"�R#YpD<���pE7�Os��;���.�o�(_�߾����=����}�I`z{k#V<7�Ȁ:䋤�YS�ƹK��o��S���4͂x�����dG�cYc�롪����أDɎX-���~m��[�D���ݰ;�ӫܡ��~�垎+�&�*Fz<��.��4���U��z����6ب�]�Ŗ|���j�8�[�,���M�_"�~Z}�Ռ�:*��~�=~�ɾmbv�2WA��r��lW�h4��C��ޗ�+<��m�ؓ,$���$����L9OK!k����Zڍ/N@ح+H�F`f&��گ�Q�̻ݴ��GP��~�9� ��TO�j��+3<����%6@w�F���:���u�ϒ	�@�#]7�*{X�o�E
ig6@��5�J�8Ƶ�~�&����m�әQ-��#����\W��l���l����&b ��7|�?�x�F�sa��+��>�H�[���!	1�(��_G1��Ѫ��_N��׍� �C��������On(S=����t�%�׋2KB�vEҁ�]���ѴTfz�|�ׅING�$ ?���^QM8Q�h+���GQz(�.�$@(�	!�бћ����=R� ��H�- � Az���p��}�o��]��^kgΙ9g�Ys�p����~I��O�%5+�Jzt��<�9������*܂߬��bW�V�9�޴f����FB�=�]�,�8V4�	�����{���Le�M�����v!��X?z���� ��&pU�Ŵܱ9�~�>,�yp3�pZ���ȇ�b�ɷ�XNt�HdZ�����9��b�$c�C�����{`���/��6�OSޖ�<#���|����
�'6@U^�YƬ~� �ԃ2�9��+9 �>U��7j��b�BJ鼁�_Ƭ�>=��2�ǿT��O�vWi�}��r�ƞg<�k���iº���!t�I��2��Ӕ��;��/���!Q�p㼞A���kj�`cb��j+YR,�a���Q;���4�UA��U��N ������*Q�/���b	E���b���'�FBu�ؙ���u��Ap���I�t�/���i����=>�w�T����m��%/7�[�m���:��z�=�t;<�v3��~,���n�y����d_ �?��5��Ǚw �l��g~������|e��E��m�I�[��BʑP�@��O�������|��k<��Dy�ç�nw9ge)����DQ��Vo���̽xՠ^Me���M-s]��ԙ�6-�N�]/�G*U�<̘���e	2���m�{K8��nL����2g������5m��\�����UɇE���k'���YS�T:�7��.��&0G��xr��iN��#u��.8<Θ\D!���|�ˏ�M`�[�0ߍ�lZC��G�Q����",bO�:Zya�O^���jݻ���Hg3�����A���hWe b���� ˆc������s�>��:V�Y����P�]6�ޱn��kuT<��������4󗨅ü���'{W�^N���d�
�\�Z1�8��n0�-�R��IEf�h! V��BS�8��X�Y�~��=K�U�"�X$�H�S4��kT/mVTp�H+�"em��JՅ7�x��@~7��æ�8\y��Ɋ��r�������3�Ғ�Z�:�������f�\\Ȍ��?�������Ջ���u⭺q�&ŭU)!�^w��)�9\(W;>���7���mA����s&�'u��|�#|�y�w�~^d��H�	6���X~}�6����2�!��5�0>ܨE�\����(J�U{z��m�g�%��~����у��?���WmS�@��������o��=� В�%kxO�Q%E��gW���y���;I�
�gC$�
&�
!���yU��"�	
���C�����c�t�k�Z7{����{{�'�E��UQ�����V.?��e����Q�}���y�
_*rR@��F�(�6O֭(��f���y��jp��g��\_Z,��;�kV��Z����q
M�:�-A�ٌ��3���.�r�EO~����O['���uNϴ���a6�&·� 7�͓5���5w;�re_nmd0���	���ٜ��{p�)B�⨎�ǯ
��S�T�\���{��-v6� '���EWPW��u�?���l�YFU��Mt�n{��{Jl��Ϛ�Լ���6����T���.�O��H#0��U	SMCBD�rݳRé$�xYӹJ���	� s-�Mx?��#��p��F��VaɻQ(8hzQ��0��N�	�w�'9k5���P��@�  M�����[G��	"S��f�V����%�)�6��!�aȋ�٫uᗪ{��q����j��~�����?-��SN|>~��W�J�d6\\ߔ{��l�:J?W��F��۾��c�>����������EnN�-�!�C@Y\ͭ�e4�CT\�g��p��*Oʾ�	9R�F���#��#�u�!����$B�;[��{/�j,k�{;��mG:�ˁfQ�B��Җ��4K�/�8\��Z��P��<�P+�G���U��������+���4K�y&̓�j���h��yc/ ���u��K�х�+��ǟ��U+wb"I�>7u��3���O��F0�ߚ�\_e
;ǝ#J+E!L:將Ͽa���g�;���9Y�0�4\E,���R������=�"�Tey�x��A�6��ʅJH��mT�]h]�H#��@��ݛ�PA��$0� $�p�v�8ʺ�n��/�?Ffć�����ʇۅoE��X׽(�	�����/!���K�d&�B��*�%���3���}��z4���Go�+2�Nՠ�F�Gnm�B-I�:������|]0�Td�:���*��Wy��U�s�l�-(U�^r����V����z�#Rq��Ӌ��Z9
�G�Z�����N@$��R����^%y�0�wW�1OC`�б�4����J�:������rkk��ײK��v����,}/eoz���;���Q�0`#�q��\���"�o|��t��"p�هG���0�������t�p>�a7����H�H.�*��z��@��s$'����L3�o�m�î&E+ԩd�nz�n���{�al̕�gl��������Bt����R�W|�7}��mMo�g�K��U�Ck�-����)����8���+/C$��_Z�8�~S���$�5@�1����Z�Z@�Gʏ�;�1 Q1�t��o8���n�YC-j="���J���&�Flwt/6FN����c��(?N!�����g���׏_��=Ù|��Xh���H�	�n�w�����<Sk�sG�I<��z��|�9Ϛ޺}��W�{ÞM��%g���j����;��D;�
v[��Igٜ�O��a��� ���{��F��Y�}�D�;ږZ 5�}T�ޣ��F�>1��KYp��X;֑&̀~�*��mw�=P���VPڊl([����� �����A�g$���uU���*Vs4����>���D���Yk�&�׶׆���a ����-��. ���ꕵ
4�C]ڧ�3�$�3n)�8.<�N'���+XV�:�Q��ʀI�Ɖ�zM8gs��M�s�wf^����$������H02�~,����|���ШC��V���=�~]��.מ��N(K�
���!8�~���יmn�u;?�k��a�a�����lWbR��n�ϯ N���Ԍ���?��FZFV��ן�Wk2?w��/�R�'GA��N�&|\,2jA�)rqaQ����R=I[�4�	%�ktQ{y���ߑfM!s�=��G�,. iQ����eMh�+�!�MQѯm��F[�zxnć��ܜ���_����r��:Й��bp��e��X{m�/!$�1���[�I���e�[@2r�#l�{�1�~�(v;��Z���ʥd.�C�/�xôݼ�����T��_���f�n�%�nN��r3����k����)P�k��F��-��B���35W��o�����ǾO��8BWr���	�3dM�*�_�xܡ�r[�n-��ت�!����tb�>IE�i����}%�u];޺�@^i��S��_�S?!�n�<u�_��#W\#��-MC�3��#"��-�]�`=ͥ�ק�]e�� �#wo$��}�Pv�7�U�c�瀔#�r��x,G��ñ�"�-v�s��3\0��P�N�y����+�D��/ꉨ��	a��KڌmI��xC>{gz�;+�f�z�9����ޓ��ի}�<��\�OE"����Y�������+#ͧC�1C������U�����J��Uӫ̠�t�:�u�7���w��q��g����Z��'�g5���R�k����C���韖�~���>yh�$�a#.K+k�:	<k�@}&����?c(���t�w6�%�[��~!�x�K+o�������W5����,з�v�l�C�����TJ��9!��M��O�����Qb;� �M�^�����pq��$t�Yv�p,<�l[�|�}2��hw�P@x���#��]�U�`N:f��.�mҧ*����ؖ��r�X�-ް��C��96vЧ�`��`}�z�u�j���x��%��~��o��̬!�iN�{�a/a�a<����VPq�2���+��cʒ�t����������a�;�
��[�����g�W�ޙ^���L:�s�) ��"n�z�u��*;��������)��G(�o� 7��E?H�CXx���y�[�ٳ1��	Y��w�=<�M��Z f��]h)̢����%��xԯ�����ϱ��/KX���V{�����P�����	O{��rJ���*�b�iO�|�s�_��h��-�b�D����E u��Yub�b��p(=7ȸ�x��_z8���7nŐ��c��Vo�m��=Vɥ��]i���Q� Z�~�Lآ��z�����3( Wx:ϭ
i1�I����\ʧ���#w�D}2&<Nk��dv@�A�I��]����E�V���Rk���$�a�*S��;K�"�n5d��~��Л��5����n
6n{%!�yi]y���Pu׆�IĜ,�zb����L�!�tE�][3������<6����8f�����~wVga�98vd�Z�wzX���@&����m��\P��6	g��PՊ��O.�ߕ�]�<�US�)��ߛ�
�&A��:��sNs�V#Q:�Dc�R�S~B�i�-V�D� ��z�z�oa��ǝI�9�V��EID�w�&�����1,P2��W.�z���$��b�4:���B�Ƥ�D*�HS�i��������$1ݚ)~�r���`R�"2������'V͋������,�{?��Q�-��=v]��*�.��B�k���|�a�w#�����N�����d;X��-�ك�S����BT�x�岨j�u��<(ɳ���sfu5�Ɣ��o����4|�q�a�����x�5qN5I��&�� "nM������BY/ {#A������wg��%I��a�/��Ow�b��r2Uw���h��@�ߤf����$g�(���~�J"Å�����y�����y:i>�q?�B�����X⒑G*���`�mԮ)i���-˳5[�k�8��o���88�	lq8ͬ�3w�Q=����aɷ��w;�S�7��/�N��y��=]o6�S���'eB(����`�&m�]��?*�������3:����2�=���9��� ><��{��V� C�|���渑�o|�]���2���*�=����� ۭ+�T�p_n���*�ߕ�3ua�$���c�Y��}�B�RoZ�W���E��c
G�i`Z��ǻ�wif�[��:�k˛���?�<dS�Op�_���t8������(�T�V#��߫���iG�o��9]`5cs@%DjT����Z;�_�����3�������'���o9C�R�*C������~eV9�iL ����hV����՗Qw��&
�!Jy`W)C8��Ø?�n=����R��K��pIj���W����0z��*���!rSl�0�;o%>eڲ�[-�Q��ДV�:R���][^�|�Os�c�� �U�F~�U�y�o�~v6O�Q}9�Ϊ	U*�)���MZnV�W<�R��U��q��~RJ�Z���.6D8E�Dj��i�����Kp�
p����[r�G�[�����.%�#WV�q�ZAӺ�e7�ݦ@s^�t���
���3h;�Єt}DY��j�H���s@��~v��ޡ�r�����L�H�mb���x5l�(`��ޛ�lW>NLF��2�dYI�ܐ�]�{��7
Ir�������u��Tޢ���mەSRz*c���,�]C=���]�����C[?����2��$���u1�:����(Q��~���.�ր�������c�[G��W܊-�.��ő�]�b�78����������ӱ�����0��s�GO�Mr�.�Y忔���˿�Z~�I���V�)�����n��d�]R7�z�2!��+U���^eR`T��43���|��H��Ѐ��0؟?�޼�w��޲�5�!c���C�ł�/�C�>8�0!]��H<�,´\�p��1�L�S $L��
�^���`��Lo_�C�[ޞ��@�ːf����/{�7o�-�<�j0I�3�ĩ�ڡ�?��3� l{��<"}��|ǚU=�H���3\.�Dh����7��E���@0��o����~k��G�ԧ��g_t�z��-��PY��V--���{3aׁ���5Q�.op�[�"�G.����p>�%��	��� ��,��؅�{���b�ths���*lE�F�+�ͯK2YI�d�!{5������ڃ�;�?H�G�+�G/���D�Vo-����A<U�$�`n����)ʻKȣ�����(r���|T=)赢���%t Ձ���f��tc뱀���}�� ��G�%��$Mg
�]?.�c�Fĥ���_��ܭ(w׃��d�0��-��[<�^�= �-�|m�,t���^�E1� ����kͣ��p;љֻ`��i,�H��t3W�R�f�IN�Ȭ�;A �X!@�?��]\N��1�\��g����i�|�sZ, �j�!�'�����ݿSt�Z�Q{~��8)�=8�������Χ��gιN�qi�V�<��b��JݼR^���R�B��]B$VٯD>��	5'P?��=��&�����]�OAz�{7��j0w}$D�����/:J1�P�
��ͷ�nӯP*	e�I_ʷ� ��

�,�I��μ�K���?���	t>������4p�	��������/�-��s�ח�-A������������]���X���m�k
��. QrLv'�d���dy��1���F�D�c��'�nng[tzV�-V��`	��x����z��dI����bxl�|x���ou]�y1��a�A
UAd�WI��,ݴ��S����P���n��@5��۩��h�a��ϟ�f8G���)����hTq<B����Yy�lQ@��U/%���	���Q�ߤ�i��e}����}�Y�o��t.:U��^���N[��*W�}�ͺ��^����[H����|z�ٞt���qUe�����	*·R_�5�fય���׮8���$�h/4k�ġ��M��-�	D�/�,��+�g!�I�ܒfsD ۙ��k1%�Y(Z�ߛ��6��aE7�i����D̔��{�7���3!u 1��a8�������c��:��I�+��bм��#��zS~#�sj���pg[r@'�`��W��d0�ɫ���+�Hǋ��ŝ��Q�f\�Z\�9���N��=ǉ��Lr�fת�7n���+A�p�Qpi�TP�|��G��X[[���������|�lX��)+班T`=9n�D���izV�Ҭ{�795�`�@� fRO��>W�p ��>G�G(\�C�}�!Bb�`!��̤FC3�V�;�j]+���>E��a%���5<����g�:��;�:�~��F�ŌPKgbO�]�I����1��
����ĉ#�Z����/}��4���wǜ���g�`��
^�f�<�ำ� R�ڬ� ����,UG[3�������*����8��(�~V�C��I��i�B�cV�k�L:c!��.�$�%���"�]w;���VǰWC6����N.��7b�
��6z)Q26H�`�ܝ�đ���S1��8���:��ݵ�B1=h���i��Z�}R	���K���v}]f�T���8}+*��,�ط�����@,�6�<�|��7��G�p�9���YRx�YɷƐO,��Y��������_��^���Ԣ~U�()�Oc0(i�h>G��F�U��kᕺ�7�lyl���ϨG��"Q�vl��>�����p��X��W�˯��?	���ܧ����p�^���ּ��gB������okqp���&Fj��^$[لT�<��|0mHQc����|uS��m������ "�����i���?~��]��;�<	�̥���y�mQ���_eX�a�^�����i��
i���rs���`�1� �&�.��`�ُ{�d�ƥ=T)SPi�u����}��&YU�'�im��א�Rm1���H��H�����]W��k�(t3j�NpmN��EN�c$�n�����y���ȑ@�C_|�Z�A�,��B��*5���3��4�泞�տ��4I�U--�I�[kU�v��<Vm^�ڮ"e(*9�)wfsg�e=�m�aS��[Wr2���d�8��*�'X<s��"��i��װ��%��أ��8�t�O�"�[���Q{�`S�G�23!�Pd5-{�
>/8; 8��G|Q9�I�ܟ�=,���A�/P�U���K�����o{���K�#�m�b0�$\������.���d�p�e�(�J�AyMiz�me�墓;�ǚw��� ��@�',�`�t����҅�M���=���v�������]K�1;Nkl��鋚�������1j����֬#[�5Q�Iי�Si++�XSU�0��Ln�_��0~5�zE�}|m�����}���MX���R���9K���c��RK����97��}#rG �߮-���A�˧u�x��N���$���M*5n�|f"o���OiȻQ�<ju�~k��$ٛ!#��q/�3�|:�U����'n�'d?�ì����A~����rN���r�}t-FU�9�!Fˁ����l��8:]��s������M�7u0������>��"1�>l_X31zt[�:Y�Q��5�ޗ��d�;!D���<��$޵d�#̙S⍣&g�q�W�u��L|��h�a��r;e�Qm����Q��a8I�&S¦�7��h��lte���a�\�+N�ĐVZ[�ū�
ǭQ<���vڠo�~�n�7+2��F���lZ(�}�$�Y?]6�Ь���ˉqH�I�R1�ƾ�&�zW�u� d��ֹ��5?BB[��t���o߆�M
x��[��,i`�d)�>q�,*��6q=m�`���|��yk��ϣ?G� �3� ��
M:���o�߂��Yg�/��+6<m@8~;������5M����cСz�}zg�o��g?���J��^��ׇ���ga�Ú��|�.v�%[���?zj����O����,�>�(K���I����	�8@���»��('��,">��Н�{�C��鯭�� dmBB��g��lZ���_i�����k��RD��+�R'��|��Mm��4ϵ:����&2ߤ���̦��x�L�ڝw�گ�s��˷�u�{c"76e�V-�\ W;l�����p6��y�"Do�`��<Y��F2����gf��ϰ�fW�fE0���7�s%y��ǨSlK���me�i܏� ^���d����f�ݯ>z;`~ �{4r(Yg@-�Ĵ���",�>��>�e��:����NZ�m{w}ȭЇ89�����P9�3�FN�%R����)�����@f���[�9�,�w��x�!�P�ڻ���3 �o���wqb����U��u�p�Y�6�A|5�ESkg6磏�ו��l����t�E�č\g�Y�y|�r�M���6P'v;Z?z�Id��4�Μ97nׁWs��vW�=�A2�s�aړ`�`X�.u}�]Y8�J��݁u�{*86�KT��(�+J6��~�d�������mD��( �>m������TD�v�LW��K��_S�pw Ň�;u�}�z��ކ{�������sa�	���Q��`�XSI�\)��67���Z6�-�κ�ꌠ-z��׶�mS���U�6�7v�2ֳ��W�����A�_���!?�/ �ek���ex��'��n,l�+�-$�v����)��/.�;��N�r�P4�ϟ�Y_���"i�/��lӓ�l3Q�d�O�e�:��m1r�	���W�O�o ��t�Z�_�6�9hk���,l�~^P�1F��?�m>�4��$���e�_(}�Pe�o�I����ȸk,>k���}o:�g�{�y¾��P�Te��!~�/v��|[̃p��e����p���6p�eN��z1�Lwd=X��q��b�q���jM��ѓu�����`k���c1qtp��R�L�+�Z���8G������E\�%��m�J�/����ȏ�R�)f�n�7ڬ��Q�w��LԈ�1#�$o��T��(R���Y�G�#W�-����>'Z�K���E~�����d�_	"
�r�O$5Tt�	4��!�W=�\��*����C�~��Զ���?���$�����$te�f��N���F����wX��D��֓ %S��5O�+�hF�,��,',��;�BG&0���J?TE&6%��\A��}�Jj�+-�7�CK�ĽCU�S�ؽH���r�v ���eg?�M-�R}X~���J��c�&�E��%�MU#�[H���\F���L��:w�K���ּ��cL{a�t�K�K!���J��q��P�Ǫ���o�����}\��v�O�d��6�$�t���> 	�����Y�1��o�������G��Q�@5_���a�F�6L�ϴD|��ȝ�⑙u�]�����vf)|t�����5�]��Vdl���$��+��9sd�	�,����z���ӐP����>/��n��&ٿz�T�e�7uj��\=֩)��*:a�n���$��n/�@ ���k':���T.� 8�K+�Vd�1�kh�����vӵ��K�6C/lj#/?�ץ��LWLȗձ���/A��JԺD&R�C��|����v��D~�6�<�	�����Fw���ӄ�$TX�J�$��7���]��^�
��+@[�����n���_���'�;�k(�{���u�3cWʳȢ>�r9�����R?f�f���?&oQ�Vc��9�"z�Q�?���ˡ�r��K�v<{�*�n�
LX����Y����"A��9�Y4:���%�{�/ ���
>+.M�7�^��B:���p_FQj�t�np���M���~���+$"=1�T�-�i%4�/��p�~���n:5�.ږ�5��(0�/�7��-#��?9���Н�m��'��"zx=���L��F{6r
cs���/\��K�� �K�x[8�F=3��K ��7-���g�*L�7�����c.�`������Oh���<�+�q�~�m��$L�c[��ʅ�
� P��Ù�ĵ�wӛ��/]��M���a,������/e-^ST��7oZ��'G�bjo���K�TO+������f6Nn㜀��|㾸>a_�_����5L��xu�o�z&���V ���x�k�d��Mj1������n.�b�Ѳ	��?�TV������d�-[.�$|�(���f�Ic]����HK��Z��am�-��64�$��n����4�R~�6F�Z8aΆ^st����F�4�_����ç�?ǢR+�EV�d&4�d��-!����2����!�ޤ����+p��+�} ݤ}���^���v(#�-�X�H����[��Bx�*�	��<58���5�zL�ח-ٓ%Hj�h�B%1 	B���N��ӯ4��_{��"��&N�oMpq?��V�����m@��W�_a��>3�ϻ $E��I���-�\9�V9$�Ds�5V¿�ܔB��yyVV����;��w�Q.*:�c���{jI�b����f�_)O�D�*�7�~�!YP�#I�0b#�2��Vw�kN��*ɻ97�~{��9�K�I�i1F�S:��u�3����B��K�羵��5���$8o����Z��-�]��͐2nI��¾ow��l���� x���mYOa@زIDx��hʂA�h�#�t�w;A�s���2��N���{"��G֮:OB!�+�����FN��^�ǣ]8�Fە�V�����G��K�����g���x虼Cu%��?6>4 �Va���*G\�ӝb�`�/��8Y�I�"bs��T�2��3
zۓ����$wͥ���iO��-���N!��
��c'=�l�g��)i����с�G�K~�S�X��nt�w��W���bcZa����J > e�������VMU�DԷ�X���w}+=�r�^ƭ��g�rE6=b�<�y��T팸`~�D�a��D���ӲKd[��`=o�|ٝ{'����/�}�����Vt�"ZtpX����,���G��t��s]�Y�Vi �\_�6�>���4z�;̆��{�>����=]6����<����E�Vzq*�
��yw��H���T`�W���x��KX�A�&��zc\Y�HqdS����h��[�Bd´�)X;d�'	d�O��l��0H�|�ݚ�Q�}I���I�]�1��C�3	#�L��UUv�.�I����ض����� RRt�,����´�$��-em���m��v,�.�(������U׀|�^�R)�0�0�uZ�[�2��|�p�m[#�����٪:��6U��Ё�oc�\�c ��?*��3�S��^=�^ʜ��Q�g�9�V�.Q����N��q��3���Q`����k`A|��●riuO�����o��*�T�Z�{���TN��������18��_��I�[�����<��(��r���N�#k�������2Q�����"
;�h<��W���Y��5NP�}kB���ݳ>e~��UFB���&����Zl�I�1�Җ���}��m)z�?�[���M�oI	����V�s��ˎ}��F�B��]�9��`qi`Ξ��VHl�/?��
Έ���ʰ��%�s��
;���UȐ���99��.�I����>L0�����H����ªE�4�~�D�z"�<������v�8��-U+�Va�$�ۭM�`��ޤ��ns�+<n��WEE'9��4/��O���һby\&۾�n��q�m��i�1c�����u��.�ػRHS0ȹ.,�+>�MtX�^3t�s.�DvR�'��8���4j[�����^z���)��G�O,͙��E��8�&���I o$C{9����q�I���L����^��{xQ^���8���r��,���\�=o]kD��SK�"�t��4�`e	Z�@1=�(|��A���b�Wfb?��ul��߬�zӐ~6�Z>b}��)��k�O�>:��3��zmx�_��mZ�Gç��:���R�6����	�^5�2�L��p�Q���h�4�Q]Ɍ�~���c`�w��*z���\�A����g'�+�cewʱ�%F�@��1�=�e�s�ڡ-ZNn�n���'_=�L���5�s�*Y��7=��Gj;U���p�1K^��}P��t+�<C}����Wʍq�a�x��{w��/ae�dd�9����|�b�:bۄ���vZi�`L��K���HS�Y��#9���G:,������pg����\iL{a��C�i�@�/�E����$����RƑlyն���+���6yV�Ù�>��ϰI:|UW�\x]�p�o|-�=��#f7Z�_3qX=���hP���� ?���-��Zl��{�9³�v�
_}p�I�ֹh�F�n���������Oո7�!��y���!�$o��k9��Q	���_�\̑��_oh|U����F��Ȅ���Ҩ,�q�{���0Ku�X���4�k�u�����2n+��P������Yq��s�Z���Ʈ���l����'�H���+��l$6ǻ����
2���Z0ܜfivU��6ܿ�7Q�܊~���*��|cz�����> ��q�1(o8P��Z)9�3����C����S���`V�'i"��ݯ�|�+�}NpX,�g��"���ۄ\n��8�a����<��X?p%��U-�A%�(���obt��Th�Qea��5�n�{�q�Y-�2������4J����q{m'WB��Ȕ�h�g�N^��gJ�̮����Y�D��=ќ��S�y�kCP/0�p��v�I�5ktV�>�=>��Cp0�,�n�>r��a\2X94���x�^�j�k=��j���<i��8q��P2F�Me@��i��<3��
�-�eM���j޸��S�r�rs~iu�*WU�g}�Ѻ��JNK�&�������gx���"�<�9�Pu~/˽SqV�o~E�:ऴ&b�C�"��[�-֘^�(ԃWXW��5�HzT��OR
�FXs��<��Yx���ktKS���|��C�Z��������8�Up�к��C�K�)Bt_����� m�C����^a%ſ6`2o��*C����:}��("4I	���3���V��J7YY$� �@�B�`vy��Uh4Y�21l{��b�fB�ޅJQ�l4�SyEЯ����q97��}ᮁL@��-\Z�zۍ����
�4��HC�r�t�1��>f�0���U;��z\zSc-��N�֛�|8������B$�D��V����ǫoǯ����}.��7�;Wm\f�6g���K����9K@���<O�^9�.��x��]�9D°k+S���
<�c8m��~��#KQ�e^�V����*�B�����"���Т�ZD���ubU�c<�����xPS'�;ȭt�{<��$����~��:��s�a[�驃i�^'r�Ԙ��<t�2��n��!W^A߆}����/i���L�|t��8��4Y�#1Q��vN���uD?W>�Jx���!@:�.�-A��cz����g�C:�p��U�7�7�QLě2R��C�=�]���$Ag�W$b�3 b���3evX`���)�5�W�SPnޢ�?������WB����h�uj0�X�Q!��B��ҏ�R�V	��넦U���ʊT����{��6����":. �V�Rd��1���׍��)D�9�0ˣ2����HPS�.>ȜC��V���o4���Z2��d�t��oB	K�(�Io�˘�Cs�-t���BI����M��Y1F�0�Ƒ&���5���tA�'u$t���	�OzÙf��i$��)vM.9�1�u�S������@A����ٯ*!\�޷M��f�	���7��Vd:+?�� 1s���E��n#揼�J8mǸ�q���$�ڇ�?�7�׷�5 X���9y��6�5P��+˾ғ�������9���%5���-��G�tfRb`��0�ˉv��~6b��rj1	@wo�ou�e뽵M0h@ؖ���3�w5%�12�Z���x�K�O�2� s���8���Fԏ��y�]Y�[v�W�Uw%<���*4�O�G�q��z߆�u�7�{6��f�K���3B4�!W���c.=�{��!���q���Y�[� �/"����pu����^[��@�A�L��"�?/ͭo���:$��2�A����ۯ��O!rs�"�5Si_���p�Y�8cB��?]�8�N��e��:I�v���&�j��p��چ�爨#�-<KR��!J��Hw9. !��	�/��\~2�g� n�����Rb��ɻ�'j�*�Ի�C�z���|�AEE(6\<qv(�5�kvrs��?�uеh�	��ڋ,��ͻ�b�F'��������5\O�In�Y�猩p�����xy�{�}c�����`�g�6uoS�+1}��J��0�V��*�NI��	w2�Ty�.�aЏf˗���}�W?}DZ�.�e�@�5������ի�tåDb9t*���Xk�G�a�"�p��g���Ԛ�l���L�z�Zh�|0�f�~eVh���ڽ�>N9}���2�z��fb+B.{3�Ho�m�l��f���-^cˤ?:p&����M�Y;6b�y��]������Y���im�� /�������2e	5<ֳ���1���
���A�5R�[�/Eǖ��b��4:��M��$��po�2��7~�Ae���Oc��HsBt"�����V����X�7�k�q����۪�TWZ�{���C��[|w�I�	{3�}GЌ�&�?��&�F�Ȼf�un�|:�������;sp?��	!+̦�$g��:����������5w��HVj�t�ۮEq]���%Pq��:-w>�l�ηh�y� ���'d��:�x����{����
�:���� ���NjL��5bǌB~��	�����ߊ��0R<jI����Z���2\��`�$+���D��i؄���E������8��wջX���B��j�����9�Ώ��g<��pe픑��J�"�Y8T��%&�πv?����6N��a��3����]�"Q�j�V�u�W�Ñ�!�����Z���S-O�L��$��d�=L�MkGǭչ�������
j�F�]���QQ@�#%��Ez/	�O鄀�NT�Io�JI�����������	1�����{���|��z�3g朽�Zkf�>֢��0[2"f�ӭ�q��8P �/�}D6�ʈ�m�c��Q�
�e��Oq�{7F#Q���dO��V�v�6�]8�Y���ve��s�?�j�эg7�H1k�_橢��s͌W2< *��Rp'S���<c�Sm���R@Q�J�'���%��Ͳ��5?�Jm��@=�
f܄��kiJ�z
�p)j��;��++�-0~9��uJwO�8��A�hPTM�zl|�|]�/���9���>_*�����߻�Py�
,��빗��:oL^ܸVe��/>�`~Ъ��v�~O�����t��D��K�(GL�&�!5/�ۗ `��^���n�>2��� ���w#�8�T_,�V�/.���;ȿ�)���QZ�~\�����k��������	�/�8~ۿ����Z|)أ�T!���V^qSt��.��ż;�[�['�ťv@����<J��&}���%�%���ɼ��3��f
v�Hb����H���q=��蚁^�H�S/��d�K�Wfy5m�
J�9tS�U)��[�胝*��Hy�̩��<���+.�|Y�I0S���C6]ó���9{��I��vq�-8��']�:�g��Nmꁫ�o��m�Ѻ͕C���)-��A�X*p����2+��4Y����P��d�fxҽ�#�?�<?޺���h���,xN�&qb���X���$J�}�d*/�r͚�l3V�g�/l_��?mP�l9�2���I��C�����d^|�g*�$|�B���}��
4�M*Ѫ�b�F�T�C� h�����3S�L}���	��\�� �e�	3�AqKQjފ���\�
�
��Q^�3b�k�7u����(���/}.�w�����/H�|�$*�qK7�D��[H�R�_�/���ͧբS�,���m�7d�Ǿ���z��{��f�ԙ��p���9�&��İC���J_?0��a<���ߪ����.���K ʛ^im��ٝ��"��Zb��O{�K�Ƌ$//Gf#��)<�n�R���i\���lvZ��{fIN>�������T�T��vq5Vik>�'4������S߭���i�_�T� ��"��$�����}��:I��v=ۨy�ls��ų�vo�v�Cmp�$�x�.�d�9��K�9��ى����ey����һ?~��qb�zfq���rR�4ـ�L�Y��s@`�I��Sa�/s�%��v���[�x9p�R��1:����{jO��Q-3��A�[)?2w�����SUy,���^ݹq(כ@.�;�4�`&�Q�1�' ���u�)sF�K���٤�V���umS�VY�}�ܦ�����y�r�<�ڵ��F��_����N~C��� ���`jC_J�'�꫞�'.+�q��uq�8B->����B��VG4;�U�<�����ѽ%�cWd��O���.
������ڵ q�;�J)���V���i�;rq�1Nb~9�Cv	?�r,Vo�׭:�yȡ���f&Z�{�Ր�1"5�B�QN��\��<���O]3H�W;�M�LR�%��/--�v�9����F�=	�ewt����=���s$ت�=VP��#�w{�3����N�5ȃܺ�ò�}a��S�uX>[x_E#�deV���*���$�>X����kZ�P��膋~NG$�jsc}�rn��E=���m��<U�}��N��,�ܚ����"Ҏp��\�SOե�̗ߴ���h'\�[@MSޖ:1��������N$�.^� r�NԲ:+�	!.AA/�]2���[9Ң��CB�nj���u�t��̻�/B�%���/��sպt�;7�.�O���M�m���p��e��P���!�ڷ���h�_[ͥ7��`Cr�0��ѥ�+a<mN�O��,���D���A�E*�v;��lU��o�wȲr�u�����ص��j5Z i11�����a��^�2�	w���e+I�?����g2QSe�r�	�=N� �S���TK���5�ܡ��u�,�"��`�ϕ$/��C�e��"ۈ���u��m	���$�D-W�rN�8C�_�0�J"��?̴p'U %���p���S�B��uy�� �%�
�[,�o{J�ǩ��aAy��~��9��Ɋ��̗>�zT�>z�?�L��Zڒqg����S��I`f.$���4�
�j�2���D�	�l��'!�9��>8`�db��/���n����M�c0n�4׃Tp���Kvӣ×�"F�ddm���n�-t�0V�/6���t�C�� C��#
����6� "��+�5I�ɟ(�{��*+��G�m��f�m)��M��
���d�����+Y�n��-�2ϒ�V2��`Q�h[�ɣ\z�P�V�B;xW�厇2��:��µōA6��x�\�P~'��3�ȧtb�T ��Hb��}s!8w$����r�_�l|��y��'�-XU�!���<�����%'�����$x;����ɤg��n�G�J��Z�ZX��ޥ�q�֋]C����*֯�AI����L횔|��0zW���A�#*�1��%���&#��T{B��m�CI��K��#���~ې��{.���Y�ټ�ߨk��ǟ�x��U>��϶���5 �Q��	�ڬ�v!\��O�ލ���^*M���^��i�$��!�(�?Y���d��@1-�$�x]|�s���<\ѾA��!��Y֧�5#� 6��D%2C�b�Yp�T~�9<;��@�i���*��������=�0?T3�r�b/n}2�m��K����,\b���j>U<�&�7�T 0X�D��7D�9T��g0<|�/S"�6���pIu��en᮶TW�-}pv�Bl4p�����sP��@c�*��i�K�8�C�絼O���]��隋����#�Ve:Si,��6��%�����+G����l[�V�Ĥρ���S,�H�F��<��@���?�^ŕ�K������̈����V�e��9��v���g�js�߼r�o�z�³2Wq�����
�8%�D�F*�ĵyjm���:H�q�
�P��%P�@�w�B#]�04�Se�����Sh�"��s���#@�O��|��Q�g�ĕ�(��i�bp��{� VϞ����M�d��IXw��m�u�а�^r������y�	 ,��/���W}��%��$U;��T�y9Ym�<k-B������w�.,Z�KP��y�RZh�b�&�%�]�Դ7=׃�6��_"����=*p[��(�I�Ed.b��)$P�3� �3�e툫rݧ��&��qi��悂l̷�}u��z�CP��0��/D�1zQ�����u�~��s���7q��-B�ߓ��� p���f�HN�پЅ�:0RJK=�����!�K�/���{�:�
i�X�.��uu�7m,�3q｢�d~5�䩔9y"��+,ڒ+�rݓ�����>�S����%/���6Я8��LQȅ��;�98�p�VO*���`j�V-�G÷��:4��R
��(�a�>A����g%Et�_#݆	~%jeڲ��u�~i���
t�7�C��M �2�)O������9��W�������BN���"�5��o2S6n,�ZV/�����[�)R瀣�]���i ���5�
J��
���O��Z���4��_����ע�[:'.�Ҹ �*���d����3��k�nM+��� �Ov�Ϋ���Ii(�S�RE�2�F�iO�	���㰓.*2���-�����y�N�ic�l����!ox ���U�ȴ�f�����4��.Z�6F�yֻ���1��zDgB����ok�5%Xo��4��etՑ�L�\��?=����F���v��Y=�Y�A��)�]o��̣	��W�i��E��z}�в�>�һ�kό11x!E�	B0����i�,P�����|�nrۃ�&��Q�^�pX�e�[�g���G�Ls�h,d݆q�F��%g�7�^`W� %�,z⡥Ly���wߏ�����?w�rIs��tPa9��
ܳ�-�S�~z*�����G.}�ߠ���>����8����P�hsa�k,��Ԍ�x˺��9�6��,�X/r���Kk'��Rx�UN��7�{W�?J�,�O���<��� M��ms𹞢D�
�A��'�rT8����i�+$��h@���{�b������e�
9��IQu�� �d����Mag��BL} k7Ε���I+l}�|�s��U��õ�j�z5wi]u����?ٲ�3���E���_a�V�S�����l�*7�����F�}M�Y���G=���{Q�=���6_����9�3K�K�.��(�|N���1�?Ag٣���|��S^F5Q��"?�Q�~X�׷{(R!��xJm�N~���̗v"ם���P���(=e�R��P���Bo�v�(܆:��d�_�*��ߗ`>EG-ȫ5�}�]q��y{%�PJ��|��s�FƲ1|��n�,Pq��Cx{��,����_H��|P;��+�JX�x�pl�Wpbm�A�I�koN�O�5�w�FE�8�#|\	#�_��Pőx��
by1����#�>89X+kUr�\����(i�S����/6���KqR$�c�l�~:�z$S�\�R�/皈X��dy}0�l�{�Ѕ%�?s;��"���p��������dI���;��
$�WD8�;�5|rw�W91�
(�$۟�ǖ�O�5�*����g�6��>O{�ӈ|Rp�n��\�͹�>Y����W�]_ܘ81��񌩺�u�j���ԫZ����L�mN���-A����#�t���,���-?�GL�*O&W�{]Xӯy��&M9G���_Z
��<��m�<xF���=�e��R��������څX�^����B�ȭ�ɗ�MY8:�4l�i,S�0[�?��֛�ex��Ӏ�F��N-�5|1?��W�Ȃ�����\J$G$i-^8E]�P�p���.�E��.����Ia���yo�+�-HW9�k�-�(y����!ž>J_��O���JShu��P����	���ؕm��}�5�\(4��εw9щ����~��Ů]��2�7Ubv�S+4>�!桀[���_�E�c����i��ie��Qb	��q�ˏ����ز�a-x�+7ߍX}���X�#$?(�@1��o:�b�Ǎə˜j���^�y��D�q�׎�"�Ii�exPӨ��0+�h�!�2)�6���� ��h���)<��������%�N����;�hO875�����[	2�l�ׄ{�M��q�)�}3]�ƛ�"�U��a�S�ٰg���*ө��K�w|�Wc>%�|"�@�p��\������1���i�4��r�tt�z�A���2c�^���a��^:���>F�"�;�;:��&�����x��1m'�b���!':0[.�����g}�h�_ɕ!���5�Ŝ!���	�^"�)<�L}����DLk1a��^r�I͋�T��Ń���c����nw����:�!g&U���Ҝ�6+��L�e��9
�����v��M1]	j,._>4�]t���2(6�$�h����Z�@��	=��೽��N��b�s�ޠ����Y���
��g�s��Y�1�>o�g��7E}I����|� (pR��I�/-Jtr��FU��eQ���'l���U��@��v���,���pܩ���iQIܦ2K��Np'Jv�8�Kp���"��N�^;^|���s#�{��=�̘���١k��d�tR���p�z�뇘R��o�-�ώ�7>J^���9���	�8�P�ã�ԙ���z-m3���qX�#t�xF:�{v�3"��۹��)gntm+������L��*��ҲG'.�g	���/8�'�7���s�7�,s(eʝZ\���_[�`%�G�}e����#Tf��c��z���ޱ�����tR��p��`u�*0�	�PC���*vx`�_��V��I�6XU���#�y�镹�&����ۚ���Y^I�<�im�E�:�\��Y�q �rP\[D\)��͔��(ї,��4R2��c�g���glJ��i�#�
�r�*1�Vd��Q�ěݶ�'����'{�"�j��/�_ޘ����k��H�[T�**��~�oi#�����j�b0����W��{e��i�����G@'��]}���m�Ύ⣂������w �� 悧�������H��)����t�e�	*z�.�2.u��#!�6*O��V<���38=d���4�(�-�30E}��k�_!��+��|�N�SAC�������d�\eutJ�p��4�l��v(X�ô�o�쉡j�E��K�� G7����4��r6��k���'��#@��̸��3��CO���ܝ�a*3�}eq>�c�-a`a�H˼Zm@�}a��R-�L�r�>�q��B���=�6g��-퐷(H$�����Wz����6D��-�b��&U�Y`�$]��7@-�'�1��v{������r��?O2Ļe��t��?�Ǧ����e����~bS�x�
*4Eq���ѻsL�@�я�!��/DX�x�B1��ʥ�q��nA/�k��t���v�7�Zc�L��Pxb&�R)�Y=I)(~��q��;;�9�^a����E�P&��j!'&���U+]Vz�>K�(%'�c�d�Ks��!�C�иN��~MI��k�z�sLݜi�&�w5�Ԝ�����v���]��_;i*�1��c��Ѳ�9���h�f��|�P�W�s�7m}�!��uG`M��l�kǰ<��K3��z����g���qaZ�O��~'J5��r����x�t�0C������q�켭ߚ�'Tv��ڻO�|�9V˖kŴ�)�1+�-
W�����ܗ.y�i�Ѷ3]��
�ҧ����_տ7��ȿR��^>V���!��r�aU�GU�&[�k��[േhP;[M�<&w�ݶ^p;
���O ��q\$�>צZ�F��R��Q��-%�N���[�3!,D������N�(U�Ӝ�SEg�'��L�a4�����|1�!�:�D�?�=�M��3"~=�ɮA]SXlz��^�4�Jc[�%�� ��yXΐ|�%h�>uE��v�R��*���u#��%�H�OF��)=C(�K"r�l 9�KAɴK&Wt�sm)�� �����#��'S3�p�+�#���V��/$�W7��`: B�n�G�g����s ���xrqb�z�1����m�(sg�ós@J�3�4]	�6ZR�T�3&�K�(W%���k�=1·eX.�#�%��Z�Հ��\��d�h{���t�-U3�?�l1aj��nZ���RX���ht�'0<3�%�><��\���r����K��UpZ�@ks,Z,�}`�N�{����m�
�5燱�3������(n^H��6rT�/8���)Lд�e�����
������ %�l��!X��W1�3�ǋ�����-�&�p�Y�=�0 ��|Ne�fc[�_�7��R�~؝�E���d٠�����!�`�}���Y�����N�|w�ϴe�>��y��!�r�H��{i.
L���I����E6�ʟ�����>����![�Y*̙>jMw���q����[�G���5\-y���Ap&ttxt�ha�b�@r��#�n-P�U�����ە�Ҥ�xS��S֓�g�ޛ��}�=�ܯ@��ƃZM�H>�\{��S�ѯ
_�kY��Io�X���{7�'��{��ַ�?E}�D�hJ*-�y`A]�卤��b�Y����c@mX�0�ҡF��;��n��H�Gu}�@|y$�S�VI࣍X"H��x��q%���X�=맅���>B'��8Ҡ�<E�c4~�D��*x���ؐ�n���l�Ͽ�/��>��������|�R�?J��F
u2� �T��0eY�d�R*��Q�KB�Q�=�Oj��YlG�d��
tv�8�QkDO��w��Mm�Op�j~����@�����ǳ�U3��	U�o����G^�C��x�m��S����>*������o�7��w/Q�Du�������m|��/�B�|�o����f�[����D�a]��y�K��O>-M$8ܽ��~l���6�$-�ж�ȁ>�^n��M�[	��>{N˓''��}��5K4}[�^ JFLR�����2n�;�k�ܔ��>�����Y�/�g�3q�OA\��a�|:�Jd�u�Z��
s%K2T����MjqC�S������<:7igk�r���j#��a�Yд��?���x�x�_u{`#���W�ޙ ������R,��� ��y���2/p�p�tw+[����e �T� w@{Ko���-w^9u���~9ȫ���ٰ+�$��)VJs|�ڌ<�?htŪ#<~)&��:�t�by�^� ��FE�2�,���he�l�J�EC�u�Qn��� ﻽� #�x�k�O��ۜ���h�âa�u�"�;�]7��iuJ�=��ώ�/�Vk�9b�Lu�1l��7O��^�̘*N��Ϙ��*��y=��a�=��&N���7�mJT���q���~������K�x_y�~�pH���v]��\�]��-�v����)J�K.�w?o]���ç3�W`�xTLAs}]g hW�)Y����E]|4�=�llk�p��eV�߄�)��߃��^�/lOLU��ֵ�d���x��b�p��<��p}��P�O��o��~�S�4�!k�ye�%F��<����p�t�#���s��b,���q_�f+�=�iBO�ԛ��q����Rz��O2��|��/�N�6-�~�p;z��V��5۰�4�v|~9�g͓���fS�E��0+��3&��@#�Ġ�q�HW��$�����덹�:�]�S|��ul�ѓ�\�W6-�F)��,��G&���T��1���2�����)��z�)��Z����n�/��1#ͧ��u�}�1t�5���U���JbϒW;�Fzϱ#���?ͧh�&�9 u�t2�D���*B�[h�K�`.̪Vg9a׾�Y���x�hr[�
Ӽ3�_��=�2��.7��V	��P�ԛ���>������RP�V��&����.�1��Z�����h���!v`������q��n�0N�;��q����� 	v6ͨ��Q�vq;P�ww��b���L�$�'��'H�l���{_7r�@/Y��F��p���;F5��tIA�.�����_�t�N�|X6�R1��؄���V&�E���}m��o6�|7�a�	%5:�iw��X�([맺
�4�b��[�m�I�me����eٓi�8ހ��ƺm\P��ƄjY�|�1>vFJ�ϕU��@�z�x�|�%ѿ��G�ħ�_E���-��_^���ӓ,�-�̱�.N�W��x]���.�C^)�O�������!�a����LՊ��{�Ө�����-߳_����1��Ha"b�F����7�5x�t슿���*���80M�O1�Y9.P~ތ��U'��9�Ȥ�*����2��e�PZ�1�m�j�}&.�bO������_�J�*�������SR<���B�S@�c�B������2`�﨧�[����X!(�ΟU��WnO�	����m������s����Ͼ��xiw��!�m;d_��s_�ō�����G[�w࿢�9�����{���p�v�p`�Y:���B���;�x'2-a"7��:��Fp��d�f�R'- p�!�cY�c��0�
���B,yC�sK굄�����y7��h|Q�2�������/<���9o��s��ю�xV�7��V��ʸ5��~:	�ͽ�H�ǝ�O�H�M�]-S[����Wj#R�
w�������+�8��V�6��6ѕ�w��oM�m�m3�� Z��?�z�[=6�Df�H�����P>VeT�ef�P[E�!Wy>�i�ɃN�e��75��K����ϖ���w�8����ڱÓeV�����0	�7.4`��W�1Y�C��,���	���&Z?!�{v�����`0�/�zq� �5�Vf'���ֈ��kԺ#�Ӓ؋��9� �s ���Ċ_ø)�^�`�Q1r68��Z&a�}Xŋ'ή�p���/�U=�k�W��8�uٴ�!�J��A^��̳η��]�䢬W!�s�fFc�7����}���I�ǳ��~�Y��J�X�QJ�+��z��� +r؁�&I���S,��;z9EF�a\��m�{�N}��ҟ	g��;�nO���ur����U��vd���	�aó�Y���q�gH��٥���9�#�-ֵ?��_��7��;S��]���,�eQ�[����^~y���O��B�l�ęl�	���J%�rs� [�;ޔ��F͂�4yHr��m95�n���p!X��,4[;H��_vqݟ ��������5@n7\�7�f���ޗ-x5�ҕ#�]���n��T`�sL�WDKҏ�;�i��q&VS\N�NT�~BdKn��>q��ЖYT��]� (�j�x��0Vb�n!��x��N��7n��<��Um4���dOo[�᫤,��!���S���mz2�\C�؛���T�1_4��	J�?�Kbp>��4��`��w�9���z����bJ�uy-��\M�)�@�K��'�v�u���-���<ĨF�*�q;G�y�7�`b�z�}�uTiJm�|*�VY��PMQ����{I����[��s��j�ם���mca�-Mrώ�MD4̹����^y�1=8�O$���[�H��L�#B|S���%�XU�d��Y[��Z�����R����8WUqcЧ*��.��C�5?�N�/q ~Q� E�`ի{S����9`���ܐ/�c�r��}��,�i��8��dLI�ݪ"J�]��f�(�����0�N�0��Τ6�$aa�>��)h�����/HcN&���Z��ҡ0�H1�o����|E�L�Wbۿ� �"s܇
�
@TsU3$nۮd"8��C �I[P���mxG���-x���h�>�e/��q�mEW)����qފC�V�>���qi���}�Ko����o�R����i�KX�=f�Z�����>:F�a�v_���ecD���	�� ��3(+2���o��	��H�c��sa�>�V�j�ϩ�;)�m� ѕ;]7�K)�����tg�r���?���
5#���≸�Ǚp�h$�ր���˄M�h�?u�{�#������ĵ��$m�|]���o+.
V��#���J�}<�,ʕ��m.W ���$%�1�}���m��Wz������WO_�<��N	��2"\� ���ܨ��b�a:�?�|'�=�W��	�N,3�����>��J��i�gdȇ��э�iq��1�
Z�kVU��Ry3��m��`���M鸲� 	�(/��c�yϾv���y�SS��z��<M"���{٥�Q�=>�U�.h�����ت�{��A<�2M���<[ԮW8����׉^���b{E��e�9�T�Ts��+��!�����ٔ���\x@�ܛ�ظl3���2���{���=<o�>A���[�;��9z�f��y��v#g����?b�b�gYvBi���7H-t=3A{J�W�ʼ����3@�'�O���%\^��ȍ���ԛZ�_�<f��W9:GBQ3����*?�$5#�9�[T�>�I�n+���ܛF��q�+��jJ��,0
W�i��~��vi�s��R3-��S�g��6�}�������|޺�W.�6,�{�Q��i�?1Xk�L�}G�������}�\����l'F�n�Dk�{VNa���v��n�\�"��>�ٳl%r'j�JD��u�XLU���������r?�E��,�<I1�a�3���o���K�\�?��!����ff��ʢ�|<�>w}�)��ƴ�,�-s�<[���c��ܫ���Z(3l�ȝ����3�[�ґI��k��������-�b5,2�[����;���I��-��[lb��o��(.+_Jn����v�U����X��Ǵ�Kwb������[���� �д[�m�=��˃��S�UR���dK�RI�$P!�΢݃��H:�uo�oYĲ~	5�j�0�/�'h�b�����ũr�����NuŷC���Kl��y���?�>�s��J�`!�������d6v��
6����$%<?J$����Q�t�Q���Oovi5o�;ia~Ug7����P=���WP��q�~���%;KOU�_���5�&Ef��)m�-f�s�����-}���?�U(���Ju��vF㟙���_��_Q��!��X�/1*F��B,��+&�l��A�F�i+`0ĺ0�U���~��70L6�z�q�QD������$D���gX���<�Q楋c5���;��.��EsP�n?~���Ws�Ũx ���}�f�l�ɘe�_�s����NY�6��JD(�<�ք�y܎S�7��c2k�i�h�6��0(�nǕ��G	7��0��a`nL�ghwk2��sT���+�EI7�#$�{)�"ZP@�<"�j5Sqy.v��^�N�%�A�����&jgi�^SL��@e%���d�b���_��?t����s�RL<5V�C�7�(�����[�hI�m}���龟$�t��B1us޵��05����Lq>�����òFv��TDJ+�+�h��9�>'~1ZF�K{m�R��Z6Zl3�v$���C	̛�a^S�	
e��S���b����À�}5�!}��J<ԙ�|²�!�����n�t_[�|!Ӝ��c(���ږ|K��Ã�d����
��ڰe���Xq����(mE��\{iՅ���X�|~�w�2n��� �>� ���^Ԩ�Ǵ/�:�����1��l��"�ζnd, ���t����?�sD����fi��&�kT��cRߟ"��j��S��ȫ�)z����m�L�IB�xŴo���|�C�W�7���F�kK��l�1�Qb�L��79�L��H�dM[`�'� "f��	jԲ����<&dYT2��Y8.��<��>U`p���u�<�]�a�-r�Q��s���8JԹHnU�˯��nLF�����'��H[x'��Hl"���Y��s[�3e��[ױn���V�M�갢V�DK�w�ɖI���X�IH�I^�"�{@��#3�4�_{
��݄���W3���5/�d\:��M0�q��ĥ����G��X�f�T6��]�:�o���*� o��w�܈�u�f	�q&"9o�s�� m��\��C&��4ʿ�q������#ޗ�+FA�;��hДM��{����)
*`�c#�i��0�F�bX��`v�kC�S�ɰ���P�d���:�r|VԗU�׶�PB�S�N��ɏ���K���Ǵ�*�S׊n���@*�v�n����1ZXZ����'2�3W� ���Lz�|6�{�u��'��������vI�m��E�T=ۄ� !0\q���k�m�oEj����O���_�4m�9[�9G<�~��\GB���n� k���i��Ps��4Uxnt:��L�>ֹ(�պ�����r���q�8�z���<�O�H�a���l9
�?��X�3r:W����0�����7���+��}��Zj_�L���m�dCe�EO�uN6?	�m?����͢\^�
I���_�(AHm���ԗ��
�7�N���%[��>w+E(���g��t�#Ϻ�5ːY�WV�|�ݎu�^6��|X�&=Z0��FN��/?PuHbhJy���4�z�ฆQPLP�h��<�֙$�P���;����OO�\^8�2qf�X�S����»suCDÓ�\=�_@����"���}�L�݇�ȓ��/V�=�I�m���d�8#�VK�ȼXa�Bo�́�^�6A
}q"�Ŝ&��9��VRߪ8�ś��>]y'+�t���&�(�E�$���I/�h�~p`r�3d#���+�K��%l�������s�(��ڜE�1N����ܥ���ˮ,?�G�_U3ܧ�}�'
]��W�*�H��ў:�ԏxMU��uۋ#���4n�[~�Hf��(?y7�y?�Aք���%�{>�.ȗX}by�s
�7W��eA`�G�$x�2_81%�U�-��7������['
,���^Ē� <�{m�נ�=����3���04���$�ջ�<>[ԋ�f���W�Zh����)�̒�B��\A�'e����,)�'��j��
�[�ߪ� YC�p���9H��H���E)��`3����9�?e��m����b$q�0�����s���xg�����|�pl��T����E��Z�s���q_]n�p��£Dxm�k��z�:*��\��i������?�h�/��0��q�h��Մc}�s�j%	36�P���������D��݈��hj��l���a�W��|On�U��,3���,��-+3%��k�>ʦ{�^�9 ����֌*K�6�
L���a-!� ��(�9�l�1}�&n��m��HF^�{�oᰅM��x���YhM�[�(���&ke��X�>oR,]�d�Y�Z�W�#��7$�m��m�������,<�����,yS�Jk��	I�g�->Ͼ�3<���V|�K�'E!�YS3��y�h��5g�
���*��ƍ�j}g�<�8FZ\Q��?p�0�`{�,��_R�~���ۂ�����epi?�����+�Lx���uh?'sL ؎v�q�h�=��A�|���V��\]��W9�ӳ�w{�=��;�
�ɠ[�}���n֜��"Y����t WpUs��1;I;��s���G��ǗZޝV?��ej��b5qKu�r����?��p����nF��Y���H���CCU���9wd�"n�i�E�ql��=�߾XP��zb��>9�	�a� hq���u@�Us/�&��SC�S�f'�
��NM�O��YU/�O/f���GZ���n���p�x9�-B�W��X�EL-����^����Q�� (�4�a9�v�l��?���R��e|����	��i�c���&Q�9��<Ԕi�J���m���븬�5�� >l�ٻM�~BQ�ĦU�J�=���+ <'!�{>��^���*���^QG���G��7ߺ(��%u����8$��\��s���Z�=���(J�OY��T���J��l$J��h�Xf6�Z������~�W: ��'f�i�~%���]o�i�5v"q�e���J5��IwwM8��ؐ�����'�<����u��|ΐ�=qd��.$1�z�gY
P#P���tr���[	M�w"�޼"C�>�����y�cǭ,ҟ�f�*�_ӟ�����#�ᬟ󭨁S�k�Nּ���Xg�-�+,�^wF%���2F��_�	�˘�p��3��>rR�5�.��Z�^���Yg��� �*����4&X��jd��/s�َ���I�G��U�I$�\�BT� �!�cn��+�����G��x�3:U�yy��%f8`���F�H��"5�Fm��p�~
��cdX���x��~H���$�s�Ȍ����-N���r
��#A�D9�9	���X�O���Ȼ 4��d57]i�=p��l%�D'V���2��H��$���䪴͘��8O{�|Sۍ>��o���q9Qg��i�z�Rr��W��N30�(;��z��#ԭ��g���V=�iB8�:|���w�!վ<�6���։8c�s����;APB���=�fQuKn���T��=�Om���E%?��$�K����2�mi�5�+�|
+hc�T��w���h����#&�*�c:�#��e�i���� ʆ��-D���:�N)e�ͻe�(-�9%����<�*\ ּm?�7wCZ�wG�ٯ֐�o�B<.Y-�kݓ���b
��겏iw7�XSlD�o���"�g�+��&o�T^��V~oğ�z`�s��NUi9��10���g`i�`~�Q�/�������W����y��;S�y��!"9�e$A�U�ʒ�&��wɡ��"`�!��Z-�E�︸> ��[N�}�0�dl���8����M�i3<�`���v��=�"�KW�n]�paU�=NE��ޗ�����`��o�-Ë	��@� ��m׉�w~������g�=0�\O	�+��:�K��yTZ�mSk��tB]���}�y�2PO�-=UG��[�`���1��c�����ŦkL��yq��j�����:6�h/�P�'sY[T��?t�������Ü|j{U��她K��Z�J��٩����>�Z�t�*��M�N����{������;�AD:(��B@�*�Ez�݀����� 6PB�ޤwDJB	Ez��"��Bپ��p�=��={�Ͼ�{�;Yk̵֜����5�5%�?Lm�]��+�'�����.�0�R7�9M���w�9*OE�����=�Rʇ���\Y��Ƹ�RS�}�G}<��F:9�߉�����'R�Ϝ�.Z�V����{���a�f�߸�lb9���F�GJ�@\�#.���+U�q?V���i� n�G���[���h��`�u,�њj������3�c�'	7�wʮM�W@�o�Xz�,n����V8/*�"��[���y;��Q���
��^��J�T?Z�<RW5��TR���3&ezʿ?7��2�7k%N-�a��ɜ��fs�H�_���1�
z4�{����b��5���{$kbb4ɒX�� �ERi!G��4�qB��|��42	풎g��$go�U��KKA�T�!GjF�?�d�-kc�Q�m�L��RkAZ��8W*��JkC����g�.�&#���_���Xm�_YG2����,N�����e&���b�`�K���"�履:D���`m�U8�[�	�)w�l�����4
UR���x�iT>T_T���x0tAk!�f�����~�X�$׭��2$b����/ɴYi��'^�)[l�^�{�(��9s�%@k�n��������z̉o�o��ڱ&&�4mx�������x�H�9�{@Ħ��û*qI��fa�������P�(����:�9e�Œ���$�;���6�%���r̫`�N�-!8xf갆������v��G_�âW^;�i�c�>�_�u��IS��^����
{��W�U�iG�L����«;p)��!8t��Cq��3�����,����ac
��'����E�E��jV��c�wg���z����k]��N��#�7��i�� �S|���)d�q2������U�)x	`�x6�0S�ZjS`�]�"�)�m7�~�������-
Z����\!��q�SX��T���E�_6U�7����k+�2�E�rlM���m���b�����!*S�)N!��� ��8{��z��4{A_ �Y6���th,S�>E���<y���Wh�S.uې�WZd���q{g��>(��;U�U���7x�¼j����θ��R�nj��s���i�+u�¯�󥇜����El����v+
�~��`��uWwb�*����p����bN3�t��&'���%�21�&�Œ���H��e��]����6��?��Z����f�[��VӶQ��m�gt��G���
���)5��bbMu�Ye����6sr�����B���.�� d��+ۛ�?f3���SԵ��x9X����W��+  ӳX5��aul.辿�X�;od|��C�.��F��.�/�ݸ���g�����C�RO����ںe�����m����B�,ۧ�}'�(}�8'�N��)�)g��^��m�2�d���뻚7�r	��l�N��R/H��}��<��������� �ܟ�䌡k�q�B�$Jt��g�)y�^�Ck��_�e3�ﱮ��Jة��m�tP��8͈޴?^���K�s"��E�`�O\|��.�ĕS��TH���Ό-A���U��:vJ�����+��-���,'t��*@MV�`GE��b�E�@"P		�C�*H�k�Œ���\�K�W�xd�p���7oH8��$oZY���">��63����"|nF~��X�x�ф��y���¶�m���!��T�`e��U'<�A�jɮx�o~���t�w�����n!�����Vc�^�y`�5zL��-6��J�����#��E4�j�G>�[��ZW�)�A$��mq�dI_���#���T�
��� ����q���(��*cN5�|�;�^��EM�$1���AT|>|ho�̄ﶒ�f2_�J���3W�O�:��BC���f��A8ؓ�J*8D���&���M�1��^<�q9�Ib6�PpfDK�L�G5�5��L�U��ѯ������=���R��EBi'5p5�	Z�w� �H�4���IZ�R�T��af����sk����ğ���
�%��=l�`��Z=m<��s���]�o�0v�����ZCW��p�m�f��I����g����e�?#`�p���~&:�T���h�)�~��_� [��RqZ���a��^�=���|�*t�/=�\ֺGڪ�r�܂M�&�` 2�#g�ʮ����ʶEe�X�3����~��JR��Fj��	q�$o0b�{R��;�r�X@kz��k~C1dZEcĝȷFP�/� �ؤ����K85���Z��!�� �&����y�3��C}Ӽ�{5dtP�Ga?@�)[��3���D����=��=�b�IL.}���*��cԋ�uE��|���x���VqZj�>o����F����ˣ^uaȶ-�j�"�K�"��֝��E�=��<�N31%�d[�9������Y��Ao���.�r]Bn��ůM���J�;�ao��ax�z�^�Ś�CP�[�W�\��uȎc�����!C��R�S/����[�6�����GĤz8]�|�l6KY�|	 �zv�E�qg�`���ľ J�Z��DK���qt�q�� (�����ԍ�'���i�z��/��\��d�����M`z�}ش���f|_uj/���{�֐z�$*�n��|�ݺ�4�6r�%�<Z��w����}-z��#)�߳�;��)�M`F:���I_�N�Sx�g֎o4"*J�?zF��we���5F��_��N�^�Gg�~��Љ-���e�y��q�-#�Y	O�cs�tI��]�B��
���?(N�˂�4.�_�Y�M|آ��c�ȧؤ�t3�rIl	�	��oa}���@���$*���;ܩ-S�!~.=�.�̹��W�����-���R�FK
���\��i�!���{�[��3���%DJ~�ݞ��S}RW���]�B���[�u��R��pl�uqXt�S� �����1~1"�p��-�Ξ �1j���*E���;�]5����=�5����U-��'�MR�������!mF�wY������Q(횤e)��;ۉO��D��c�0}��,ZiA<�@v�ku������v;�M������5�B����D�qv���1$᩿�6|���x�����������iq ^¨�T?��$�[�Xjefk�����.)��P�2QE�^�^Z��6�qJ�H�N;��ƅ9��~��j{��Ě>
fwb��z<�fy���G!ܗz@�>Z�5���ӝ-����iV	�#x2��>M�p9������#���j�=��(���w8Zy���ķ�2�ǧ}�t�|�&����[��a*Ռo>���w�kM�-�U,ד�3�7�XՕ�E;����t8���p����c�����x��SK�`V������2�)P!�Y�щ��aK6Ҥ�B�|K�9Z�*�[�5+�B�H2��o[�a��ve8�ڈ
ҾgQ���zD-�? g�L^˫���y�j�y�r{�z�2�>iɻK�+S�/o0W^����]6�PU�� V��y�HGؔ�v)���s`���2�z�*�� JtB�����IE��G�҇ox0F���u�W���z���*U�銤.R��������<��O{���PU2�t�WW>��3���r��6z&�_��n��$�n*l�RO���/����8���?�:�V`�R?��J��О���G3�����r'�`���Lmb|�ц;EY������d��C6�(L���/�5�{Ql�mJ+0Lŏk/��6�����D����=2��%�-rU��;L�][�G� ���Q/�!�c��L��JKc�T���R��!g�<��E!\��pP�ΚPGc���w�$�Z���d����~��-����w�P�9�S���P�E ����?4q��ݐH�����q����m��pN�o�`	��hŁ��Ʃ�^���\d��|�|�h�>����p�c>������܎�ټ� ��Avޔt!kk?�W�T��u$�=����5���.E|bʭkQc	��M���E��5���a�I�i�S2�Ƿ��
C�6%�ta��� qӂ)�7ΐ���q����mʼ����������Ǐ��rgb�s���Y����#�Ä�p���۩bI�<�]��U,��h����<���ҝ
�h�/�>".�[*��	�g�j�ģ���q�j�{�1��7zj�NK�px��N��fDެ7���5����*w�4I���v�ŁN���������w��?6RTZ)*��T�^��r�6�l�\��+m}�oж�+i�N�\b������}������F�ӪY}����r��������%F������C�e�c�*R�������C )I�U����&�֚���W@^5����+��m�>�&kk�$pk8[���n��!*q4�F9�Q�ޠ�2g[h'L�}��C��J�_(O4��X�$jO����~����	T�{J�-
 �ނ�F�S,}�ׂF��v��/~�X��q}lgɒ��`E!�EJ��D��,/v�Í]嗀��׏f�6yJRkd���,��Ү�r��	���ܽ��Ţ�����Rc?p�K/
.�{k�����V[����`���Lӳ��w3%�m�����3fx:|ṻ�/��9M��O�K��v��U��X����Ae���y} Xeo:ڤ�g��='�Bʽ:�*��y��pQ,�|n��&[Ł���(���% ���ĢX�¼�����%�ll�4� WB�`H^ �B���]����}�.e/�N�5�O�:��
qyF���4�q�K���vɗ���:���LY��|��٧��Λ�����嘢e�z���kDj�>�h>+����ŲH? ڲ��ru�;p��,'��i���i�j⿋�I��<�����ߎ�����-U(�$4��'^��=�9i1j8�aYe?����gP�)�0.m�v�P�]�����<�E`-�lɩ
��=�!��+B"~GK�qc��W�Y3C�r�R��)H5���z	
X~�s���7�o/Q����A��oA/��r��������N�g�!vܿ�^����w�fe��%�������w6�����w	�U�� ��5]��Tkwκ�!&V	��1���Y1�s��n+5Q���j�lBA_N���>�ݷ6+2�5~{��C �9^G0I=9��S�\* �J��؀��/���|� �`�hA}�u��C;�Z�����6o�2�[n@�rs�:�ȣ_̌W𣏵� C���6�/��1�`���5�/N��?���S��>���	�n.~2~P��p�G��ҧD3�tEE9�%CN��5�����j쮀e���^7䩧�ʒR�q�3vUIxg�j�0�~�٩P��C�4(��4{L�WlkZ|X�Y/�y���s�Wz�K���.7d�4R����ϗ��O,Q�:[��u�M	��k$��Nn���Dv,�ʪ���?�m��>�(��2�e�z�C��[�{f�S�)���V����Y�x7S���:���:ÌP�V=RF���oË�?����5Y�&��R�u�
b:�;E�����5L�M��޵?Q,� Xx�^���v�8���\Vyl����������pa��g��B�DX����G�{q�#�W������"q��) T���^�w������n#��?�Uu�	z�b��k����~Z�ͦ1L3-|QlQ0�~,��z�ϰ"��(bMmӛW^��&�
�mQRq�u0j����^����<�g��>��h�u!F��E��}����էf�����BE�.�#��#��3ɴ�H(�,ة�f�9�Cv��}Z�o���7S��4u\���"z�[��-ٹ7�`B	�贽db�j�(q~�x�)k�u����Q�q9.[�>�^�4f�c��u}_��1)�G/xnyf��%p�O��(9��l:�~?,.k��2$n���\�뛏Φ~����`·�OW�E�;O�z�ˑ[x�|�suR!G��b��ā5�;>6��H+�S�98<�*��݂�=����0�jC ��������6	��C��P�$��rp@�S���e�k�������@ �b�C���3�P�S������Ⱉ��`ӎ,se/�L�ps�<�Dl|�Q�{Q���ɘ?��ߝ�N�^B�Fp������e��vJ09����|pQ�.�:%s���۪����Yy�[)�W�M���[=<�K�����Y����N)�.~܉�v�z�U�I�q�a�z�˙Uґ��^�Yһ�aIiqz�V��N��/<*�*RN���U����%�=����TΞ`M^�{R����v4��
-���Nĩ�a�`�F�I��(�(�g�9�b����zK3��.T֗����ֹ�[0�OźYM�`|.,,|>�	,n�� ����l�8�/��
��Q����qQ��������C���
||�e"�^��ho�n�I8��ñ~�8�x�F�������2Wq�Y~{D������:�#��^��w�b��|�5��=R�	�0�� ��F�
,�~�b�d�ň�����3h������F�O�/�8�8�y6���ԓx���3�K�ݬ@Qw[�*{6��AbbSV���d�/�Pg�ʐƵ��{�̨��C� ��b�Z��^�lyGEP��q�W4m
�T/.�%&C7�E��Q�\��ͧ)FF�mg|��8v��5��"��jy����TA� �݃��A�C�!)F���{*_F���)W��G	�v����AQ�/�PW`#��I��	x�]��e�Kjsg��̾���0r��`�t�>�ҤW �&�[:w̠�Z��aȚ���-�����͝��ǒx6T���/�A�fҤ� ,�-<�Y�j��2���
>��(��+�F�[��(cM;�Ȧ�BZ��%C��n_�w��A{�A�v��%GT�0q��e�*���*�m~t�|��n}S(����67�j�t	0!;T)�i5�ZС�2��P��|jZ瘟��l�<�cOlC�����#��]cG{�[������9I]��ܲ��@K!w���XP/n�e.UB��Zo�Z���Hh�j�3���6��JҞ�Z��4á���S&<����Oe=m"��k���R޵��+2�F����e�}g�#��[����O�c{�Jp������QB�׻��]p�\�v�����բ�{a)6��YO�>fm�����$lU�ltSddT��~4b|�+��x$�!��41O�Q�!!}��>�3ܒ���h�����2!�y�@�"b�?-ͨ��S,_�N�꒸|8�3aIc�ݧ�Cxg(�]OI8��c�C���E`\���K4T[u����h�&��������7i�B��Ѕ���Aʔ�V�m9W/X�zzc�~��qީp��T��a�w��R�]1���ڪVW���(Qtݞ*1;�;Nhū���%Qr�b�LJ�gi�V�L�z��)((�4�C׀\h.��,��Bȥ����$V(l19���@8�L���*l��_�����D�����ᓾ�1Az����1� ?S;��9%���8�k�x�&y��P�� 0��~yL��}���e�1~6���#�;U�F����ƛɞ����`�3��aC������Pݭ��j�f_�N�:�S�߻���avl`���'\;!Z������ב:\�ka��?��q"qHl
��#�m����CW]��O��)�НP��=+����wO}P��7����EA�:C�?�@��=>�@u�ivj�)�F͈��Yx�=�J�]f�{�D�I�j�M�]%��0_m �a�m��7�-ˬ���!0�a��j���G�1��)� �V��7i:c�wR���{���,�H�Ͱ������2?w�u����Yu1S�;:��}���R�;��K���/��]�n�3�����R�^/�!�����ط/����
N������QPg=�R���I�l@FX�h*_	+���߬r�ғ�I�N�",vz��x�#M��H'NE���Ъ�r����w�)Rո��JG�{����R�.S���3��dZ�RH'�E�cmk9uY�%��Ћ$;�.�1�Eb+kv뢠$����G��O��]"���{0��"�*�
��i�h�9Bf'���hw�%u}q�D��p�׫|z4��:� �\����is�Q���� �V��0�pC�͉�I֐�6����;>L��q_�W]i�Ԭ�6H�2��E�2�͚t����%t�+�������R��LI�V�e��V��#�4 I^*b� Ѷ�`���w��c�'���'̦^����E���O��J\��9ڸ�fX:������<�q�O��1��3�?��X\����8ר.Vj�{aI"!�f��c���	���x.�&�ы8��;�� �d/*zJ{G�r�pl]:s�ˆl^�ӓ����Cb���;��~]�k��g,U8ߙ2���_�	�ɝ��I���V�nS��5�9�g!�^�0��wʷ�yc�T��xqB�]��J�'�1�9�]@�E��w&��C�9z[q$I�`������J�V�?E��^>�jK�AO�/��7+*'�l�
�Feua����0q�q;���=Pʍ�&Ka+�tu��+L���覟���z�@y��M%�� ���3.$������e����o�c$ʧ/�V�#V����}߬�{a �k�S|CϽ��?=���Xw�r���I�����������0�C~5���o����Εw*,��]���%Y�F�g͌J+��PL�KM�8G��C�	g|E����=���Xt��{��`��YF��3�$��F�C�򌃈�%u+���@��AW�����vb��V@�q��7k�qy�/H2vs�B��~�7V>%�(�fQ���1\ߘ��͂5uG� z�F�0� �1�q����f����v�U�X�\0>=��R�O=s������л�xp�SA��ј�Ui���h�����p��U�EK���������bUM�B���'y0�WR(��,B�<p�v��4gj{��Qgؘ]�LM\��MyЕɓ�����w�����8ϕ��km$cn��d���|�M�P*�h���%ln7G:hgZ�%�c���������������P��B�^���s�*un�%��6_s֌uy��0#j���L�����f�:�E�->�j���@���Loc<I�ީ-N�^�|6R")�f�TҎ~}O酞�@I����@w�?*\-���?�}�[��k�-8�b��9�ʱ:Hz��r�v�����č9��ز��7�����@8���oV�B�Ђv�.?�RkL�U�l`����K's<�\L��3[&�[+!�*�h97ů��5J��4��ۋ�_��y����87!�5�)���_Jd4"��J���^�KrU�������A`ۗ|�2�Υf����h��QڈI���G��w���h4�v������r
ة�?,������].�D��a�O��zJ��%�q�텄�֕����Z^P�g�\uA�.��Q�S���L�$�շX|�ΗN�E��S��UsT�
n�Mb�_�M�`�� [�k�Td�v�l&D�����@W�JfEA�|��GjwO��1�����?9eCr;� v�N�Sx��P�8oI�lq�&H0�h�m�s���F��>���8�Ǿ�k�w+���uFN�Բ�#�c�CG�!]����黼��$���;ޙ����/�{:��`S�EI�B�0������	�n��e〫�?t���Ŵ.N��9��v�/�R���a�+����['v���0=c�u28���ڵ>oc���]���_�I�9pU�.8�R|�8a�L�����B��t��Г-�K�6�C��ww�t�
��1Fx�]�E�X�J���	���/UH)꽭b��5����Z�T���^>�w��M������%�rX�Вh�c�z�� ��њ�����3t⮙��F���G���Im���޾����s�'������u��t$,H1����)G
�X'6���G1�|H�jT�mo�=#A�0�c�[�c�}�:��$��9�Yh	�Z�(�j��;N(לo#�d|g���5=\
�ykh&t���OC�'��R�E=ޜ��>(�+|������g�`�zR���Oje-h���tK4�������U�c����^�GpU7�?��4F̃��r��f�F���#ʦqOz6��$��]�8:q��E��w���AM�sU3��q�G����	�a���?A�|?n[ٜ�����8�

��իV����w�x�TЭ�ކ��?c��0�6wE���
�=\&�Jik���j�]�L��u�9ZgZ�x�h+�X>�̧��ϳù�X�S��~������߭���Y�_p�E�A|c�On��Ҋ:9o`�-�M��[�	�y�����|a5:P��� Wӷ�Wa���i�f�t���!'�Kw%9�������Z'p(��8q@ًВUr+_��د�#��%XAɽc���o{�ܰ��┆�!�*fHEyc��.7~��)�S�� ���S�Ƣu�Ś�>�}�hgjy��Ӟ�i��Ze�H�M�������	�5�2���Yk�Nw$Ae��G����b9�X�l`�yM��fa� a�=6x�k�zvW��i�	�)���gS���#���~�7��d���
�(�٬����`�o�0T�nK�����:u����a�m�oGc��DCq;�D�����&D�0���g�:��[���s�iS��#<�CMv�B�@�Ȁ�q�c;�=�:�V�nm,4��[�D^^]0��*N�s坽*���Ѳb��kg���1y8TXN��^t��司7�2��W�]>bQ�,P��=����Xl�\~O�~)l56�p�[���gt�
�U�]}�nޣ�}Цs�GP ����J�WcCח���W�,Z�nb�y�Y?�y8�OW���?e���Ve��Ϙ��iե�t������N%�߰	1��h�]���V���*����>����
�I�OUí�wC��,f��vC���D.Fs�̤_N�=�fbզ����"��.0ws�[��B��J0x:h�6� �d#��1[-�G$��b��7x���k?�)�=���Ag��A	.{��o�d�1��`��1f���k��Y���� x�v�n1k�ݎs3�'�&�d2x��a��,ԓ���6�TBEG��u"}���3�kV$_�����S��砪����B�ᷦV���D���a7W1���'���v������N�@�0eo?9���U;�F���U���M����������?�+�Չ��oh��#�GRb^��FJ���@�B�?X����vs�L�scP
2�usC�@��ۼ�p�n3_3�f��@%�=�%4����[n��ȵ"�
P�3p�,'�"�0� �)�:]��c�:&PQ�w���~���D�L{��a��C�X>���jk��#ⷖis�t��O;�g=剦�Q���l�*hKx\|V���bh�����,��R��ș`�z��D�9r~uX�(Y
�K�P�n*)�]�y�	:�?�V�9�D��'x�k���W�Z����1�#�V>��hh:I�,K���,���ufy�k�`#�̺y@D����QR�����6��/XU����B%�����ߒ���6�CC��d)�R.����1�Ps�Z;�2&w	�3#YX��V$��h�"�0s��Uq�l{���P�aX�}��a<e|a�q	�i��9�F�6rfc��Z�I�K��ʢH<��n�A�h�G�)��d���U, G4Ӫ�?�Ω=We�w��F�`��ܝ.���5�A�C�����e�յϵ�ҝ�R�u����ov槀��t�.�E�fύ��7�m'����q�ɪ����{�VO|XwN��LC�3��o������5c��P�tG�3p�@�ԁ��؏�[��z-�?�q��{�%������K��M��� �H�`^^��x��85e�8�v�g��w�U��8,��������q/p�;u�����~��D�ݬ�e��.7?��
;�AQ+]��$�����X�w��˔��)Fj�O�
u/�
�ʟ�_d�cx��i��do���7N'�����n�͎K�3���{&�1�3ۆm0X����-A���]<����:�s3�^��
�X�l.]H(��h�آ3��LC/�<)wco'����^�k&�����ZS�ep���7^VtR���i�*�ƾ
D��ɿ��[��k�Ij}O�;B������	?�7�Rʣ��>W���(ե��˸�RcU�'�ƫ�����P�vS|�aߪV��b���i@j��|�v�G�>c���W<?4
�
So�z��'��~D�g���\Z<�pћj���,f�e�]���5��~�V�P�B��E>�Z&��R6���/䴉���K��k�k7[^�=��k���'�)z�̓��e�&�F�\�,�^���5Q���̝!gh��a�
���O���`0��//';��o�c�Fy�R�B5I���Ww%�$��:��,��¸����ʝXڧلg5�I����G%�~P'!~�C�4��@B�P5�����SQU�Ɗ��TB�N�J���i�_�2}���a6�o`���5��U3!=E� �%����أfW��J<��X�T��Q^����u���*+�>y��>���ÕCy�z+@Ѣ �d���X?�Z�~�E�MC(�9���H��ѫ<���2.����R1�b�á���/pE���� �KWl&Obr8�؞�I����C[�\�v��ze��bڽZX��igƅh3w�	_#Ǚq�e�X��U�����pX�HZ���M�۶������h��'��NK�����ڂ�
!N]I�� ����I0����ʲl �w}4H
�<��]h�*S��๞�PӀK �}K|W{��=N�!>?�E���y�����-x�X�R��#g�|�i=�<d�|����D�kO��п�Z�ة���-
�Cw���c�,��sѓ�DXr���^�;*�U�͋��֥w���=�G�ͺ{���I�H����]���g
53�G���a;�u�4�v1�㡜���k�n��h�7��t'Λ��ڌoeJ^Q��ڴQ�o'�j��'����-j�e�O&!-����[Гݢ,<thy�{�* jt��i�ۮ6R+ҩ@B��J�4��Ҭ�
�t�����&�PZ�ϩ&2�F|;Wk�f�&gaZ�4{�(%�^l�/úS}��8���9w��y�ŭ?S�@��MT��i-.����N%�+����B��h��j����a�H֠�c�&5��lBY<�!ݘ-�?@�����|��:�ȝ�0�M���x��E5:8)�l�j��;h�G���|i�3�;�i-J��Z^�~Jd�5V2���H ��������gw���U��m���7����9�I����'8�&��V���f:��|8��`ڟ�f{�-r����Ŭ��c�s@�f�ƌ��vn"�hy��U]�ZYZr/�aw��z�Mf�`�Q��T��m((�0e:L}�{���E·����K�4h�ז���Ւa
����x�O�Z����*�<ʌ��.D�J�5 �nX4mOw���� 9���M2�����E#_=zŕ�)�(�TD��=��1ȫ��>��B�:?׆_0g:A[�]�A��+���gUEw�LL''��l��z�ǡx���/�	K�+�TG��!��a����[�nz��:�m`.�q��k���đ�m�a����3C��Ϧ�~7�p&�Rܫ��y+Hʿ;������%���_Z���x�Fj�7��-4���z�ā�G�C�!v����y��i%�kQO��䆾���u�VL��}?|v����F	(V��9A�+[��kn\� D��,�bybk:'���ƍ*�����m��L�4\P@0���%'����FQ��t2�v��������D�<]��� �{�^��i�׃Y4ƥ�q�4�=S�������-'���V�;Qs�O��4w5� )7P��ύ�m�[єk�l���&�Չ��{f:���(�F�a~KA���#}�����@�N��Dj���� �G�K�^i�[B��`�,.�{�N�ă�k(�ƵUo��,�k�?��>�?��aT�U����D� o�=ƣ���aD���-ޝA؅t�%K�����,��ТbAw���bPp�&[5�u*��>@ة��<�V��3N��wo���A.8�Mk!ufP�t�=qj��0��\(cO����-�*r�����U�R�,��L'<�'+tU+�W?*ݎ���`}�� �� 2g��������1��4����L�	]��c�*n.��{�0����ϨL�u��bGN6b�e�3�`�;��)�)��n�O��y\c�Z�3L}��5�����(
�*h�M���������7�s�<o��a6my�26Zzb�c�{	�\����*��|���$(*Ńb5��y��a4-R3vZ��i

#��ͯ��&V�0ʥKCk��^�j�D���̖�c��)���+s�(X2�%��d7��r�F�d��;S���<^�ӟ�f}�;�4����Rw-�����:[�k���朐�>>^�����A�]�H���tv����u]�g$�'� �5�/���g#�k/�w�����V]�ZD׼�y�moTq�6�ݕ�«8�[��yWi]���
FK��{�y(ɶV �uN*u���Ձ	�m���t$�Ԉm�w�Gdi�	�a$�u��9}$�f*�Ϟb)��]H�STM����3�G�ۓ�WiQ�����f/Oc��ll&��E��`�y�N�����OK�.��Z�A�X ��$�g����c�)3|aH�*�7�a����I��OL��l�tI:Ѝ���I=��).��8��������������7�O"K^�^�l���|[Q{��:��D�A������0�2���p1�X�2�9���ŗ���'A�3$��
��QU��ۮ�q���zk��Yc���%�ZO������vY���CSۙ�%�_���s��S\?���[	4��R���q[#�G?(/�3��G��$�K ���$٧�����\l:%��<�z	Xp�h���}�s}z	뻮Чx/�}���t	xV��˃��K�
��l�͇��M`ˠ�����}���9*�1y	���2�K�!���C�ߛ��j���V��.z���/�`����:4e��s���:}"_(r��غU	�?��tcE�y/_\���'\5c4�cnd�����R=$���X�T��?���΅�$%o�1SWZ?m�P2���D�'��8/��PK   �<�X���]  [  /   images/cbec1558-c992-4de5-91c3-4ac90e5ffec0.png���S��i���S��>�����TJA� )��:��8I)�����Ox?�������~gؙ�$���@ �����#_>z' �1���<��K������������1I�n�g����q�~�����r��q�?�g�����VS1*8($Me�^]9�{ؐ���D7-;��ݣp����ԸT%�Q���%�B�ބqT��|>Z::o��x�A�4�3:߸�(ep�t����� ô�r���7�][7��G�ч���e��Ӭ��P����?�����dޏ�+3� ��O�W���U�����{���R0��Y��,��.����/ES�X��㺐��7���ZO���qlll_I�
XZY�ɩ�������/�?�?Dof 1�͏��>5U6w8��&(�l(�K��*�iyH��MU29��=�,���N�z|��;"��sQ�\BJ�<P�����kt�S"�*��ǘN�F,#�O}�T
kO��0?��s\�#������k(��u�д�F���]:���	׹b�w�)�5��b�r���D6x���NT�n�O��r�f��a���������JR�1m����СUPJ��1�6_��]���~Z���.����B2��Ŗ�
�S���Pp$q��%�O�k��[�ph%T�v<=9M#*����[2��}qA����h�!�0TT@���IC}o����	��� \Wv��v�霾�n��G����H���ե�ہ,2�D̍�Mhq�p�A�c�.P�~�ϛ�S	��E�F�,��J�:��@�EA�=��u@&�I�5���o�sg���J	���q`\y�#t+K��7��&8&�s8��$��ag�bY����L�:)p������m��9QG n>wU��	1cYNoqc�������'9����H�o�����(�:��_y��YS'��K��($H�XJ���Ox��\0Kr�DF�>J����z�?�7E�:�0������If��'S�6����Z��j�)��qZ(�>Tѻbz�_�J�K��sX��7vF�T��:P1������vf�C�a��+��,dK)�#���@�dy�\�ͫ2��zKB���\�,����2r�<�_u��^�U*�!��6ut-w5����e	L��)i�KG��I�L�r�S���`8?E� xaaV]����0���k�\&W������s�ؽ�*�-Y��U�=Z�����[��}�xOy����:/�P���r��s��+�w��׸�b�bm�F°�(�hj�l>b�S5��)���3��Oo��/?�?]e��F�_4T�R�0�}�u���{���iѱ�2=��CS���rLm�w��TA W��5^3�>����w���bܪ����%y"Mj\�2Zim������_�$�p������~�����~�:�������׉����w3(M;�ᬣ�L�GBҗVp�i�>�V�\.���e�êJ�/-{g�>8Z�w��E��O����ȴ��N$
��b��~���z����>P��לq�И*��L���ka��BƷ�'���̰1�W�)�у��#�|~B5w�5lX� �2�߬Bo8�s���h�I���ٳ�Dՙ#��?���:�Қ��+&�6y���hk�[�f�m�b��=f�� {�q� &�
ⱊ%�Ɋ��s���3���ט#�HA,��Ӛ���"�~�8�����#���q͞2Oz�Jg��`�"��*|\R���|dÙX�z���Q�Q6|��6��𱹻�����=�baf������������w�� Ip�8WB8���9��Th��ې�<*Z��/��' ɶ��7����d��� S�//Q��O��e�O���ā>y9+UJ!E�qg��:u�����5��{�������=Ҭ�Sd�l}*V���݄����aQ\���P��jO�+���3BѰ��:Y@����a�4c���ys�x���e���{ⲳ��n�mg�n#H�c��A��`�^X+����7KTVV���(O���熇�;�6^EB�1Gtaq�0J��m/�74+���%qF�6
�>Y,���ϟS���b P��O��D���H�;/ܗ766�m�p�L�a:�u/:*,$�%#���De����L9�a�M�ۓ������DTr���������z~>�s��͘.�[L�����͏�#�	nb�,i�3���7j����j.��v���5���WB�@��f�,��,rc!�?��αuZ�w]^9F5hC�444Έ���5���32��8Y�����S�l��[Q�d�ǽ������%� ��N������s��	�����21��33��#gg�CD^|�y&ʛ��E�:�e�����T��8;�K�;I3�IF�d�-gE�ao����z
a;}{rrrXUU�ܦ(��XFN��<=\ٙ�+�\��q���pR�{#&&��������&�M��� U�lv��όD"�!� �z@A�N��Y�j���_��^yz�>I:5�3�'[1b	�3fiJ��Wb1|�J=���gs|���"VK��II�p����w`[�ۍ"n�a�'�^s6����+�-rF��H��{���u:��d?�`6�l���$��`�O-5ޣ�w�LyÚ�t�e���ί_�����0?d� �n?ɦM�;~�}�T���-.����2'�z�Z��zS����%I#Z4[)���AR��-�j���z�/x^P�|�IR�Zg�5�ҏ��S�w�����Ӻ1@�V���D�JulM�z���>2Oo%LX+�IkЏ.��,��v[��0]vv�z�{$���P��_
�j�Z ��e��D���#�ͥj�oj�z/����6�$��n��܍p��4�D:g��'/�Ϙ��h�����f��[�We�\������N�+a�^�PӸBbXE ,D��*UPV�D} ���L2e���|�L�5:�Zjim��S��F�,F�E��w�B���0�ߨ����6�K���MS��:� �5�A�__�U!H�d��q�����1�M:��b]I�svVs����2}��a�7
;��y?�7�����n���Z/�Ifz��݁��/�*,5L��@n՛�"rT�[%��Q��}MpRG�����Qj�=1�=����'!��Zm��5���������!��U�>�#�5ߥ�(3}O��[�t80� a��P������-��Pd�����Q/��>O�\V�~��v���奦�W-u��5b��Z����1�i2�s�/_�P�����1	G��ks�"r��7�%s�jYL����_K�C��ɟk:l�����Ù��sP{����B��	xkJ{E�Vn�ί�_�4Q�/���/�uY���c�����cZa,ǅY�-��W&��]����*�n��Q})뵠�-+	���ڠ� �"SS���	+�"o�o��{G�ɛ���2*+�d릑�4�Y�ɍj����?KO`�Y�
���p�I���@��߄�gb����9|��wSp�?<��=�}�:��d��S9Փh±�Y�f�2S��ͧ��0�2�ܚN~�|W�I�2��b�PU�5�~��bm�F?�	-�V�zY��.\��U�S��veZ>��L�k�����������is��^��.���yz��t圕\�H0�3A,z�:~�Z�4�5*��Z��¥�������(;c�9�V&��"�Aq�TΠ�?��,e	��i���c�-��¹��*�x!F��Y\K��1�N�!���<�ۨ፩�6��4��'����K]Q>�<熉w��V=}��O<5��.ˈ}�}���y����b���Љꉌ�rdZ��.K�4�w[񧾿vf���pq�]@�e�me���3��޲G�zCBc��6�J=�|a3Ύ��$-��`9�w	��uT�0�����QaNMm0�H�5�[��DD'��s�!�����j0�6�ͫW;��YՋ��ͳ�ɂ
���a�7r���n~:Qفs�YU@�]�������#�o�$��/�Z3by.��R*��w־s����&QU���p8<
�S]GW��7j�Miˏ�-�/�:��?��Y&���*�R�̤�v?=;��В��	�JHHX�*ڍ5*�,j-��� n7������1��l&ۿD����Y�M����F�a�L�_��=$�K�b��Չ�}�n�z���O��E�@][��)�>�J����<;;$e���3.#���Al��ǿ�0���J�;$���:j%��'5h-�v ����<0	�4z>��e�r�A)]m�k4���[p�~{}Z |'>���#L�jll���W���%73�3����L�ޫ{YJ6~u��0�L�yq�(�,���r~�|4������Pͧ!�/��#�$XC�j
����o��(A��n`�ʳ��*
���&�?���Gs4]o�t9�	��zyOH�ˋ=��×j=��Bv���&��5�߭?�:	�� �� ���k���i�L�E}Vn�Y����ϗ?��'�Vo����{X"���BM�c4��(��L鐳�@����u1#>ǧ�Lm(�a)�RXۆ4�/�~S)�
Q��	@ӱK�ISe0�pj�?��;���fS}(�p�?����O��Nl꺲�ɟ�U���֮��6C���3�p�v�i��8�����p��)k˾�Iqc���O�	R�-�dy��k���!���T�tI1�LG�*�w��)z�]y
v�\s2<*��bA�IC�.Đ�����	n�!�wd{=����ϰt�E?�<R�w�_����pE�Oa�T� ��6]$r���^������)�~e:Y�&_� ϏH�,U:��`��@-�
���Fӭ�M*m�Z�X�Ž�I�4�C���b�P�AR����.�=����5��I� zÏ�=�"�	WNt�5�z�L$��Wn@�Ḽ��K�+]�_�"Ti�_-h2�
?��(�K��0�JG׮`�H�r����bGu�#�J�TJ|Ww��8\Wj9ͨ�~,I�b
c���M�Ƒýaxh$(�6ģ�|?"�l#ļ^�w�\CڞGpV^��X�~ۯ�	��.�);v��ZZ��(��ZH}O�y��[K��>S�垎%U�!t�,�PRjg�����#�pn3����\זM�H�"w�?��&nqt8��p��)��W���L�p���up-������t��	�ęշ���$�gP;i��C��u��w�OKn�S�W:k���~�4?#S-8<2 �֟\����Ӭ��=�D�>L�W��h�����@1�PK   �<�X	� .W /   images/cca7adb9-3a17-4e0c-97e4-0d979b0e08a4.png���?���?��*t <�H��F)�ӱ�ϕ���3�)	!)BH���ͬrJbif�Y��m����>�>�?�w��vQ+]��n���z��47��}��]�=��?��|'&�Y
<�6�m�xD�{����G��d���v��X[�<bhb����C ���@����?�P	|��֕�G�����a��vpk�\Κ��o�Ğ����#�N�y�.$��}�lЄ�ԃ!��5�cm-O���577�5#�-B��N���T��?��������B���\i�H}?ҿ��T�J���s_	�����x����M�j��5��.' p�o����|�m����7��I�%�S��nW��369��o��fF`ټx�ۅ5���ɷ��:�c;�N�n�;��c�P@�ɨP������;�b�+�.6�h��6l����]�_�e��U����Zy[&�K"1 �޽-�d�U�hT��wB@`�:�d���ܝ�!p�*�[����	�[K��B���b�������+n�۪�<{�joS�[_�]<��%}p����d��kw�=�w-���G��O���?���}�Z���fsc3g��pD�?���+�gD�J$5���+��-��d�;$��IQ:��/V|)D�d
��'�(]|{]����1��1�������zn {�wQ�q�wo��pF�֏-`���i���1���R���Xl���Dn���}�s��o�\:p��]�����������k{�/���������3�JǤ_j���.��z���q��5���c�e`�}󦴰�>����1���B�Îs�Tlo߮N00�t�έ3g�Ω���-|=qD"C��~��X���]ݧ�ާ�VW��K-�++K�)���`�0Ԧ,զs�>ɰ���?������(��={D��J2��-'RWu~�� 
n/p��#�ܹs�2"e?H�}+�&dg],wҶ��>F@�w��ָ�:h�ꪪ=�ҩ�?<z��|�`��fz�>LO�^ԯ�
<����p)M{W��5闯�Z��ts���)I����ٹ|�Q����6�����}��mIK�)�f�6��\<Ǝ��T�[H;V��8�$����|ODͼ���������O��+ӽR�**�>>����]���6N)�*3{��t�w]	�t1��_�׮�SR2��}o+-/���t����ƥ�ѕ��p�M����<}k������5%x{F8���G������T�$��Ur��1����Xc\�U
��:c])OHh�����Ǧ���˫���ӽ��<�*�|
�Y���ˇ�߿[��z2Àw�h��4�tt�Xm㻰]��_<z$Sn��������C���^�X�F^��6vve�(#��h[�5�X_ۉ�@�'O5��^+[����ր@�����Y�)�/�܂�,ufM�w//.>���UH�VR�ot���8w�d3��[DN0��B)<H׹���V���w��Bz��87�����I�	�������R��+���U
���F��8�Q��K�~�4�>�8�d��a��;7��eeyy��{��'��<Z&��i�&&�������KOOO��m�$͏YQ�tIK��[���MQ�/X���$3�������4˼�t1�"jڏ�k�K����)v�������ޥ;�	�,��#���L;�;Vi�nW��n0�Y�u�>���o��bkk�qU-�Q�dfn��o�&������di]8��<\��xKS�tNT�'��ڄ֕���X���7�2E������t��������kz�1�Is�;�� 
�k����Yq+�c���^���c4��C����:����	������2R������p�=;�
�vqH�h� Ӵ������B��b]�E�Z�L��7�I��*/r��ijj�bJm�Fп��z���;��T���m:H�&_�1H�m���������i/���NP* (?(Լ�������з���_�|��ȣK���כcys��f²C��z�HN�����$���=�t�J���ʲ�8B}����O��kĦR:b�5��9�lj|4�y�����iW|z���%�sl��dp�OII�ɯ_�,H-F���_��ִ�,*�0�(���tTE ��B{m���X�������\��w-=��ׁ��te��o:��4/k��oz��%tL$t=�J�Tq����UTظ q�����[A��D�z��e�Lnd]�'�]C�c�g�׵�W�-����@(TP8Mq����Ҭ]��'^=.�o�ľ[_,o�?�)��!)img��<p���#`����]��b] //)-Mjj�8�<�v��uGGǈ�[%+�YT��1i��v$�[s�g�ddk���1�[�	6 ��6�>�V��0HE&�'�������Fp*�k�����cO�)@���[�7�,+ g#Xx����d�A�U�F�:%�����SCO/w�>��F���'�_ \��Ci�9�࠯[��̱13��z�*a�E�%>�v�D�^���&ئ��Fe�ꢒR��L��/-,�~�k�|��ӆ�����.~:Jk��\f��+�ΫZ!�U`������9:��:k���/����i���<yr��|���"y"B��y�`� ��Y&�4*��p4�d'0�N���[�tm6jȥ���5�^O������j����ޟ�����o=�>�ho����iO/e�����{� ��ܸQ �-I�9P��ӥ.� ��AF��YOC��?�0�SZ����a�'kb.G+S�_}c�D��q���p@e�[Ӝ>܀0���1�z82�]�e��2�����Mw�I����g�R�66��q�AQ�{��8M�{jj\.-)QZ�R��shh��@v�aaa�G�7bb�2s�#���R��K���� b��#ll� /A������Weӭ�OK�g���=���Z$�(3��� W'JA�f��e�����v�����-��]��%].�b���XO�V���;�$c�%_��M,1p�;����?d��|U��xѫ�e�@\Vv��N!�CI�^VbɊ��І�˲��j�dR��p; �YnS#r�>;�����su�z����kh\)��cfa�f?Y�����:���z�[޸�(r�r��<PP�S��_����HF�+����??ֺawv֗Ei� Z7B��Ƽ~д�+ؗJ�f�nle.�
k�~�.�k5?ǖLbs�7$�{xx����9���Խ�M^RFf���W�t�fݧrF�mb�&P��������Ib����![ B����S��+<�JY`	�#6$�nr���'Ws��*���Z�]��G�x9�����{msSR����4|ר����#���-���ȝQ!oNN�KJI�ۿR�R\^��5�N$��4��h}��ek����L���Lru��J�?� ��K<�(6�ɉ����(#�� ȓ��l�rs��wK�4o}sι�փY��!.*:��g����!��^+��-�-�/|������7nH����Ӂ[ۺb���#��O��Ѱ�@���p�� s��q�C')%m�!Iy� c'@ڤ/1���C�#�#��Noݗ���;7eF	���;���	J���7��j�C_i�壡��k��V�}l��y�J��Rxf���f�j-��ۙ���B�+;QF{b�� j�_�dΠLId2z+���j{�h�D�a�a@�J���ܑ>N�m�>U���c��d�\���\�aҼ���ɓ�\��,�p�!=�	�ٙ9kc/���b#c ��`M��\�����X�`nmܭ
DN��E����
��WI�i �!��X���)��)��!��%�o7�V�|e_(��ÆD����셉����Y��n�:�}W�u�h�'i����!�%hk�m�.iʹ�~���F���n�&��������{�޵]�n~aa��/E�Ǝ��|nm�VS���
��b@����|����t�G7�a��t<���Nk�:�������l��f��=��rs�}H�` ��ad���}J���4)��Ap�:����l�kr��מM� 6c�T$�K�8N����/�R�O%%��L��o��m��/=����XT����A
ǎAfkw���sw���2�1��h�h楃*�!3�*��3����`8d���Î_��!�#t�)���l@<��:��T_ yj|�3�QNt�V�^�˗ޏ8�VC+� z	X��ҀB.�����Fr�Ǐ[�z2�B �<���I����"}��n�ΟG`�`�-���Ɍ�FJߤ\�Ǻ�c�n^0<Լ-u��Rǆ?�;�V@��$$�#抓etJ��!�U16�*,"�����z� ���/�1��]���uf��H�H�S5�	|lq��^7�-��#�|=<�o�`
��Y����qk����%�J�ʞ�+Tr�3O�\'+���-8�޺8�����}s~d*3��@��F�gn�}�^̲Ď�ԝ��� �Su�!�E�zK6�� у�_�l�(c�<%�`s�v|s/�)p����f���+�?�+�t����4*R+m�����
圪z�F�^:U���?8�E��^�5lI0� �����?�������X���C�Z_��>c�lR��%x,`@�k\�wL<p`���P����[�By��7�T�\����1'��󷇝�ը����
�ʳGS�d�JtO����#�B)��ϯ�'�!aQK��k��}�>(	�#?� �8�E�M��j�)"n��YX���(L�k��o�)^0�K�*�QC[�cN�D�Uj8Oh�a��d�,�����&$� �!Lk��g��5)y����+b�#ܽ靽F�#�ؑJ�����0r;W+�&>䢪�VT�^٥8�C&��T�����M�Z��>���j)YU��ైcȍ��D��Ĳ������͖��2`� 7TT��=ڟ���c;>'���:� -l΃X�j���T���V�8v����&ND` "EZ���K�P�R�(ۀ(�:̝j bV<2I�}�]�!�K��l8���׸!�������Lf(�^f/-��k��9is��d��+�� P�#�ue�����;ow�? djG�餥ͦ\����K���=;w ƾ� �ʣ{̬�O��f$&ʪ>�8Q���Ub>(E�-E�M� ���-T�������O�����'<�:��W�ʊ2Rl�1M��\:d��!�x�&���	�Z��'�|�d� 7y�kz���q4!W�4��c���ų�����\�!��#:W�U:�w�b��_0�.HO�DfN!.h}i�m&G����r�s.�g����\8������$���n�B�������I)�>��m�����p��8Ѳ���+ �MɃ�:{����S]�cX	l���h���>�q}�?�����;_}#�F|J�v�/ߐ��5�Z�x-4e�~���{�B9�)���J���`��)�7��y���􁍏v8���1 �e����'�\�+3�U�(��1�CX^��r��x�$�$L����d�F��󿗖6��}���X�/u%�:�3bk��<��+e��j�b�`�����+Z;9��C"&��$c\��]cc��"���lho_�Lǒ�
n��ZE�T4����������/��MՈ������j�/�����$���
��m uh�L5g��ھ�>�li�u�JE���VDc�9��u%)%tT]�l��b��k�*_h��Q/@&ϴVʊąnN��7 �����t�wyD S���a�[��~�-C�M����n����J�o��#P�)���!��"BC`P��O^:U���`�M+�̃.���c���>��M���I��<ѵ��Hfz�Kۡ'���t�)d��jΉ����A��e��\��vcW��B\��~�-�Y;�N?`��]��)����G, ��/ �gXp�uNن�cV��MM��)�%"e5��Q��3�_{��+��We����+q��o?�ْ+�c��}ȏ�'~����V�����ѹ�f,veӡ���2� �%�O�Ц!8,/�%z���S�CC�ru#
��--��J���T 4��K��n��>܃��)���^�u��s���\cf��V�T�c�Ui�z�YE:-RE�V`���0"<�J�S�N��r.\�r�)
���MK@. �-VJ�nb��>��Q���Dpf� e�jw7�^����pxC�^Tyw��w5C[y���ٙ+��i�O�I.�5�;w_��
!cX�(/�ExhI�����|�f6"�P���n�H���+6���y�	Di�Tv���@! xP��+_�Ph5.l������d�#cA+�LA���L�Sqy�~� ~��X�w�"))I	=�w���'�������J�/ǔ����2�?���^�"MK�ۨm�4��"�:�Z]"qm�H�K�5j+c��wx؟��-�b��va�<�/ hJؔ' C�r���1��2��G�hH��j��OV}��}�rz���o��$5��u���\S�8�geg����#��Xt�W�K��	�k����իo5���/�"\{"g�AAw T��ܰz/��dLv�F��&��iGM<s��,N�(���W�Z�k��PN����x�M�DC7�]W�����R�;yƽň�lZ��źwBk�yî攅�|��.�_Ӵ�q`}$�p����3�R�m[^�fy�����Ο'�[)�N��](�X)u���  ��-p�.��{M�[�-��E�����lc8M���7V��o�]R#�an�{gQ+ϸ/^�D7�ǻ/�s~�o��1��G\m��֊�h�+�HuE���M3k��_�������S֕"�\[��Y��Nȡ�c.uu��L���E'X�G�������6A��ɢ�;�}���qrqA�ՙ�3~Rth�;�0|F�Zu�KFcnE�S{���]]@%�Tf2T�Kq.ݨ���ϽA�R�*�c����cz-����5�be`��?~t>Vߐ�2�J�|�^��]�[�������Af_�(Q2��(5���}Ծ�l��H�м�?C/b6��2z������:�8����3dxN��ډq���2 �xi��UJc�tr"Tϩ�2������2�)� �E�J��S����6����`
�G��������k�����3?OY�t�j�抦Bdw!��C��4��Բ������*мҙ�0�w�uѷǾ�ZTcW/Z+-�RG)�0< bA2��Z��4����V��r�HAS/��t�gg}{��jnł�9yBV֎�߈�*w�uз��� %�T���J�Y�B(Vs��ڝ����J*�F��V*�Y��3�C�(|CcwW6��~��+�_�z�k�VO�p�8
N`�Ƣ���{B�pf[xF��������^��N��B���N�K�0�a�X8����e���T�`������L�b?ʂP�!�R�<%X��<����.��Z�C�Ѫ�KƧ��Ԣ����MN�_�������V�ǝ���;���]���	9i̚��宯�/���<7�?;`l���^�5�ٳ؁[�;�wJ&�i�g��V��6�?���N]�����vs���G:\���ON`".�cq��z*���<"����ʂטs(��W����6S֟�1N4,@��c��;�>q�8�FK��oC"V-U]��+�_R�qU���5�,2V���������Bs,�r�j�)a��a9����4��#�+
5�w��`���X��TF�Ye)H�8qC'<���)�A�h�B�p��1�$[�W-E�;>�@,.p��]yQս3_��[-N�m�l��5�
 ���c�s)@��o�����\��j��(��thX�{P]]�ǰziq����.✎�'ľ9��Ǩ�w���=ո\�4������0��5~)���!(���P"��� ���NQ��㧻*хV^����P�>q���v����B�̵�8<4Jr��������8���Ve�����d�]���5'G��wG]������\nN��]q5N�~��r?B?��[�iN7����P���!�x�M�~X� �t)<�#E����x�uAK�y@��0%�2~�����Jp��Ђ�v��3 py�C���u�S,��P*��̀�z��f��¤6l�1�$ALJR�eZCwzH �(��}ys�2�*��Ћ��4�mr���9��qx��!�'�s�+Ih����^���,�,LUY�Ĩ�
���ApMEeu��(�nm�4�iv]�����گ>��z��)ۼ�m�C����V����mYBv�z:x0�
5��l�x���`�8����%7�D���'�����b�]:����1��|����ȬB��^�����t�B��<���A�j{�Ys<�\�bBZ�$}^\�P�~<�"W�cK�Q���e|�bȥjk�N�^���v��%q��΋C<FJ�iu�Z�f�G#Vi�Hi��o���g�����P!�?<Y̎
`2C9l@���u?[hΕ��B�w9�@H6�_�vI����
��ؚw��k2=fN�S�L^�iTG�.�b��+��nh'@�[/9Q�lg:D&���K���d�?~¦�
�� �b/��K㸾�����Ƅ���kx�Fr�樴��^���H�Z��ɀ�U�w��C�Y\�t��_��H�����$��^2��1]��� ��N�kv���O�#��E��}����K��kE_��^�*FQ8�ۖð�B��A���
X]�B�$P�qf�'�����{�A`�����?`�D�Tb&���������>[К�T���U~�7����J�m'��ۣ�������?*nE��i�-�k4��6Of�t�G,�Aw�����,>y��R���g��/שMH' 69�g�oǈ����=��a���@"�-�/�eM"�  �H>�ҁ|�81d�����YK_Q�xl���9^��]D�F|�����jxf���_���0m��@ j�[��u�a�P�޽ �!��䮘�\�9��l�0b�;P���)++�؜��������2򸯱1Z�r,���ub�̢�K�*;�����^3U]�f�f�s���RnR:w��l��_���kZ�~��E�$i���Zo��Gl��>���5���%X8���C��&�RB�WվQ�����H�L�dW3b�~���#6W��EU"?���D�]����F�p��a�VsQ�0��fJ�r��#6�����QY��4S7��u=������O#r\'��8t���ANE@�o@ ��X�nT9��g�V甔n���q�#�U��l�E(sڬ��{�hRqy��!��*o,~pO��3)wxR���q��ƾX�q�x@���ʚ��d#R��l�}�I��4h�vƫj��V$����o�8�e��fz6h{iC�6���|j��:�u�=t+�%E� �+��7� �1��N�%`��A�;��B�������5����k��s!GGv=}�ɇ��=w��?��,�ݶ���Y�����u���X����wK~d���0Q�TuGp2��W�@7�PG"���C���T������l���`uu0`�F�_Cޓ�'���%�YV��{<��j�وM�%ɝSV�g�C �?�O]*l��3����J]��zzj?O������RCq��әE��2�V��Q*��Y���C�\��d�@ |���ɜ��u���8����Z��t\hYW̗c:�99��%g@YI�So0�Myl�f��@�p&�pW��N��C��MaQa%ɤs�����hG̽30��� ��������&�y׹=��0�Ò`{�� ��Iޘ^��1�'V�[S�p�5�㽦���zr��Z��K��M'TM~��+��C`�8�+Hd1#�����]a���<?����/BE@��>©�صpjk��������6a�q�𙹵��:?��R�.�O~m�i���E�O�.4P�S!�O���#{-�`��%Vx#��Xz�~w=�J}�>�e�>���$�j.���l�4���?���k�9�����Hh/�!fg#>���z?��^W��ܦ�ks�H�H-}��@�1�9����`f����h�6=]"�h`h�PT�ٲ���n�̇�����M�Y�t��][N�~;���l�A����~9�i��9���D�a����M��>�]>Ɏ�TN�m"Ph�S��јT���_�;�ĉ����O��X�LAa�Mz_9�7F�cyT�)_���ѽkq#��΀w;t�	|Sa�p4������H�	ޖZ��+����I���Rr��	i�؞����� ��?�#�|�@�zf��'���K�+��Ȓ��i��a3='��q_J�Z=��V���S�#
����À�1(���\�ZBwhp]Ya��Ւ��h�h��^�umL�B���!��|�9UQ�hQ���@�Їk��a3c�bW��o���P�����ݡ��Ǥ�vK F�K�x+H�;�B㉤���ƃ%~�T�'�e��kuz,GE��j�	5|x�F��q�,�"�9��ʊ��L����1`|��_ �����{����J��߿;?�j�:*Z�ܽ(~����@�0��"�ok�.~��x�#��a&�x�imkA|�����U�g(U�i{���f���l�Ro���*+)q �o{��2�y�Ȃ8���q��{6�`�N~_}Z�Kb)�-��%��c�J��ݰ� ��ϔ�`	M(����>�H�2;���p�+\j�/4C�*������k��^Z�@~&����N���E��xR�#(����v����=a)��Z^ZZ���-p��.@N��5����]L�K�������}͆�}�򡑊�nCo�e�uW/Z	�߅e4��l6'1������FS�.,),i�H���c����|ѳ*'�������cm�oN��sM������ �l���"����խ�
]Ot��W���kt��)z�L-� +��0Rxn�!r�^�]���s�zS�`�� ~���;cf/y�_)����o�ɨ��
E�R�5�m�o*��ُ���H�4� J�V�����"�B����� 4_K���y{^�-`�0�����[Do
�މQ�[Ҭ�?΢2��8y���2�y��-	��9�s�b���ݫ{Ӓ�sW`�q��ah�y����X��U��,Ĭ������Dⶸ�mW$�ߞ&D`T��݊�ee& ��y���n�S�f�I���Б��� ��	J�=,?��t�S �G4�?������?ה��RU��ҍ��[������&�V�il����@�֩�tq5�g�T�'37���Oť�si���Ј������4�Г�&ֶ��\]��:�`��w< ,Y*�ژ�ѡ��1���k�z��GqK%�?��~t�Qq�Z�!��q�#,6%\���F�u��u�n��n>т�����}m8y�}����h��������f��G3%O�I����K���W�/���W���KI���ih_*%�� �tv�ϒo����̈զ/G��gQ�/K����:A��V�C%x�	��-F�f)×F�C�&��,v赵BQ�������E��qἵ�Y�p�߽���N����'��[^�Cn2G��n߃�d��8xN+E�d2&��v���M��йՠ=7���T9���_��,��ܛw�z����I��
rT�
^*-���P}��WD)�25�D�#�w��1� I��PC.|"��^�jvÏ�Ȳ<���Kݗ��+#	]��x���^������o��6�����K8�����)՟�O�A���5�w���H0�����0�=wRD����eW�ȒZ-)��0I��@��c�n��I� ����}�p��&)����K��I�ژ�-�q��a=���(^�k�~Cs���tB�d�>*�x_/�7�0�{�#���0;�p3�~0# �c�n]��O	�=Ҽ����T��}���ѕ�D٨������G�XÎz
y�n፫ڮ��\�0���*��'��o�w���O�/i)\�^։�]B2�C>ϴ�Wp�$�Ы��"���X]��9'`�ϔ>��˸���[Ƥ��'���6�Ea}�X�.�,*�y[�D�x�͐%zx�r��|B�;��ޘ�h���q{�����}sQ�Ү`p�M��(�%��{�~0l#�}K����Ls��vJ�|��|�IZ�QD"�!��U��8d�n$Lwx���5z!̹W�w�������=s�n�M����vђl䇏r�]��o ʻ�q��<-��n���HC`�^K�m�&)^x��F�2W�muɇؤ���ĹN9�L�)$#�������>C�>�(�,��B�)Q�g ��^Q���b�X�W���r���/�(��Ib� ��wjo2�wk�_À_����h޻wo� �+�!��@&P*l�*`���[`�?'�T\Xl���TX�/|5��1
5����&j`Ӿ�V(q�a�q��TSթ'�&}x��
k�eV�����r̫���1���Y����.HZ����ւ=�a��t�ZP�������l�,+<_J�<�D����U(oL#�\���=	�݁�ty���o�� qC������L��KE�6��6Lx�"cax����Ԁ�<�>
5�Y].�;���*�~Ի���u���(�yX��1�xE��N5����P��Z�v�Q��HN2�b�&�BQϔ ����!�Ji�~3EV�n�[h�����t	
8�[d��-�J�`#l ���G�}�|JT"K O�j�\�׷��I$�c9m��-��h�6��\ʫ��#��xш��)MI�
��+.�����^��D�y5Trs9 ���U���&f5���`Sr�y�꯳%E��}��9�}y	6a�M����*.[��DgGH~Yy9D ���K���d�!��Q?�mhhk70~󘊫u��ӕ=]��Y�2�##,���|�8���v+q����A�_��*�ثg�L>�c�{l�C3����h�U@ �J��0,�c�����E.q��"�y(/��}�YXCM�Up��8~ˎ��۹���Z�<�{�QFp���t� ����M|�i%f�%��6{혛�ۍvIY�l��*����7�N�!F��0}����K0.�������P���`���%�R��tw(�v@A�eE���0�S.��~g�}�<�;��8!_�R
k��T����x�`��jO���Iss/1��8�}���BCC�O��W}b�m]2�+%�ߕW۸j�`o
���Lu/��{�/�r�� �����-BO��S�0������4@aq��ȃ�P���n�/�.P�v�J�%G){]��t�9Ev��cI��kG�4,����^��v�i�<�����Z[]�k�����Ԧ`��7F^O''z	hD����!�#�������m!����������2ΰq�;��ǧ4�'{�8=&@��K.>V��Um&ר	s�[la�?Iᭂ-{�N�Y?���ڽB���C[�B����>�|cM�'ѣ@�����8���M����Rǀtx;�A�%�ow���~͆ڙ����^~�_L�V���0(�U@�%�'p�G���0�	u�-:_9�h~Za8��!-c�)"̊���M�������:_��ԡ����Ü%�n=R���uQr�*;[�K� 4ԘU ]�g B�I��0�� ь�~ 1��o[�5�^j�F+Z������[���-�v�zm_��S�|˿H�����|�Mvv��U����?ߋY����u4����M��%h��cbaD��ڑa�i5�R��p!���_��a����(f� �-��4x��)6Dk���V��Y��3�*��	��T��v=}^0�o8��ĕ�W�s�@�Ghݼ�����",��X�0�3uq�s������AH�S��e���\�Ĺ�CCf_(W1�:���@R�7�/��`x��V��0��zv;��o�kR�WsO��5WZ���><�J��>�z���r���n�O��y�[��r��L{�U���={b�����;�cWՉD�c�'l���T����~$�eG榥5����7��ܛ�ca��L�Q/���3�'�<�|%J��y[: �!m��]�k�ڟ5��p�JwE"Ӷ�~�U%���γ�IѴ�%������8ٕm��suY*E�5_g��1��@"ZARD���K� n)���瀼J�
3jT����So��b�x�����NBW��f��_:M�u�����b�zQ����I��ƶ�G��n�@�P�M�܎�Kл�; ��c�NO�:ȟg7~��H����p��#.c���s�5WrC\�cε��U�T-¡1uiJ_����];�̨5rtۋ2I�/�l/ci���c�S�;���g�.kl�\d	��D����M��J+�Ax���ț�Q���x��T�{#g�#��-��&��@g�����ڄ�F�{Q�7J�(��-ۀ�����v�~]����d	F�z��9<�p��+8��-��3�Py]�y-���keRT����1�6��/d���;��@�3��A�I����떨{��;.tt�z�\���^�}*Wg?}�xus��FS��o�G�DNM��|����9�_���M���P��ܤбgZЉ����#���������,��4�.�ތ6Z�W�e>2����{�O��<<�ћw,d �u���&��9+�lT�Ċ2�C�g���J��}��e԰���)�/���<L��c6%6�E_O~�b�'�#�ѕX5ڰ8v��� ����he�PS�(�Mͫ����b�ͅ804�SK�&�Uf*%O7),�>�]���o�R����d��-l c�8$  ��{�`"��"�23}�����&�8'��5��
�Z8���b�2��'��U���j>���@�;��ݔ+x���bf��D�Tך��0��y��Gٴ�� �	.E����q2=�)3r�����B������ڍ��Y�r6m�V+p�g�b
x��(�xy8í��)��C�l ����$�aN�Q���o��&$��%��F?q�w��剏�Ii���96��"������%��:B��p��e�h��C���Nv��F4C1�iNZ����l�]�*�،��w��_������ūXa�-q>�2K��Џ��>�U�/�X)ѿ]ɳ����;'g&  �r�r757����Vg�O�j����E�8�):x�ݓYJ5���h�)���C£I<��� ~��t�K�6;�>8>�]O�&tW�pB�+7��/x�Co*��Z�M����Rx3=74MJ!9g�QD�%C � !Ee��\j�Ү'����)8M���#�;���8��ImZڈ�f�@��ߌ��\�rBB��� �nȢ��怮=�İGU&��E�6���jg�ż�R -�I]I�fn�?Rc�-�1��Z�l���N	����f�[�$�x�^����z��������J�@̞}����q���4�:`FIX2+$��0�M�W�hs��ql�����Ʃ=u �ۨ�g:֗k�x|�:�8)%���3�tm�g�,  ������ϣǎ��h�6�y�v��z�"�]y�eł鋓��T�~BW��.�vU2|`^ף68k��������M�����Os5���)���	ăM�[������Y�P�7����*�4����(��b�\od�C9�Gt{i���j�|+`-���P^^�9��~������C�Z��N˳ ���y��N�QpMp�����ֆv�D�ė�y�q����P���ugD=j8�&L'�W��G	�m8^=Y�N-���`gE�J���Un���Q7";�jDv�P���	�:����1@���Q	wR�G��4�9��bq2��(�T�jBQϸ��j��z}N��d�/scܷˀ�Z����6Nt�j���IffJ)����.􋏅�,Y�%\�1.�s���H$�v!�2ЯIɇ�&a�]��,�@���i 0rX�=;`��mL��'H_�h�̘g��i�iV�k�ϨZS�e����\^A��vg-o�
pi��HJoJ��z���$��k۬����z"�}1�2���W�:�B�H�Mq�X�T��v�����e�����}.Z�ݹS�xM������u63py��.::Q%z�{P���Աj*K�J��m�U��@�zm�c	#ɔ��o󟢛�����{�we�mL�:]���8(�������#՝�9�H��
�k��C���2��;�B��7�6o����&����̉Z��f�d1��J���O �����
XZ�E���@���R�R���}y�4�#��xV:q�'J�b�:�(%lV�Y�Ɇ?�?6-�q�!#a!nB
�͌�\�֡_52��78@'*].�S pI���c� �*��s�0���U~a�t4[�y�t��I���%��lRz�.��r��X��L5�ڒO�����(4�^eeJ�q��@��!�~Q)u͟>~�t	��F9�p��'�־���Ͷ�&��`��ڼ!������2�� �pk�0N�4��2�>�7et��$%lmQ���3����߾�e�Z[qi���۵�=b=,���8���`S�{���Qܾl
��5���5��&�hHtlS8�{a^<��u�{�)�~��k�����[K���J�Rܓ�o�sf	7$�����Di�9w
٠��1M�.��0��u@�N�u�8��y��m�����ɴ�K��Ro������. {�K�xۺA{�^kϧ�c;H[����`E�?�������C֪C6H��Y-<��ʿ�ĩ�B�[;W��F�/>���o�`�c�a��j�_O4?Z�$����r���,����%�۾��[7�K
?p��D����G�K��?��h9G�t�����f�������a�B�N�ם6��[��E��z�o�"u�Ț�('���\2��**�z8~Ű�p}n����l݁P�o�Y�$���do*�"󄲝y�YY�J�����=���g�ᜳ��s�?���������<��y���󞀜F�ZA~����$�^V�Aޙ!/?~MN�B{��M��>�I7D����g�/�B���c��~J�-(�����%��b��j�p5Wܚ���N��+��(��U�%�_��Lf<�/��
|'1��:����"J�� ���xԵ���g㚺�}3���� ���m~ F���3q�AlL�>�룈q�s:*��"��5	���v��r��=@F�s��g���o��N�r^>41���'>����6�u��d���0���
�>�)1��u�~;�&��G�B;�.�Ԅ�~}�:���X�}@t�%����M�n��qH�(~`�����-ȧ��2iF�����D�Qٵ+LJk^�v��p��.V͇gB����������r�'r�R�����K�pQ����ߪ�f/�FW�%�#��b���=/�����v��p�=�*%J�d����]��2V�(WyR{~W���7ySH���zÓ$�oG�zk':,�.C�"-�<U;3�&m D��'��	�ʋsF�xm�����O�6��8�)`2%'��j1ؗ=Ra)pW%�{��񦔴��z_���H���fz���-)����0psêV����?~�x�|�ό�`Z�p�Y�u��:\�� 3k@2Z?����'"�䧇���L!e��H�/l
.�*��� ����N7d	��qf��T�������n"����Y�)|�l���h����N����{M�C'.c�$��FY��Ū�����	���Y�SR�i>C��x�Q��9�ʿ�Y81��x�C��8?;WN;��_��������8���}�dE�� Ι1`����ҫ4�'\���-����q�/8������?���B�D����\����C-�K�Ђ@P�oc�ĕ�t�#�:�IX���LA�~��n�;i���
ظ=�uս]Ǻl��
�,�M5X�Ab�<$��&�8�8&
 ����i�����djCg�F�tI����/Ǜ�Y��7fv�>U ֫�g���w�)��߯��`Ѵ����X�@��~_�=X{�`�տ2g���Rk�gZ�����%� ��5�δ�VX2u����`[ {�[H�<S��R�7��L�����%�.0����!�6<Y���ĳ���&Rd���Q��ޖ�_a�uЗVV��l��Ϣ�q�����[�'GY��ܰУ�$�M�H���[��:5��i�SXSG������[���{�`Q�m%�:�R@�.:��OrC<'b��� ,Ac��ØW"s��iIp�G3Sn��d"T�Szz��_�^n�/�,�\�`����A�u�~��)�K=�f���q�9��:0��
Dp�h@���]��¥�]�k�����ӓ�T2��K���F�hݸ����x�㇯����K�&��:is�'����b�#�cN���@B�ʞN����n����Xz�d�����hg󹍠�߄�T:��|B�{!� .>Q��f��*1�y_�"�p0c�~�ԗ! [�&}����9�/sT�I41�N��`8X߰�vq�����h��#d�n��ׯ��C���G|�M=�Bg�w^?_��'�S��Y�ӷg7�owg�6�R��1	}�U��>�=�c=F��t�K��ޙ�k@(��r��1�B�7�)�Sd���ZL�v�"I�|�Y��x���JV��g��ƫ���,����!�J�y�N$�N�څ.'Bk�Y�s�쟪8��tb��)n$.K$������=g!�g��R��ҧ+�T���:E�=E���������m�C%����
���ץ k�{��w���e�n�q�qݿ���;����.�����/���a$S%ɂ���s@��A��݊շ֥?svp:���� �c��'�&f�,��^_��vn-���9�R���밮���C�2ȴj�N�]c}�pP>��Ÿ�Q�w�Oۯx�hH8d�|E@�xY��R�o���8X��A�Uv����F�B�y��_���2`
*��K���g�hP*�d�E�h�e�(�U�We�w�=d;3[�UJ��[\@���.P�wP�V>E��*K�˯�b�n�d,����no��¾
�+��uR1N\�_� �2�{�I��Y��&���b��C�3Qhp�̡����	��3��|؉rvs��x���=�證3O�t8|~ͭ�[%�hG�-����@<���n���\@�������5���ye��!|l�����Q��\<��EZ��ƪ���[zKA3��]���ڪ�רgʊ����^4{�Y�H�h�-�w2SM��>3��ȝ�-���uqXҦ���xvxJKJ��&��X�����c (.-݀ �π�%��?K�u�$B]}�A��x�
��I�.�{��E��8 �nqPx����+�����+�	x�٧kCz�,�_�L�W&���l�H]����cm�6>�a�8<T)QE��/�`F#��1MZ���ls���[���W�޷AUP�v�qf�nЌ�.m˧���!x��"Ӳ_vV��x^^�|�?w���8E81�%�r:�wUkz]��<T1\c6 H_��@Pm�u�W_W���$U��*��;��#jآ�g�gb�����WXp(9���v���ב�3�{_t�ޛw?���{�����]²u�Kvk^�e�oY��y�f�f�|��U��������K(�L, WHQ�)�4���vK�A璡G���?y�^�yc�����A�-�uyl)h%|>���^�H9q\?��|�,�?���-�^�E�� ��.+w��GBk;���U��-ڜ�U=Y�>B#�<W�ظC���h�9$A����:���ς���|�J�����i����2d��[����H&��GU:�7�Jh���o�	X�}�0fܓI1e77�7�m�w��i�� ş�P�W�����w�Z�	34mRs�S��7��k.ٍ�;�%O*�q�HkP���*�cdD�Q�t��f�h���9��ܜm�,��/�B�>==�`��O�K�AI~v`.ds�����]��P��eFV��������{�c�������x���-Ȫ؁a�nW�nX��^w$�;�L6����.Z���}�%[����Q�)i0�{s3^�3�w���-�)n���`g�[����7�����D�&�$�W&���vE������A?��}�5,.�D0�ӫņ��*���Đ�"|�ˑ)l���W��	������}{B4���t�V���R���`���^���5z����A2��B�
It.��6��k�_�RvVW0�w���!Ju�����S�� p.:X_%v�\�3[Â���JD�XxAv즈��U�pw�L%-0IR�o��!���oo��S%%Ô;��K3]����F��l9��ڝ��~�	j�|�>�ڄ��'�����w��u>�FX�p���fַ�Oa�Liv�2!���r�<�៟j(_jZVܖ�Z������J�
~�t�/b6.��^�l��n>cB�(H��w�oO;d-v�Ịˠ]��D���s���8<dϓZQ�I��� 6�����Ȯ�*q���m T����Y)ހ
���1:&�~1�E��;����t��`;�_V�;)�)2L�P�x�9�%�v�+B�cm?PN�������1 �ݢɑ�|��5LM��fK eqD�ԓćyn�RR�a�
��U��ِ+�ܬa�޿$L�T$��#b��7� $e��c��Mx�	� �<���L/��}�B����O�G��+*��׺�BO�M��]�)P�u3y��[
D�4-�Z�g�V6T����������dL���zX��,���� S��<��Q3y<���'�'��e��I��#�ߏ;��JH�H�	�C� �9�����v��X�ټ��Ds^��q��q-z��o�-���Ar���c�u�����䄅{3[��?:Q��j(5m2w�ޞ���Y�����A�����?��4�e��ov"��g*	��U�1.��3�ޏ���l��(m��g#�i0��֕���aM��Ԩ��]AQ1v��5������&j�R��B�/��;<�Z�l�|WӾ	0�|y���	�c�L	MM����F'��ߧ����*��2X;sh=���*������"�Y[������Oi	v���e';�C�^��'G(�����ph���s����[�i��p�(��J�eӲ;g��AY��u�F6a`%�%�*3�-����m���K`�.5ȒށD� �~_.�S9I^�����L���Q��b���%��0.|�O�-_20���;1|�b����?:#b�H�T�f[=X:Q���3en|?"��B
���X��)puR����*���-2��t��g�8�IP���߼ڴ��ay�C�y|jw�QoG�n�}>���� 4��G5t�]�4�'�^F5�����%�I4��g�(T�)��n��@p�V1�%u3�����5b����=ɏ�~�y��w߭)�^�|���-wNE��7x�z�'╺��Qr�E������]o)���P]э�i6�G_%˸���֫��[僮��y��Uj�sfgU�k�!Ł��GQ��ͺJ��6i�x�'���0xz�M�7�!���	o��oww^�;���^�Ų�`f��qa�<P=�R�v��z.NI6tq��8��i.�߄F���2��c/���y�6��I#��ԗ�IkJ���˭�Յ�I��?iT�n$��[Pmh�AhR�\m�^�4�X�2SvR��:f��P�����W���V4ٰ�3=9"�r�D�(!C�������f:����!7+}��0er��=�)@W���%�7���/�6�Y��bL�5��e���V��<�C�B� �Z^�_U��Iɑv��ĥd��δ�v��C�J��$�rI�?� �������*R�lEe}$nΏ��dz8e��F�2Uϓ��re6)����G�h}�;/��(��$�0���B�K� vH@,���2=&C���r�z�:���/oo&o��ɱ��H����-�N�!F�?�g��j��un��Z�.��Ucd�Q�׷�1e͖<����(���.3��{�y�}����A�\6�(���B;�ۥ7u,%�/��c뭼u�b�����K�ͣ�ff],��8dhh��0�h�7�d�e�ޥ��e�yo�Yw�Z��q�B�0Г�hp���3�}����@Q{^SGk-��+h�$.X��[ U;�lk��Ԭ��T���$<I�ă�i��7S�R����Uˌ�Zr���7j�I��ST(y�D�wD�j�~P��jz��jr�V�M``��_�)�.�+WA���]��x������ix����|���ޗ ��=�H�}n�n�a��c���^������7��y��N�P�f�и�;�~φ5�#�U�q5cS���qM5d��&��}w��
҄4����3v��Kw�j~����|��$�&*��<�m��{B�ᆕ1}E��섔��V2v�����ZS�q��=)�X65B_E֚w׈%��p����K���B�V�2�����fi��$�H���4�'�m�N�Γ�v$���Q��POB�9�_��{m1���yJ
��_�P��$)�\�'���L�\��(&�ӝ�}����r�̀��#&�4��i�.�Q�!�Q�;����5A�y ؁� G��O<v`�������`�t�L�M1��TD9�I�7�oEف>����PݝK�|����	�L�iH�Aրy�v�lL	�ş6\��B����Z!ƨ.��fkJ�����U�}ZCW�(e�����x;ݏF�7I���<����k�����4�}�ib�����/;���|2� w�YU�~/� {\J�%�xN[�Q[�6S��[mL�21d~��:��Y:|
Y<�3�P2u�4�Q��B�&�#�ج�w���nX ;�>�X:�cUX��ua��"��q�R��q�9_z���˓K�{?�6�!*T<v[��K��M�q�%%���HP���m�'喢B��~��z��qu����Ө/_8����ؖ�p��,��؜�����������iO����څB�̮I78g8F���G��qZ��������?>�V�(m�$UK��C��P��^M�n�4����O?�k2�,��S��s��rgM�k�������G��~�&�y���N< �G��Rl���wSC]Jc�A���T8C��r^�9i7��I�-�y$!x�zg�<���^'jH�[�u�ϻ胼�_��y�{�k��@{�O�Xȿ��f��� ��4�r��`.0�soV�0q�5YĴi��b��5|�#;T�
�|�<��W#�����4#�y��ܰ�˨�j�*��MZ��K�v��'�Xm�i��.d��홟l���N����{?b'�@0�S>Y��3Z�X�bE��y!��?��Fh
R�Ѝ�7$����=�A��3��]���J|P}��MG�F}}���w��(���IRzK�ГԽW�~�p�?g�=8=r8ڇ����\�6��mNCX���{��A���������d�M�e
�{������B��R�[1@W�/��|p��Z�"���?j�Yd����%���f��̋QKm'$�h�JB@���n��tb�b�Z�+Bi���[���"%�3T�.��u���}�$���*&�7���h[���?��ϲ�7p��U�a�s�����ZnYc���0o�R�����:aB��]� T����X�U�WT�O�����;�m$��l����H�N�~������+6ځ��.G�ж����f����]ώ�f+H��l�� ���_߲�RZ�v��X�C��u����m�Rl��G���6t��	���=����6
�j�#���u�'���,�/|� LIW0��M%��j�b&1�g��6��)�2WY*��A���w��/T\׆�Q%�AlGY(�N~҂���ҽ�x=d�F���_�x�d*�g��M�9�-xA�O����'@"@��>l"�,�V���L��Va�Nۿj�����]m�������ȍ��Ɩ	Ɲ�Wr[��d�qM���^E�ܚ�z?��h�D�Ί@�nu���A4&ˢ�ꦄ�&!���e�K%%敗�F�dU(B-�ԥ�-����d��v	^���{�1m殼��
r��w�*�E����ü�TRRR���ӄ�4������>�a&�|�p����R��aIq�|Tj��Y���.�(/�lu�e��j��gW�%�O3(ޘ�� �P�7Ƞ�K@b�,���V�u!����,���un���U�Z�-�T60nȵ<5����G��M*���xw�)���~�5��k�����!��|��炨��{�����#���Iߏ!
�;n�+�ʎ���_\d��u�k���+����y9_n9E��-�L�����]�=_��q^x�/�9���$���#���]��MD� �4��fY�$V�*���5K��9�*�p<�LU��p��{�즹�'E-��H�dw1�{���6G>�x�-,�GN�"�	Y��P��*���$?�����ۄGH��$"Zʭ@Uc����Mí���9���|W�%��N�*{��{����1����r�ъ<��F�۟���7���Y��漻�T���c�cGGJI|�q����)ˁ�!�A��0L�Ou�:���!�M�/j���ͮ���K��*�n�$�w��~�]�Y�E{��ɵ��l�Kf�t�L�v4O&a�F���t�rlL%(��L�g�:�kJ�i˲�TnB1��U�H�!I�f�5�Ĳ��>-(8��9��D3��pf辙~@jꞢ����bZ��]���� K�Y����j�7�K���l\�^BXl�<�:?�܄N`������!��P��D�@������ڗ-�]��l��7�(;�C^5ӈ���jt�:ZƮ�P~I����;��I�]V	AZ7��-�:��A�%t�n[��Pꇩ��K�U�4����o)\���z՛�2$��px�d}�1���Qt�w��i�RvS�;�����ëqgj�2�Y-�ʘ����X_j�f1B�޲�̭ �0 BN��-��h���T�o;���~��~{���C��ǌ��7�x���%0���K_�����-3�N]_�tr�ٞۍ������P��%b����V�~�Ұ�R\J	�o���|JaT)�E�nSFc�.Áqp��.�H�Cr���H�NK��z�^��Ɠ�=����$Q�3E�+��n+�e�IC�f�
�����؁_Ơ�o�0?����p� ؀���Q1�O�/���0��������s�ų����>.���׉u�=��\!��_;8xoL5��G^BZ���9�����1��gW������t����>�>e����YM�A�JJ���1�W�@�҇_�����j�ꫝ��n�e�!�ٞR��V��\�
5�o�y���Ɖt������a�s�s&����
���	�?-ģ�hq�?k8�L�$�0_�Ů0G����Κ�.�F�BR���l������&�F⡿f�Wr�H��A��a��3�h	����
�z��ٴ��?�?�/��{wX9��t�T��I,�����5�n���ً}�Yf��+�/W��Z�6䦨ku�Z��ٍV�{�j"����a۪5��w2��YfJ��}[�c]�w��C��c�%�gh�~����G�;`����D�-I���IEZ;T`B��ؔ�ˁ��4x��6p�K7��E^`E���R ��~Q�\�#Yym鸟�g}�>�h4>;H 2���2��M�$f�u.�I�ܥ�Є��� ���1���/m�F%-n)՞��}������py�-~����VP�;mv�c�3��	�|v�l�٪��N%{ad��s���:��H���5���Wf�Bv 񋎗+���R'A�F����|덃0h��&��!�f�Ys������.�֚|
�Rw\�]���E���޺Q�ڨԡ�=t�?���n��I/Z�= �`�����B�L�c��A������6)������wk�6&�U�TN7����V7���f�u��+�:&�v��h���?���)��/�$?��T��e��_�7��-�(����\T��gC/ۏ%��k�����a�� �b�,�v#*{XX���9�	��I����v�D�A�5j��+�����n%?�T�V\��2zj����Ņ��;��*6R���
���+߽{�W&9n}�|�X���ms�s�m-��3DR�Ŵ`�:�,w��~�a�o��Zo����4�ޤ022�/�Vz]-��8�tj�j)���d�+����<f�N{��6��2ģ�5�RGO��<���KQ��C75Daۙn�
�s2�e��b�t���"ڛr�Q�a��yN~�e�N"����l?m ���q=����?Ϩ��|q�Q�j�����&dhڽ ���UK� �3��1���J���|x�����h��8�i������¤�K-���@����z��%G��Ŵ~��������Ų��)Pxl/=���5E���E<Z��(R�/��7y\:|�D�$�S�R	QԐ����%����<��P��ȼ5W���ˆ|@� ߊ�P��(µ.�dĜj�H���6!Z�g����,-�]���v�-�M�yC��$a�>�(�%}��J�/�" "$�/��K���%��3:ޙ�kz�r��݄�IH�6n����+�Ɯ��\D�"�Z*�"P3�ꠖD�#lŚW�� ��i7!k�P&����=B3�Ů;��Z�z&���U��Oi��������6���O�����3�1��e�Ջ���K�G�R|�iC�zY����DHӺ�����<���6�_�3�͜e�Ot��FTޑYr�?�᥼j5AW���6!+�P6��|��i8�q�����3G����˿gm�F��ڣW[�}�W,����~,B��`�;ލ��b�M��.uQ	��z�!I�J�U��>��b��b���d��L�-�X\�w�����F�q�Zٽ�*TQ��a��#h�8�=� ���dش��@Px;�E���c�hU�M�eB�����M#݌iDtvU�F��7���PZڔ4U�.Gn���A��HA�#7��Ko�����Y�d�|�wX�X�z�v=ݮ�(E�����X����)m���u��>��Ekv����+���ZMM������ˊ�2���lS<!<� �ˈ}�����ђ�4��40}1�C|��SW�Z������V��sAa�Jbh3I������S�pMcBz6g?qo9�U���M�_�s���i��!���W�@^c�5wk��x�덃]48� ȷ���)���ҡ^��xD�K�ܨM���p��!Ğ,����3x�[��ݟ7B�?7��[1�w&?��������G�WD���a.f����o���u%=��&�9�4y�^!����B~�\�|+/wg"J��!O>T7�j�k�,���5����1]p���Z*RQ_v>5��������͓��_��痣M�Uƫe�C���s������v�S�`�>6��J�)�$."�pc�+5W!��q�~&�S�����G��3��4˵���\h�c.t�q=٥\�8C�ͫI�E��'��}�%��	)2������Xz������˨~�1����[͵����
o[6�&\�-R��:Kx�K���ucͮ���v�!�%^0�F�ˇ�,�C��p�{�h�{��W� `}%o$���\X}�j�Q��q!�̮����*-��ݕ��|<�*�� ����F��k���������t7��2mZ�T����mNW��e&�� ��ӂ�Q<;eo0O敨�5jSnt�at��}eFx5��r�m�S����1�ݎ=�N?�c+�n��]��
&[t���������D�y�L�K����}�(O��VL]d��MY��*�VH��a�Lɒ��Vm�C
HH��GFbG�+��pje�n���Q��B�O�'t1V9x�O["�YB������?|Ƨ�(�Zd�P�TU�K�ջ�� _y�w��ܑ~�k8�iGN��fu�j����.L�Z�S�ah�*�nK�R��UM�_F���N�&k�	1B�����+E;��^!(���LJD�P��k!Ty�V_�q�].>���-�����l�W��#���`�J��?��]�r�1'��X`�ύe������ ��� �~�x�)t"���#�n׶��"J������-�|&��R_�OX��u.5�;��K�ֈ}���YOG�{�����f��G_��\)~â�t)���Ag���UO7k@�xX�,p�+�+�&�p9�j1�v曕������+S�h9~	u'Yc�����[����׶W^�Yot\�QL�ZKb������
b=�gk���;����п�p���b���*G%JB���	:F�VL1�S�o��/¥�
��څ�m��������6ۗ��]IC+����6�aZo�S�Z5AH�����fA��R�y�k/�6�[}��r�
�2^��˒�k�#w�	ǭHI&�g9c���4�	zv�g�{6ϳ<�q���'̷T�B��֗/%6fOq��ٸV �z&aX��]�𴫍��lꪔ�I�F��߼M�]A��y�&�U�jE70�"r>��)����u����x,���S[��g��X��OV1��G�7�k��+�.8mҊrQi" �V�(��J����S�����Ѥ������ڙ����E�"\zض�ޕ������������H��캪W�d����ֻ���&<s�fd�40��}�C�ᇌ�0�������3�RX��/K#�K���A�ۮ ��|͖b�[!.��|�ZU�H|��Wf�q$�U���<9pc\V�ۯ]m��>iߍ���e�;�m�-9�����V{9$,���ɓ^�B�Y*���]����W��n��{����v�CDpZs}gz�H-|���T`J����w���V@���(��N��,���jo��:�BE�L'�^]�����L���
�-�>4�iZ�"��_�-4ω2Ly=G-��{,[��c<�Űl7ĕ��� Z{		��v�4d��d��t�?����yף�!�OP١��(Lad��pv6\|�3;�\|�e|��1;*�-jX���&�0�\T5A�8�iEۊq8���ę�x�Ih�h���d��y�x��e�o�ˬ��9῎γ�;���J~�}�9��-�2h$f���.����7���	W��M�jZ�`-RV7��e��ٴے�l�5�O��AI6�K�)n�R`��h�V�@��9�����.�"6|4�0�ܗ�ON}ۼ�B.$�2j�<���4�\���h~�����eQ��R��ǟo��0r̔�Y��=��;%�v���y+���QK��
��5���A�{�����Y{>q	|j<&1��6�!p���lO���,5��[��p�N�ǫ�t~���7��wY�C��X��:�k��*�h���ߘ@jNl����ƀ�2⅃5���`����a���.m��=���'5�m���K� 	{5������I���.��z./~��I�Mt��\d{(����=�<��[+��������O��r�F,p�[CC%�q9����O��M�J�)�'X�Q���#4� 	���6��E,%��Xcq~?	�Ά�a�Dz�v'���v51��p�z1��������TD&QҲ�?��e�0�	J��q�	�Jv(:���K��]j�Ĥ�c�A�Q�0�l��u�{�v���f�V�_xJ�i"���������SOZe'�iܽ1�dJ��dH)��;�n����9)��d��'��,��!�_`K�a_�� �԰SA%�ي�C(zC.��:E����}f�嶏v���Kc�i��>z�;�$�2�%��}n��dD]��5ف6����~�^X�&"x-$�����ć�/�)��ko�b�����g���J�0 jŚ�adfO�Y�MN?����)�5K��Wt�(I� ��z��(!�:�@*��~��̒b�hY1�;�MV:�8N.CM*�Wy	��讟s �����ᘧ�9�P��d>��X����x�"+���ֽ�h��Y�P[xS����_��O����O�X:p�����&��O�����k�<cf�;����p���aH�'���{0r�4V�F��S3���P4N�ey�^������'�4��M�R+F����k�,����_�k<l��/�?E�0����'L>���JW�U͒�6��� �����U���������{�|)Brފ��4w˓�������$\����'5w���K$�mnK����� ��ᖵym��|�D^�vME^>�|�4Yb�wQ�/�״�R�_������1E�<7r��ttu�4?gfZ�N�V�ɿ���1������Gޞ�_��X�;xos���	��0�=�®�C%z�����#s�鋎��w>(&}H������'�t.��)����Zr�C*͏dJQ>v'��1h���[J�Lm�w�˒&iD�G8?�ԑ��]��{d%MCܻ2X�����zB;��������[Y�N���bW�`�̊���4[��e�)Y[Vş���x��ٻն��,h����JIEh�A����P��POT�
U�JHr���"�G9NUX(���3��|�?��gQ�A��A��wT}��O��ْ�e�A�SФ��/�� 2����a"�NW[%V��f�^I��(�|�^q����/�iEyAؤ`x:�rÅ~4���&�6ۛ����� Y2 ;`]��vrf�����d��b���O��8�e;�h�B���$��<ԯ K.>���|�!�����M>�a5�����A�i������J�f����7��H�a�(������!���ag9���n��	z{^�~ɰ"�gP^���;0p#^~�H}c��iJ����nXy܃��{Fy�i�4 v�u��?��/���N����O[U�ͨ�'1Vv��4�Y}u��?�Ѝ���M~T�h��D���5�6��zi�1=s)� ���p�q�}��I���h=H�K�4���١�X�� ��ύ�J����WX�~� '��@[UDx�����:nZn�$|�A�{�hH�:a���s�璏��w���,�*;����l���׺�.��&I�/g�pѲ�o.�P�,k8�Y�JP�錄�V�@]��Ų��VK��T8G`e�&����oIs�X�'S:H��CzT�6	�Yg�[iZ�}Ƀz��0��2J1�H��!�ݮ��|���{S��=�v^*�a�XjN<�=��d?����F0��v��$ئX(����:�	|�6�9Q.���0�0UpD2�7�Tn�6����� ��:rnh��8��#�o*��&&�����V�gљ��c�.��F�([�kp���p���-b�<z����5U#�������e֑R����p>nO:�n����?;#!Rʛ��H�/�g�՗�lώ�ΪH��(��=�:������o~���H��~�v�U<f�}(3=��k�3���Q
��b������Y�1R6�c�HS�x.}5���٤�߬}��$�:;m�g��6򵆫�u��Q5?a�F#���Ԉ:�T��#҉��d��(v��U�Ǝ�G��#@��5��C��ʺ� S�ma�V7�0��8��i7�Z������_��-�+x`�׎\� Jv�eb��v%aR.$��b�����`�5��
)�71]HS�y�6�1��2��c�mY��}�p���V��*M+���r�Ԥ�Ν�oL+ɜv0��]�ᮋM��ev��_�w�n~�zJ�����p�̊5���OJ����J[�]��
R�L�X��" ���1�B�ѿM���@�_K��H{��ޓ������M�V���ns�k�`��[l�n�wȹ��i]��(�d.w�ne�-�Z`>�?��)
�L٘4��/��:��#�L������� �L��J�{�nU�*�(�T����Y`��㤨�gP��-]%0�U��.��m���c���hǃ3촡6�%��Vyp��{�썙��1XVOf��z� �Q��}O�5�K�����hl��À���g�աJ�8x�z�
ݧ��{�e��??="!�TO.��k{�C〡(ś�7M�q�+xd�xV�j��ߊ	�ʬ!�.K�ɍX�~/��������¥QV.#�����Wb+r6ז8�5¡WZ�3ydc/Z���.�(X,��K5U{�<�ACTq����d���7�_��J�xiC8�����e؆�R]wD;D�#�MLLD��4��!�r�U֯��J?vZT����b���y6�Ĺ�l`�MW4^"��������$�%O}Ƃ���O�\���߹���4��7�Wd3N�P��z���!�t,/�!�NM0�OM�_�Мowm�q+���8�`�*π� ^����!��G^Q8��O�j�eR���P�0��^��qԏ�l�l��G5اSL�0}�*>���֪��`�-�Pn�����4�r���0�Vs�
ߪ�@(�Ө3�
�%���*�]L�ܤ#���K���+��"�xh���oUֆ>��$Gb�I��8�CQQ�y<�]f��x�1�L0Qt97�9���/P�TzY]��ױ�$q������/1'�r��Z5���--��kٻǐ���ZpA�Z�������f�}�ֹ��|�xe=2��0R>�n'���L�J�4�^]Z�"�*�\���O�30��JΠh��A��U�Ț�P!���솄��IƮ�#͑f�G\�����c����qD��փ����Z��fll��/ʐ>�}�G����6���ϼ�Q	�.$��7�_�h	e�5ܪ�~g���;
x�A�0�dĭ�p����ˮe�oQ��O�FT��z��!�I�d�HGԆ0׆��k5��»��ՒdmT�c����6�E2ɻ[�A:��䟸]���Ipj�x����p�M��~�F��X���-e��N���rj�n�P�'w93���c��U���x̲�eD$�醊~^��a_��^y`���\��A�^C�տ���~eX�N_a����и%Sa����o� ��.��� )�5JB�X��o&��˄��jy���|��^��{LzWz4 ��C-����/\[� ��Y/����?����qO���w;�%�VMF{�G�٧��+�T��� 4�� jG0�1��(!g!{z�I�Ou�3��-�Tzt=w[�,ݯ���ފ�!,R�+��G���[��vW���Qs�L�1,i�;c�K�#s �|��?@MkP�Rͼ�"]��'��מ{q�1|��u��7́�$F��+#��q��v��9s�K�I�����p�3�ǫ}pp��/\�K �)Η��������	LZf��L:}�v�G/��n�����|N!{KqTt�o��j��В�3�	+em}Cu��A���\�L�&���~��R��`��+3�r~E��GL���:�����]�_��/E�7�%���pY��a@�P{�b�'�ц�m6�a;��Y����֐S4�L�Z�3�m�Zw��ܑ�hHH'���Qb��m�ͺa`u�@���W#�32�|Jo��sX6�9�3��&����ox��.�^Q�k5e���hkӤ�TVV�Qo���������t��H�4�Q��� �)��HKK��0b�(-9�F7l4��2}~��u��s�������{�p�#��ߦ+�(U�����c�������7���;�#v���"�1�Z��*�a���{�F� �d�`̵��=#vǇ����H�J�j�B<Y�!exWRA+6.��£^�IM3 ���L-�R��|�KP�n0v��6"���J����#��X�]�8%v己���_���󗫟C!͙m�c�ޕ-�Dԧ��,T�s�	%�DF&�K�*�a����m���۷o���z2�׸O,v�J�x�\�+8���d���bI�9�%��ըA9Zh���o}�|�AE�*����5q[�(\��٧����K��K�Hf���S{-�W�F�~��+}BEƗ�<�'�`8s8I:#tY�m��W�dO蔌F&�j) �K��|��s�`���������E��dw6��'j��؀�����-�?S����g��ͣp��s�{�,P�	X6\�hE����$e�_\\��qrO`���Ү #� �+�L�� CpG���_����
ؽ:_�m��[4�>d�:.��Ӣ{�:P��7��{s�+�i���w������"�.��z*��ruf� ��g̞p�P���U)[fm��l3�_Rޭ&	q �]T<*.
�K꒸T�S�}�����`���&YQ����g�$0�hW��EmK��.Ս�Ɩ��`�X�����;�B�D;I˞���/��o�vݓ[�I[��@�|H������������nU��x��"[�vڱ��G��eq��4���T�Q��������x��Nc>��Z����Z]���}@qR�/,��2�O�VQ�3'>G�s������U����G<4�IϠ�F�V�Q���@9�O2�^�
����D,�ns~�u �=]����U�5��9̛M���v`��'�b4��N�["t�GI��\���F:��ZM��5�&�ӏ�Q�@q���2�!r��6�7�ڋA��魮mytu�s��~{�w"�̡�ǆ�;Z a�Ƕ�򧤦��_2`�gg���2Xn�`r�G��6��}eY]Ґ���Qy�ʈ⧈�~g)�T�w���A�-�a��Go�%�,V���!�`�9�;��j���o��_��d�'^���s{f��Vx>�[����ݘ��7/TǛ�{3?���tǘ<�^����*W��PD(�Qh�y��Nq�xɶ!:99�ϸ��Y�R�;��eP���FGcsv��A0VT���J˷vq�wDFl�+J��4�h��T�Ⱥy�4�mI��1�|����,�*Ҟ�)aS�>���n�;0k{�~y�r2X��c�F~O���]oS�-O�$Rla��J���S���[��U�a�>ϝ�.g��}y��T&C||g?�r��M1�^�?V����h�
�P�Ø7�\��� ������?R1�I�ӟm��OV�>��82 *%��w���Ƌ_��D�u$��ſK7,�J���"E{��S%^|�>.�k���:���܀��:"Ո��ޜ*��'��&�A����?�0�̓�]6�S;�ÌE���|�*{�#$��=��K+��U�5�m����LMM�K�V��z}�~E�i[�	�/�.�H���V��e�ȧ*��6F���?���^�T�,x�
�x��X��v�.�u4��hK&7�G�p(F��;<���U��XryR\\T����H
q7��'���������(�>
f����K�X�֙�F�&���{�����k��_��ۺ _jJ	yﰈJ��ZmubM���U��	Ứ�޷���!ׅ,��
T��_XM�7��B�-�Y�/�����&^߇�K�,]Li���pה8��xح�m�l�����7��L�K�^0T�����N��J���\S�å1������ݙHB�;�Y�C�R{��#��b��W��E�@ҭ͓#��*RB�撡M�7�9#h�Yz�}��`3Ë�͆^m����<���Ȇ�M��73Э���� ���?C3'_���%�,>T\�Fܚ����ը����s�](��Ls�ײ�HI���cT$'.��������]Gb��MrQ�Y���'�?\������d���]�g�c��P��	
XIgf��.WDk{ɒ��*��7)�9���ڱ�Ǎ{�&�b�̟}}d�U8�����F�S�{�r�(:�H���N��UNށ&�p���.�ĺ�.��珕D�B޽���b�G�$���G��_NEZ�[uj�:P�V}�*�OC4�V�/��X�~��{�׸��AV�3:#R���\�$w[�c�����Xh�Ȧ͚+K~���2"o�d�7�G�N�����
���P̑�����ҿ��,��~$P�f�<(��ź;+׎�1��1�5dd�-�%a�cL����ԛ�l�^�+l�N�Կ!-ґ��,
x2"���<DOk��P<=G�����]w��R�l�H���MP�Epտ^�w�o�D��~L^��-� ���(�
q8�ЩNF<p/c���7I=�w�g�TR��?M]zJ�@�ry����i.��ǏdLlҾ|yV>A�Q!�1�~�nfc4i'�.l�80C�+Lӵ�~5s'1��m�ΒHc9�R;���$9I��R�Qӥ�����|m�GkM-�����)0��Z{��}�����XCٜw�L�s�#��J�x�4�B��S���&8�����"�����]H��1��>�Y�=&s󲽳�s׃ʖ�c�P�5�w��ߍ���*���p��]��ȼ�6��F��Z<��e��@'[^�W-sX��IQ:�H�m�-�1�:\��hI6����ZS���yx\l4=�����AD����ň�J{�&9i��,C�T�N��Y���M�G��h;0�~�z����q�v��1m�,MV�h�0���n��. �J2}�i��J�~�Ƶ�mz�E���b��g�y������� �6�����D1P�@�?X��oگv��gs���c��j'�Xz�)��Lr��v��r���?r��	f�Hp�4��k1m�d��[��ݔ�%��g�q���>��w���,+-����66���J�5�m�~�f�#����w&�~�=�P���(K�YW�V��p��!���߁�����!�l�������,Y�zD?�p��Xg���.���5'��k��f��Go؁*�G�p��r��1�D��6���-v����˳����G�n�%�儖���	ut��,`ʼ;־6��=gX�@��!v�R*�,3^�7�?�_��S�w��
��6���F,���~Ӓ\5�c&5V� 2�<h�'�h����	�0��Z�p���heg�Hj']�G�u$����0W-!���km�1�V�C;�n��qN�?��K敀�?H��w;G{�/�\R�##L��yeIߖG#���,�X9�rP�NΕl�I��p���n�<G�He�E]��Vۯl���^��m��m��D�s7Mt�<�(���ݎBNG>R�y�\�R<�3ss5h^����>]:��9fu%�`J}��Y�j��ײ_�|�� <g
�`|���Ff2��H=�?���u}e��`R��E�6�{c����b�[6��^��2�=t\`H��v{U`�Gb����/[D�?��ٰ=���C���$�+r"g��|�s�Y�1b�c񎹄'Y���-G�TS�r��#�����5��>i[�����_�1Uw�Wγ���1V���.���O��Pk���:�wC��iB�o������nK�͍f�� �J'1qW�}�;Ki��		���6 D�V���,�EUi��B��W��Dg#?�gY�Q��b���|ǅ��I���R�w��� �ݎh�
‛��o6g����ԇ@1��r9�{���?�7��������4�K+h���ױ�k�܀ؔJֶ�{���Sa:����`��Z�����ԏ�}�I�f�;��M����C9��{������N(�T�yw�RoMc�n�^�߀L��`���꡽i�+��,�cvx��3�vD%��U�xs�y�o��OV���c����Q*l��_���M��K?������j�$����!���͞Gc���{y��y���Q~��9&!� �O�kV�Б䒏�M�`{)[�ȸ������˳`Y'J��9�q��B��;�GK��3}8�Ճ�Jf��ʕ@�ʊrpv:U��9x����Y�ٍ����l�~��
OQ��Տ@��@��u���{��-�Ey@�)\�$��~M%��'��'�2[ �����I�������r�ֽ��(�QR4p�c���۱�7j�������!�UUW�䰐V�)#U�{�b�� �������?VͰ��͋3>c߸��ܽ��$׷��;g3�zM��@���v�9�#���͚.}u�_Yc�9h|ܥB4F���~i�=� ��r�훓Hz��5��7�aC퓺���͜�U`�/'=��a�yQ�����/}`�v��f�uD���'�@�7+�U�
~�)8�GP�N[�X�����]��]滨e;\�/iQ
��������e�����څ3wŤ�.d���"�b�y��4Nkj/އ���m'�}���te�KZmm�-�v��{�7��T�T?�%YY�7�4��˦��zK�$޴�;V�Y�,;�_6���S�w֜�1w���"��]��ho�J_�����AIF��/�`�������}��\�Z%��|����3˿i<��q+y�dT^��7�_�ra���S�G����:�������x�v_���r�JMm����ˠ����[��n�gf��ۓ1���WS;����qq�9"��Y�:�M	V�I��s%�h'�<�Y�|%��1�3�
��0cWT\9g�B��EI�ʩ2��r�#�R����Ԫ�1"r�Q�JwG ӯ�X3�j�{�Ug�|c�7㍅ L�i.w~�Ȋ���.�K��P>n��߂Tt�'/�w��+-zc)0�zf������\��=I�:Aq�H���X��	%�� aE��F*�f����ٝ ����o|�7Pv�-���W�k�����o.�K�}�*�ҥ������J��饂,���A���8ertx��/�Z�������x*�QA����Qeg�b��A+[?�����9{��w����ǱG�3��4��⊿*k�q 'W�����ݪY$WH5��/^�@��$��<��Xɸ�,)bݬ���-m�||Yʎ]�#��Z)���3��x<��_y�ȑu4��ɐ/��<���\�G��Ÿ^j�.K�-�����É��p�"��r�6���~�ZZ���Y.,G��+�o��W����߁V�@o"����3\��)��&����Q[����@�Jܿom韲�R�V��*���`cK�hpV�Mܷ��aє	�D9hվ���]�5#h���[�g���cs�O��/�IkO ����X#.j�N�XLUAf⫏�Z��������U�/� �E.����1�/
ꅙeoJ�un��B���Z�lm���"�H1_�\��x����c�布��!+��a���9Q�љ@Ҧޔ
b�;\M���n��[NB/�ӻ	��?''�C��5qN��P��1�����%ʫ/�q+�}D�`������Y#H{O��N���6������HԸ�?޽Qʍ�L�(�'��o�ʦ!ګ<��G����k�3���$��Ժˡ�P�ֵgD��d�6�I��+f[֎J�H��0}�D���Dɟ�2�/K�tz'vR���������e�tk��ɘ{,�;a�}jXA$��z+Z �c���g���"�*��}.�@CakDfA93*��U�
�R��۵j��:��.U���c�U>�?
R�5tÞ\�%/�t�E��T���,�D��Ǻ����K=w
�|��\�Φ�:렋��m�˧Eu�❳�<����Ψ(�l�O"Y�M%�{������<�����S�}@�YH^�`��U��V��jZA�'j�/�����/��Lŀ�L-Je� >s*�fIZ�vQ[J	�zc�}��v�ƉwF}�$]=�h%�D�ז{2��#ZQH�Y���P"��	�,���_Ro�s.���G��S�ܮM����+�A=��3�8�9��ʸ�3c������yw\C2w��v�ڡ"��s�Q3�=~�h>鷷��?COೈ����>ssR@f���早(/�O�[�ҽ��4��l7��jT��5P{��	��կ=��6�l���Gt>�D�W=r9�*D�[kV%���{���,{5�OK!�*�[����&*�S��Zrׂ�2�1��Ax�t�x'����^�j��^�������󻦶6&�9�_NN^O��>.��Ǚb!�[=�%o�ZY������Y�j��=Y	�1�nT,��#��BL(�XvfM~I�8��ѕ������Q���dIu�m�Y��J�{�pYJN�>�c�׸s�r�ɭ]~���(��eUS��d	[��`��gdΦ�6��Ѧ�pi�9�T�P�i/sŵ�+m�W-C@��|��.�Ip	ZZ�\�Ѿ3�g������N�k�dgR�ΏH��(�vv�f"��G�[	���<�@�D,�����ji^�u��sW~�A=��L�w�+c�o1v9$���2q s�U��5�JT��p�&+��,�~����_^�9�߰zR9=�*��so>՝�XG�O`UbC\�凅���԰<�&�V�}r~�ȈB�n_����۵�w]L`���V�C����A�lYv�+�~>SX�������:�GP,�(7D�gvNY@b?j������5�~xؑ�8y�UcV��OP�3��ڼb��<��� �G�ċ��N��+�z�MH9j%�§D��&��o��Ɔ���rdWޟH��0�6o0t���ֱ�.1�U��x�~�qW�xbXC�ȭ�M��ӝ��0�KS��(��+���b��R&�Dv cC�:üKYI�J�4�Ɔ�G�^.�;7_�!_[%ά!]s��͘a����p�Ӄ����*�xX����LgͭR\#��q]d��4�EL�엛���8�9e�u���!�_m7g��y]��TX�iT���z#Jc�ڐ�J|��0��ab�=��鿸�id�G��g�{�Ɉ�����6�|45Xa�1��_����E�Z\T�~��c�����l��0#;˛�{�r�?��
��1|uԭ�����],�n;A�d��s)�(mz��Z��ݮ�H&����4;<[>M�Ǜ5�a1tWZʫX�0FI��;�7�a����X�澢K�����6��Y�<vRy��-����c8oxDi��d��r��	ԩ3���Q]�����_��pۖ��y󨰷\�^]D�Y�ړRK��k������<I�}�l���c��O����2n�YRǋ��!w�}�S�$W��])錹�~$������fds�eY�`3ʯ��P6^�`3=��Tv���-0��/��Ot��$�����C�2A�n̎�e�fc�2�O��[�z��ü�&�}��������e�l"jZ�����|�7�W���vϜ�ݶ����O��y@��Z֤�j�a�ҭ�4���}�BӞ!.�^́�c$�-u1rm�L��a�-��M2Tl����D����Ά�PK�Y|��`��}��s}�4Q�)�n���X��4JR�{��,ˁkX�F�MV���OB����1�]fcq�̰݇)���8s�ą�B4�u*��	�9�Ѳ
v3��ND)~a��B�m��̔�b��J�,��ϕ�rxHa��/j-_�����f�=d�-�O�QPz�E1��v�;�S[լٵn�iVl.���\騔!7P]�5�M&D��@.����i���|Ա}���z?�[����>�h�Wy`�a�W o��F�퍒۹������G"���{ȹ4g&��m�x�3�`��,1Rv�xb\�{^�
�q�|���6��F? ؈x�q���^���B>�=�b�l�`���v`�
�h��kaI�g��^��ܬ[b�)���!Ƿ����V�y�O���4�e���t`z_���,v6��0����E�S��Lߟ*�����D^��0��~��v�����x�:�Ju�|�VꅄЈCs����q�Sύ�%X�c�O+�汛ě�JH�1}��b=�����֌e%������{��q�״���]x�s/N썳��m���k��`�l}�ŝ,fM�\�>�vQ��u��8���7;�u��/?t��]K� ԝل��=C_�i�)���bC��_2qY$�5(��Xi��u_ ����J��d���k�8����PE92#C�G[���zV�C��ؤ�	�*�|�Ҡ�!�/�;�f�NÓ����֗��]���Mؙ��^e��2�����Z����x���!�|�`���Y����9�4{�SkH�l��۵6��*;5\A��(U5[i�k#�pL�_�/��kS����'�y��t�pOw��һ�

I��A�<w�����QU60u�!��^�z����f��d.Q�4�C��/9�flwj���(�I�ԾvXJ��2� @b=-���z�Dy���럭#��P���Y�M��ѕ֗?��>1}o�S�T��M[��"A����o�*|-0��i��&�,���Ա�Z]����;0ǂ<���^��QN]K3;uK����9�-�W�b��ʶ��StS��^����3�Y7^(���z�6 )4�TB����|l�J�K�z�5�M�_�{;���]��b�uL/g�}��6^�����gb�����ōk��u�Ɗ&�ū��pM��	5��ߛ^Yì�`;��[;��"���>���o�
;�:�,�����'�b��Iӥ{���i��Q���Y��0��h�p�l��u��Cy 	��+-e�} 	����mr�=>���|������,>���}9t�w�s$�����gN�zC��B�	R9�C�.d�|�c����������_�z#=�tΪ9�{��f@�To{�T��]�Ũ��H�n�ʕ�X�w�fOД��Vj���@�����BP>o>h!N�*�MC��_�j]З!��n� 7�Jx���F��~�j?+��	�g�X�۷�Ba;W�^ìo���5������%�k�y�(gBxKx�v9������Es������e�խ����'���_��ЈՑ�����YnLZ�!a��)�p�g�/���e��.\Iޗ�������G����Hf��S�J)���	 S�VT�O˂�zD�A��%�w�R��DQ�k��g����韞���;���]3�:Z�a�G��}�Έ|���͋��-d��J 3f6�1}�]we��_��m��C;to�.�@�U8泅�xSL�(źF�*��R�*��Ae=Ř?��\Sϧ����2%!L���e��8�����M���(A�k���1憬�eXhl2;��?y/y�m_���T���V��?�:|�58�
C�U�e��bgxe���}�8����NlPX�J��T��b#�m���-q>�0��#�ߑ��m�7�U���*���ao��o����!"sxkUJ�D��q���&�/�P�da���=�e���I�~�l�� ����J7]ȟ�C���Gۈ5pX�[�y}^��l�B/X?"�	��U��X�����UTW�d^�f���K�O[�7ʶ���u@A�vr��j�j4 7nJ����qUy�vn]�p����T�ˏP^�o�':O?G���TgͼyK�L�8%!��r��vV��'����o$�	��d�Z��h�S���I�G�0�~��PV���ٻT]z>4�j�������s��h�>%a��8�n)�lIt�(��7 ;�]��D�5�H�_q79�٭!\A˽���Gq:�l-vHQ�)�庲W~���%{��9��#���F��� (�ޛZUy�r(�@���(L2����)=��3^6"9��bi'���^���w��H34R-z��WY��2⺁�Y��]^eN4�Y������:�ds�-��W��q'�9�CuK(�o�����@���T�/�d�v����"=���ض!-z|�1~]���c(ݪ=��Jj"uF]p�T�Q�@�@��O��.P�gU~�%�N�Z?�ٗ=g����mF��,��]�Q������Ҵ�T�m��k��X>�ل�Ug�"R����i���#�o��|�<������Q['�;x�~ `�7����S���ƧT�s�aT�Nێ��=cU�;*�J�R��5��Bfq��@�X���%�K�� /�4wև�&Ԫ�WŴW�W��Y¤R����5������R�{�ٗ��N�|�e��r�Ά�߬��=�� E�?~C+�� �Z�Qh��$ek9��KBwx3YRwN�	&utm�!W�_�[��s�V�<e���S�}��5l�_)S,��ԩx ��
��Ok6����]�]~�D�|.�U��A]4z�����u����[�h|W����^�,�ԡ;��#0bD�#�i_5C��2�����]���6z�ypQ7���{̆�po�%�9�j��&�n�N�X?�'��e����x���Y��z_��`���z�WV!���yp����z��ox���%��۸Ise����s��(��tF�U�%3�ی��[���D\͘��B���A��00�Ռ��G^Ț��L�����O�d�fW�Y�ٲt����9'ã��I�`�[���r�����$��>G����T-����̩���P��)���נ
H��:�/��76���:W���8��U�n3s���HC����[�Ag���7�z���4xKԈ&���Uqz��� 䢏��U�>Tw�Қ��}D��&7�������z�����ג�s0��H>���&d��Iz�Ay�r۷�p|7���o:�2t��B�!��i��!�d���ϱ�T�ɗ�;�M����n�v�!O���9]�;��w|�����[}�CzF�S�x�b�m�?�� �t?id�3�pF�mz^�3����R�L%�:%@
c��H�9�O�O���Movff�5TL�:��p
�+�Jo��?��^Z����L�m;wn؉E�jI��<�!C}PI}��^)�෈���Ug+��LrK)|�֨��am����;���מ�='d% 4��*�ѼQZ:��b�SHY~+i3̋���+S��)Qm�����	Yc!�C��.�UV��C�t���B�d%'���DU�JS�m��k�V�_��>G�.[�z(V���m��	w��g��Hc����Ⱦ9���پ���֭���P�
�q+}^N�����9Oi�����w[�?����qFꮞ���j�aM��%vgT��]܂ǏzGx�'/[�:`��DO�(e�������v��d�"�~g�m,#A�K7lx�-�����S��S:Jۿ�nӓ�Ϩp����ޥ�ݳ�F����鼐���P�pݣ����[�����{��W�c�GR�l�E��a�=�iUlU<���o���B���mE��ىn�*�@2;`u�/<��9�����y�E�u�V���Y^���E��A�2$���?�?�<���J��z���'�^�B/�����i�xK//��J��h����H���"1��~�*+s�=�^��ʖ/G}M��M���wa�3u��J.���^���2^�2��IBv`yx|_��Om��D���3��>#�j:�7�I��_"ܛ���*�ɸ�v :���`�L]C#N/f�[_��L������fPD(��'����T�5��4Q��F8�
Ȅ���'��`K��+���W�g�P��[<�e�=.F�g-�v.�/�F^�=.̄�lz�p�+Y^R��*�x��]�����cAtC���`t�j����FP���^Q5\D�h�c��&q���b�^n}כ��;GQ��3Y�
�"��F��qN�BQ;�Hp�
b��7�9�����E�)��p�eFD�~��3�a0֓�[Q��L1���/���_�4�G(Ǯ$�ds#X؀#�	�d����N�b�����lL�V};��X��Ӝͪ5a�:�qx�������2O� �ɸ#��Rقq���I�OSI�u/�֨�J�`e���Z������`M��/M?#t�#�����;�Ch��c�
��;3���e���L�2���ć�7�|��o�_�*t��:�����{e$T29P�)!u����ݤ!aΑ}���욢Ѫ�%`<�����}��E���RN<ϹC���_J\I�-T��f�����Y�w&�R&�� �r:���?��'Y���ނ_�6Q��-Bn���.%Ltaٖ���0�G��R%�%V�31P�C��'�<�U9�T3X"����s��J�����Y�h>��I��Y"CI&���0|y�����41�맸һ]�YV�ʍ��Lg�V?�j� �֖8^�X"��F�:.fĶ�7�|��n-xy�_�O\�4Ol��y����E���ml�@5;�ڨ��K��	C5e`vЅo���M��^'߱�e��WÇu�ڭ��m�+?S�Mw�żՌ4JHH02�c�[I7�e?�S�35޻y�I�s8T�~%����Z9]���{�+��d@W��@�z��(��{��f�ĘN��\ �u�T����}@�]��ߺ(�u�W ���t-�����L|i{'eG������.t���4�R���Jm�e�I��Wh��M��L�ѿٍ�� !��Q��@.ͱK�V�Ҫ(P�60 �����~�2G z����O��x{����=g�C���'ŵ��fG]�BUv>g��B�=I�_wT2B�?�ѐNJ��6��	�1��������	)^�����}�P_^�j#I@ćmֵ �vI
Ⱦrvjʛ.R~���H�i�D�3�*�3����Q��ѹYa��G�������	��~x�Ñ^����"&�,���ČFRv�	����X���c�7!�:�9�m�	u��(�s��p1�����FJ3����w��uH���ܖyl���g���ו�[+B#(7�A�{�K�Yo�f5HB�H�����Q�q�#���U��-FY�k܊�}[���e��hgcY�8��b��Tt.�4��v��\mw����Ӎ��Yd}��k,�:7=UC "�-b${F�g�����7�.Ր�4�&1JUI��>%�=\�_{sX�E_G���[ivn΂���@���Ȩ����G�4��1&�{�3��H�m�
"�c=��]/DN�^1a9��7��Ѥs�	�"�JD�=��ow��^��V� �k��3*Ta�_�9ys�d�h����_���ВW��	���_8NIM���Ap���F��1B��&\D�����}�\���D����WѢ�GGݱ��J�n���	�w{�DA����S�� 揋P^�]�vu96ne��-.��et{�8gl����lMa6Gi=���D����7�'�2H�M(��N�_��h�O�1Ѕa	��)�Y!���mбdR�q��՛{�3e��jdA$Qs��b�d��>���*<�����ۮgV!U�oI�+r���'�A�
�'�x+��l��'�[n�Y[�+��z^�5��o*Wl�PJ]�m�����x�G`�O�%���k���n��Q;f��%v�����7��:,%�I�d�VhkR�qN\F��[�_y�z�0k�p���\�]�*�.���~�yƾQ ��ֶ��������X��
�����V5Jb��l7>S	�����=�SZa����@����ي���9��n�e+$�}�F�3�*B�_��<&s�͘�V*��v�����y��Z��u��e�(u�&~E�m�QR����/�$��~�$�L_R��	Dg4�k�Ng�`Eg��&�� M���91O)�6�;��6{W7��ߙI}�q������P��kc�ф;Gv'��̔����)>?�Ur�{>zf76b&x�xA4��Nk]��#6�u���~���a�m�){u˥�T����H�����f����'?{p�wC�B��c��� XI>�~v�Y�1 L>����0��|�חV3�S��B�"�,o�����(&�H��壖�it>��j<x�)�~~�Cr2���c|s�� o��H�C�K����Ry��\�2��J�
'i<�s6=����(�8�B5m��kd�T8S�c����y��u�)�$�Rʈ��L��M�r�w��{�S`5�+�j�؞��8�_z9�ѣ;���Y��`~��C��
M�כ����=��I��3^:j�#��܏4���g�@�*y�7�syOMx�e����3���t�9Ň��e(\�?��8B):oH�u�Ӄ^)b�׾>v�BJn�}�$ʅ0�U�0VIxWl�.FrJ��H���lS!+.�H/��L��c��r��o^6|�-/ȯ������*c��^,�\ZS���E$�犞CU�t�W��͆���>���暍���������4�z�MU���_/[��r�6)�n{�o�n��3z`:�#p$3.(p�%9�Z[w�V&dY�QhS~�a0�o�
@�t��Cz?��/~��o��Ah����l�S�sA�Ò����>)��^�-�<��ֈa�s��x��Qf�&�@�"<'u�%���n����#g�@|�S�&���_�3tO��Z>��Ӄ4]ZՋ�j�%��a����ߊ�8��鋀�MM?"���g��ŉ�h�W)No��Y((�X��������j��7�� �Y�s_{4�f�!N�^�/�Kq��[{\H1ڃk!�X�+aB!��N��:�l�<{��̑iPA[�0����@lX��ו~v��rE�/	��i~����1B����_k�lރu��gDx������6!�A��}�r��,.�~2:�f�E��U��5��H�T�a[���bW̅���C��t��R2��	g���J�G� ���xf$4h��픗�9�3���"LEkBl��Zf<������Ͼř<w��=� �#Ц�;�]�]�`Y���{i6���L���;�n��u�a�����	�a�S4�`�
�f�i��O���E�B�� -�a���s�cdc�<p�7vO$�{H�{.߳���v��J�t�p��S�^��ٜ%�l��ÔJ&�V�Ƹ<�C�h}���V	�N_�U�u���t`7����ˮ"���V��s}�R�����Q���ro�{�$K�m��{���4�ϩA���N�-��0tṸ�o^��Q��O+���6F�����`��z(���7�,����?ߣʃ��Z�ccI99;�� �骏�\]m��6-A�a� VG���W��Q�� ��/�o�᷼�ІTP�JW����J�(s�zJ9���P|�����"�ȓ����	�L��[K�2�oM��%��xS~�[�S�b�Qj&yy��K\xOn�i�{q��V��Y�	��G���>�B���+�GZi����ZwJ��{^R��d�͇���4�F��o��]��zV��dgߌ�����,;%�/l�i.�9��G,�s(K���ͽ*�a��p���a�r&)�����P���}�ptź���7�k��3�ؐ�M����o��he�,�\�給�y #k�x�JnZ���`�&��P�c�'le�����Xz�)4�f�ݼ���6����}��Զ�c'�aDѪ7"�(�	O���dEqڤ�xt�{���Z�}�0X;�K�Ng��GD�)B&0�)���I&�}:���J�ǳg��߁_�������+��'N��7�+)3b��^�GXSow�����z�:5/��?r�|G�?|}��-���~Uo~%�<��SdIUC�{P����AsO�ܵ�P���tr���<<'c�u��7����?���ﴹ��a�)�9�s����^?�r�L��>l�oߟG�:wRi��[w*�C��[�
���l�9��Qʟ���͟	��
@4���Q���z�^G�_C�wkS��Y�.�L�sK�ɿ�i�}���(�@�vupC�䆄8��ѷ�P8���~�^x���H�����	{�T��{��B]��!����u���!�Vh1��� �������'u��`(9������)���>���g]��%V���G��i(��� ��b�f~���$�����K_���ב��*���@�H(g���E����T6ml��BM -P·�9�(^��j�^���hN�2ҧ�����>Ǔ�D!#a�UYy�"�J�b���@KJy�Y�h!��k8Y1�y���J&�)��M�[h4
�{U��5���:j����D�����������" v�9ǯ|���oEz�HMOFK}玳���K3�us�nq'Cq6��1HH��N�	�=܎pY�mI���<�?}�]g���8��Yr�iؠ}��7d�������e���H	a�o�*]�J�	ˆ���8^���I������G>,Y�~����ﳹ&Gb��0�!T��@�@#-9:��~�Vw������/?���� #/[e�˄O�W<���R8[���nb����ǀp`�D�'W"�r�kq��>�lR�l��ѽz3?M�Z��ǖ��Yv����%��{ʦG��xm���Z|3Iw벋��6�;�;��n%�շ��6��ҥM��٪�M���h䆅`G�W
W��?��;�7��ޫj������tش�7���j�V	J��Z{��W��"f�;b�������/�9�s����{��}-BqWq�@t��s�#ё��Tl�>w'[�k�uW��$i��a��~��/�T�H�:���i�E/��?xĲ��9P��<q_ۮ9X9k ���ڢ����n8����[h_`���u��x���4�r�%Cw�rh�+�k�0��,��U �&�m��S���J��x�I�h���z��!����%R�Bw.p��}����s�)�Q oAy�� ���4�����*Fpi�a��d�}�Q�A�&��~��K��fԀ��u�ύJ�uؚV=X����ո^̼��F����%�H� ������j�C_���_x���PzF��7i�V���
U�1*��m4�hx�]2��<ь��I(�t1x��#[���2id�� ��]�o��ɮ��������A�n��#�Y���<��!(;b�oT��EU�|�y���H`����'vo��qNK��MȪ�Uu@��}j�u.A�,E[ߟ��s�oI���W�~��Ә�QZ���x�7��+M<>��@�Y��uZs����f֔jhy�����g2��ݾ���__��j'�G){0I������c`���#&��$J26���,=�Q7]�p�s��v b���>d�CA^�>���1^�r��ڞKs!�Z?M�������b�?v��5�9�7�5�
D��V|@l�ĈV�,��s0\��1x;}�~B!e#d�U���;���-Rnu��� ��,
�ˉ"5��Wn!q�.��`[�`���\x�����M��V���W|�����ٌ�(f�J#R��mE��,�H�l,�-j�\�R��C[��b��m��h?����7��.s�	�~p�o����Y��H�]+�	�<�c(�C�sW����pys��6@���U�Mn;��IM8f�e"W��|(�x�~t${�_�Ҏ2��*����.P�('��FT0zilo��d���\uC���
��;��Υ��4�4F��k��s�z����}~~ʅ�.CWϾӨ Rz7j7�(�j�!4`�両��VCG9͙�|�����3:7h����	Y\��t^����ja�7�H��?��^��9~��(�C���n���7R^�KFT�'ɦ�ʢV-�t�V����6��?Qc q>�ڜ�_�\J&,!��[^���X�u���b��A��a���(.s��GJ�M�k���Bf�G��z[��d*�F�`�����?] a��21r��Z��v�ƣ�A�9�JB�/ȑYk�4�]_B���?o?�m�|�*Qu�c��hM��#���4.��Nx�M�=�1j��G�d�iC>Nň}��w� ����ϻ3�ˆU�����>J��؝9}�����X9Ҽ���k�����r�~�����w@�+7�'������~�j0}�6��Ѣ姀1��������A�K��V�o�]`�n�.]���>sR#̨�48�^����3=~ŇZ�l�ȉFC��������-f�7���1��uE�+!f��=� �]��Ta ����~K�Z����r���?��X��W W�u'x��r%�&i�4k+Y'i{�Zo�(��Gm濪���ϭp���s�����@>��8=�P��w�]/.�������A��d���N�d\%�.!���d�8�;�cq��J],2��	�9t���
���.��[<
)~+{Y���#��-��J%}��g�������ʦޒU�C݈��V�x/	�,�t��n$��VΖb�C"^��T5W��5��Ԕ\u��aunr�umAǣ6X��b"V�����5.]�7���|ޱ������۟`��9AU�������G�D7$r���d)�\���I_��N��»�Q��p��d�@�	�lI��b��k/����w!��Ŏ:cά?�w�;an��ʐ�&@fc��@*��("M=dNz"�V�h.�������Q�ԕ"��C���dE&l�Ȫmӆ+�Np~�5�x'��X��'�_0��X-��ܯ��0���.ӻ��n�g�A������	����r�\��D��~��^����O,Y���3���Ӫs;I�0�Rk����h�t�0YTh��I�%I���h��5� A���U*���?�7t����@�j8��c	���U�w��E��t�
��S�Y)@|�3���	s>ɞD�`��c��>~��zY���=ោ��^ܸ��P��\k�� �������dW�������w½00�兢���.tܝf3欓�b_v*dhS��u��理O�Ф��3�1�g��~�iRE?���;��{j2�M49"�7֎cP�0���ϖ�"bde��.��B����?o��gA�i�)�h�z�/㾦*�o�µh��P�k��dJ���Dm�N���t�4&�N����'�}nr���Oq���UO���oc�����:���!�3|t`8���ډ�ꂏ��D׵Z0qS�,�<[���͓y��I��+�a�����I���h���r��8'��f�� 	�����ū�Q�X?`W�,�&6���Q=�Y���/֤� M6v��:@�8�qRv��Yq���m�<cۢ�Įr�b��)Lq�Y�Ԥ�����qx��hjյ�6R����}@7.�1^4���z��z��A��-�E.��1���m�8��%*���oރ����9P@����ω�{��;0�Y�;�c8��&\�U 	�d k���z��G���|�n�>��8.{�O��S���S6��'\w�e���"��37������~~��]�հ�B�2�0�Z��?ū��sx ��<�-����K�/�=U]WY���i+MV�-����h%9[Y�ż���i�$��#<5�I�6����&|�4����(�J�m�o`�'_�2]^0��1q�;�����B�U��\�3��>��$����H��x�]�&����x6F1����8Ϳ�&�9S�е����rz�2v?�
 �l�����2L�[GH��?�3�Ӄ+�qȷ5K�(�{�~,'2YݯPP7���)�xf~�M������0�\��)�����,!��68ԍ5���r)Y�����Üc5�5�J
ޜ�*M��z��{ߗ���ᾔ�F�c:o�J}@œ$`��vwux+�!M�����=��<���Ss�"�����f��%��TX��R� C�o�8���p�mNO�[*tbn����Bc8zt;>⏨�s�\�+dk}A�Ls��=m�`�k�L�������VDX�5��̓~K4W��ZIM7�M�7p�i��o-ſ�����������ځ��ۡs��ς�*�'N�)&�gy T�����E`oM�D�'����Tt�΄[�F?1?#2�C�	��W[?���?�1���̜8G �����(�G͠� ���0!-+�1��>�ȋ�b���r)��b�⸚>���U5'����u)��Z]j�Up��$ʦ�]��P��8Z�kg���Yȱ���l�JP��v��a��|���}툶2+� O C�6��f��]=8=}�8�M��p���ZC���0Ml�#hB]���H���$�?�t��-���˒�P�ںxe����$�����1(��n��(��n�3�����q �׈�X����0�-G�J#�PV$���e/)�s�.	܆�"8OSG�Ͼ�쎃�U��L�m�F���J&=C�6�o�w����ĵTZ�ZȤ2	4���
u[���څ�35^�/���ϸG��f�f��qoڈ��8d���1x���&>]�2r��r[�+�����t�L �j�l鬵�w\_5�V)O���5��_��L�R󖜔!Bt�����80��)��q����[�l;�G;�JX=����
���t��_7���)ҵ�����^���h��EИ������d�XA0�hƁ���m����$:n�3p��L���Ŀ����?����6lR(op��^ �|���K��?��V@� �:�Y�b����6)\@��`ڛ�r|��Ѕ��Q�j�wa��Y]P[�_�qg�ޙ�$�FK�Z<r��3����&Dw{�نwt�	/p<�0�"Ҽ�� �F�1�q&o��!_����zF7�g�~i��D�xI���Rn�0M�b���.�*PHд���3�ɴ����QυK۵�mi;9�F�@���Zu�r%�pFi�1Qp�b�jkU�ĸڅ�6>�*�����#�\��o��Z �����l H|T�w�`����"o��M�#���o����?Se�M<�����+����%�����l���f
).�d�~ً��5�RW%��|�x�N��E;�E���w�t�uQ�[�Y�j��e�������.�#|�X��=N�%�)m<R�ǉ/ȿF<g+H�=��pm��%f8'䐞���k��&�/��3:��ʀ���OS�`���d�W�6��߮/l���qd��8���ؾ��l�üڀ�Y@���v@L4�Bk �Xn�u�����]���g$:�N�M�/d��L&�Vng���Z�SP"������L	��P�K4*H*|�zz�Ҳ�ll�4v�0d0����1�
z�����9�g>0��OY����%�Cм�>�������X��/uC����|ݽ}=�O� 9��9�C���kn�ef�د ND�6�=�yے�It��!�{/�щ��q���lK��� ���uw&��/"�M�- ���,���hh�/����6��l��:r��c�)�^Ȣ������`ZۑY���~��R��Z/�'SDǄ���i�!`��K{�M���������.�Me��f��6���d�x�	2�O��
�v��f�+z�w��&̰T�Bd���1Ю�1S�o[l.8�����]�A����7�>�~���ۜ�}yt�:vu�1�|��Ja�o��\�w/��[ƣ�����%�p�Ԩt����\~h�`�R�F~�I�;e�٦�x���Ŵ(K�����B�;n�@���f��h�d��?�c�r�z�����Y�Pa��,��/�*��i�Z(����)������mXN�U���|��E�si��苶qv�#��o�>tȯ�4�8'�����~~ɡתL���r�8��˦)돵�놜p��\/�ADU�����9<nr�`��������O�'b�b ��>CG�ңL��O�j����)�/����������
�w�bs���d��&����x��:����[}�@���O��޴	SC"�3�N�2s�@��D��ķs��h��4���L��I�τ�MC6�c_q�I�➮�n"l_z�r��"��u��I�:�k3�Z�>�9��	���������D*	 z���h�R��dPGv�`�|I�j,��`�&�cԣ�	y�ng�Үiه�(��gŦ����.�D/��ߠ4T����W$_tlD�=!�c�V�cQ0!>d�Ob�͜G�Y�Y�U|��!P\��Q~�b��Y��8�D��[*l��[�,����VRW�����0,����X�1�×;C�"l�ۦ�
�ɢ��-s��Ǧ���X�@�5)�z�S�pz��E����^V=�̶�q�:,#e�X�����D�Q�'��KwO�Qj�_g�l������)�������n���Z�)�9ɓ�d���#�149b�!��m�̨����L��Lo*����E	&��GL��� ��p��$�9�r�b��dY��JV$����zJ�/��3=q72H�І���y�vZ}�	.EEЕ4�f�M�$*Qx[�C��vD���`{��}7�]���vsw��l"��0����=x�Z�hm��`�45��*��翭Y�t�`JbbbϿV���IW��#�Pml��ϻ���^�\�����g6�x��[��b��7�9�7A}��!n;=�R"wr��e�s�#���o����p��8��Mzd�r2:'8<����S�jTB>���X��ch�4��4r���zx�k�1�9��:7�zj\x�2Lrf��Ӥ��]�X�WwC��<
��	�������)J�L������!L�)�x�1SVzWqZ����3��c��jc$�/� 5�F4[a
5���H�� �{~��7��w�.6\a���4&��,7g�j���դ9;�UC
�:����m-���W5/D|ۆL�� �nm����G����01��|ͭ�Q�sF���E�s?(�ԃ���s�2TC��j�хf�h�������%6d���Ml��+w����$�t�Nd��E)ک�nX˚��o'��>�(�l>!��)Q�^	ڰ�u�X�*�1Z�*�;�S�2��di��5�>��:�M� �)
��O��|c	tflO�o��t��Z�~X�Y��[d���l�^=����`���6PѺBB�#%g�j�@k
o��W�^�i�ߴm~y_f�D����޳oېx�T�!��yf<w�6�.U)�U��"+�-pA�ƿI��
���G[CwS9��<��t#(�x�
ʻ�A�У�k��w �˥��e6�U5��%Y��d���rR��k����+0�����I�Ω=h3R��;9B��P��l�l���`�j�ܦ��#_%�0c�	�IRc<4�N�u��vN�9g�}�
�AڵJ�Jwj`�]n|\�2�Y�t��sҩ�^�v`E8���]�J£��O%�=޾��<m�z�$�Y.�X�6��-Q�����h'`�u[���y�V�=2��F�_d&2�Eq�M?V����؝A����4�V�MAo�u"�XI��/;�= [0���O��VF�44�Y%h-�o���騟�ꐰ���3���
��7�h���s�m���)��Yվ�P4NV����h���{2��`�]4 8g��b{�/YI޳B+�v`���^��}���O�_�遨`4�H��%7�ez����V�ďm �w���<�4H�������c�2��t�?��6��G���c���������7���;��F1�<���@���y��.��Y����,#[�*�4�����-�H��9F���� >�tk���-2���hvu�/�w�|������\,�3��Cҷl�c<S��bjDh�>(�q����.�����x�Q.Ǆl�aY��zf���X��Pj���P���1�υ���n�:ì��L�@ClPj�������T���4�Ǫ����2M5�go�x�FP�P�� ;��L�OHN�O�H�o�Wk���f�ƭ��*�Lf�Zw��ON2�uw	�N_��B�N��~�:!�M�uC�����lZ��T^���f�w[p��U��$���f�~D3o���+K�Z]�;;�BV}_{Z�j%ˌ�#I�`gn$��"?�l7�����?�L���)Z��Vg��k�)�F��ܤgӊ�黱�)vؘ���R�Ҝ����e��Ù ��]��?�ȍ�qm�m����-��W2�7#��ѡ���r���s�l%Ri7�K�#��� ^�^���ޡ;�Qe_=���V�VǗE݉Ag�d��ɸ��
Y�"�[�{1Vʵ9jj�)�?쟴��gO��H?U%]�3�E$�$@���Rk՜�.)�t������-Yr��<��K���oq*�GԺ�+�'�'�c#����XV�h��|���r���+��p�>�߹"lz���~'g�.c��.�b����F����֠���%/��ʊ~eA��zU���*��q������E��ܵ/sf�'�Gs���_j��9w�I�����sKv�K;/{�zniz�?W�����5{�ܭ����o��2�h^Iq6�1�I����K�ȂE&kV���_`�\��}0���ܾZsri��@�����
4�坧uq{v8^�L%z�(#���_��uJW��0��>W���q������0����k)�N{����)H9��]�t
�T6?s]��Y���*[
�e�A��n����Z9x��!��Hc�ճ�g��B�v=�Fe��JC ���_��jl�,z��e܌��%C��{�Q�&�(�߷���(͸=๿�L�w�� U�p�݉�1뷟��u��@��n�������`�>����{�j>/�һ.k3������"3�Y�U���q�B?�}�Ψdz�`'qU�e��fZ�%�9`M�	����9sS �6��() �pI�G4��[�f��.�Iߦ@Q�ԡmy�^�L�IJu��(���E&LV�`A)�O�V�2�_*��O���.�	4J���!K>�Z�3�Ճ u cm�,؎��C����;#��݆���L��ȢN���-��b�j�_f��%�1�Yp�H��H��mc7�nd8ES�v��[�nK��t^,�"Z����0�Y`�f{�Nq�
w�Føb�o+_=��/UW7/y}S��f���-D��s�O�	�t#/t~��`;�&�D��H���G��F��-��a������n_�u��np-z|D�T�3'��\�OPY{l�n<KC���Jw\������2�Sm�7��󵛪Ilԟw��\R�Zm��wkH�d��d�R��5��[a��*~V�[�c�3�1x]Z��U�c"AU�i�M*%��5M	=�#�D� �ˈ�GNi����i�_�	�S�B0��.F�墘�*���路Yȣҫ�N�u�N�����X
�?�R��Ճk�����͂��Cy�'@_����&?{&���(N#���zo����M�0���8c��=n�Lf�|baN+��b��JU$a	$��gz�C0�i!UB�K���4[��B��r�U"�:��?T�����B�]|b`����=��F%�U�+UN�N�/Ta����<��I��q�a�/��p���"���������½
�[g�+�?6��yj��-L�Q��K�0�3�:��"oa2�Ճ6����w�5�˻FiM�P�f3���������xs�u�c����k�B��yE���t��ۭ���/��o_h�YM3q����ޡ.�W-��L�	~˲&�������{(͕f#����T�$D\�Z]�ɻ�-Y"�5&��h4��	��Λ��#2�v*�K�(,OC���:�@����]O��q�z;B4�b�3���䳭�lSD�ҋ�ǚΫ�l8�P�S���_M��5���i�:���<RB�VM$�Nb���P^���!�V�B�'`�d�+`]�_�6/ۉ�F��]'�q�*I`\�L�Ӌ~��n(|0-����~��O|K���دCb]��5;S����.�����T��}���=��k⌟�&
t��he�kJ$e��d�5���[ә~g~ ���)cc��������񵗥�6���زO<�T���g�='�]�@����
��מ	��-k9'�fh���F�uT�a�/#�. ���Vݧ���/e�{��(>|����	�vZ(�����9��X-^�i=U��i��~U�`������W�|[�=y�ڲ�A$GS�b��MpV5~7K�T�&A_��V "v��[�m7̭e����C�����ԥB3�i�c81��uժ�`�
�!"��ͮ%k��[��,�fR�)oJ٘�_�����v�qd��=�.Rz}	�rU�*]L��,��'P�>K�M������Y��7�'_�&{��X�"+<��O:y���ß����&���Oj�<�k�s`xz-1���#'	S��~�J>�<kT�o{��3wnV�|�#��C����?V-p��ޅ��N8�����1��D&�}�ʈ,�{�h퉏n�7�0��� �� �Q0���Hc���v�V��	�7�^���0z�JwF{(�:���iOi1��K��+S"v���Fܠ��<A��~Չ���	�)�UL��5[���:�M�r���<?vvrrBU�$���_����Fe<���V�0��3T$��<��#%&�!����P\8-��{��7A�X���%�%�!o`��5�6`�}����j��ѧ��?������V��k%XY�^2�̈́�/6�f�u��~��/��IəZd\|��B��>z_�^�(({y2�4�)���赀�^�-O4�� |A���sb�ڡm6����nZ�����a�w�6���F��,��?�(�FW �� H�sW�D+���@M��ք��O�=��@�$%j���~��0L�������oM�A^S����`{�����p�C�a8S�E�jH��B���Oh���Bf)ڲ�v�7�Iq�ឍ�]t��g�f���1k�5(���kr�����h��ճ�sQR�-�"$�`�к�L�w#}�AC��K�Y���QOQ߷�@�5��}��j�H��s1N"!��D_!s�����W�D�
���P�T&��4O���J����w�&��B#v��h[�KjބU����\��[$�)��Y�c�kP*<��[^�IBڇÊ�W���G]��$G/N��9����=�G�;�)* ��B���@}t��]ik�X-(}����EE�w��Z�f0�V"�!wj�k�1�t}�悀��Ÿp��܁�ˈ�~�����_�(5[��E��M�j��U��0Q���@%Xhm)ve�n)���Į_��H��v�1��?*~��F������DJ���`��M5���������IkZ�RG7�l6o�͛w��gjs��:�8�%$B�z>AOǅx?�y�F5�t����b�O�(G�v��n��P��D�j�����ݣ�l1gOC�c$���uWI_�}�����(̣�Z�Mʛ��5&�� c�O6���E�s������tf���7��޼��,�qq�:>���vV�4�u!
ȓq����4u4�c@t�)�Y��w6g�3�������t�"�:8o�W����R*j�s�t���}��.���Gw�5�{�pjy�I�;w	
u�k�mH����c���"�CNOb"ob�����2d���	�� !6��4�32G�R�S4MSk���� D�Zu��s�گǋՓz��_#>6��]�Dbp>M�*?�ߨ���Z��o��@�Q��Rw�C���1Xt��}�
]Q`Ndi�@�����Xw��yf�/��٠t������W?�R�Dq/�o�G�O��:��)��ʮZ@�9��y7F���Q�Fz�z޴�O0&�G�^��]�}�Z@U����R���H��+l�������aNo��_�X���`B�������a�p5s�:�ɖ�R8����N��/�sw�uTu}���(`zy�hA�rE2ǔ,M
.�6�'���&@ �/���Uœ�TTT���M���B,l`/�moHm�Z�ߦ��K}5���wO�ݹ�u�A�v/,�)�8�_[.�'�NE{[fP�>�J(�n�(x�Z�,�U۴��զ�}Ս���éU)<y2mA��
�[�v�a�����B\5��g�2��'am�-j2UQr��V {���oH�{�"�!��J�a��(�V3�!E��lm1ºmKO�![
Z
O�<(	��M��I;޺�vj��5������w�?�ە���Y����o��0�����m��-�c�������:\����T;z�?FH�i ��-p�5�C�3	�c���a�<���*v[��2�I���
�ڎioɾT~��p ��pv[�a0|�G�?l<������\�ɀd��tA���h�aP���Ξ�/��SNci��z|_�r��f�ٷ��4�尧��!�y��w=�y������`�#���!9�kqĂl'���#�����RJ�ߎ�ɋ���>��l���jg���%���̏�W{&���~���ygښZ�l�J�n�n�5��.+�m���dYj�`q�[�N���=��K@[J�k��L��Fl�*��Z<�r@�o�}�)${´�a�k�p	YtV����[�(�dq�y�������[H?#�\-lu$�K)�
H��W>�d�")���Y��	�R"�
��x���膶A1�0G@����.)}~Q,��Mx�9�������{�z���{�����L��?�^\�`��U�'"�9��ߵ���E�zP�gԀ�i�v�!���"MM�&5N����W���f2"��S�6��`�5d2��?�:�I��Q�<�d��܁�qx���G��U
w�Ȝ���k[;ƴ�$����.ѻi!�_lnɩZ���L���mzh̗
�N�J1�D�'�Ϙ8�����~	�a�(�5���X"مs�Z��/n߭�V��~8����)�W��B�\��d�$r��Tq6U�I�޻h��'e@O__H$�h�˛1�	"Q�4�ƚ"������ń�^1��]zXIQe��i�'��/X]������t2��nr��^��Ǘ30��P8���/K�2�D=�T<��܌8e�c3�k��;-H��C�rS8��{ǉG�z���U�g�;����8��8���>˰R���5���������������[�-^[���IM��6h	�����y���!t�I.�����G/�;ϥ��0<�?gpQª��Ղ��N �J�����+�� ��68��p��;z�Ɩ���W�S����0ߎ��~���_�����cev[����[${ ��>i$�Y��u8���)ώ�c>rmd/#�sK�B��%%�+�nt��d�H��ӓ0ni���
¹���uM�I��~��wnj����ou+�o.Z�eO�uf/S��K[iV��z���1�A�<�M	�ǷZ8��j?f4�^W� _�\���Y��a"v��錎�v*|��i�Jޮ�	�[��6�'��[)~c���_e׭*1L��b�/Z�U�fد4�A�!-��h3e����J~��ث�b���������?�O����d~�J�mL���s����x/u���i7q�~�����.R����2	���I´�J��9���fN��U�������t5��Cl��}*M�����F��'O-���U�x����>_���O�qrB����mᣠ���^onY���|�L�C���W �����+p�3���c��^U���I!g�����}�l��L�?��4[��x�����&�f�-����m��(k�a�Z�R����/?�3�\��vi���)���̶ 7Fkx�D�/�:_X���:��k�����,im���z�C�
�x�P�#��-��|˳g>R�`M�&�L�������l�F�߶��+n����(��3[�N7l�]-���j@��{4��%����6[��I��s��'�a����}��#zp�A-(u���c��Ǟ'��y}ƺ�fPm)�Ws��1�F��z'�ɟ�x��u��ڟ��Ơu~����+
}r���b��m�z���}�Ů.ݍ�`hT��E��	�,�Ii�M�����-��m���2��K���o4PF�w���Z0q�������{>���l��B�E�(y�v	��GE<d'1�tК��+�w���B�y�Z�ϣ���΀H�����ѫ�T��b ��,ϮH�4C��Ee�<>�νL�r�7�?�p9Ļ��z�(`���I�\����qgx�]�+Nf����2�u�^`˙W޳ф�C?6�JƦ�j�'�����=�d�Xh���B�,B�H9%�)M��]�r�H�d0�6�_dv�����ϟL��m�a�3�KcD�w�)R�x���\w����_K�ڈqhm3s��hQ��߇R�(V�p�9EgZ[��μ�#o.?��WO]�����a��S��Z9��XsQ�#My	Y��t@UOZ��W;�3��Ub�Q�1�L�۩X�#�C����a�hZ����Je�!�+�D	�;m���C���ug�w.�F\w��H���kd�KǛ�N ���(f��z ��C����@%��D���u�z�|l#�<cGS�?;U�RP�Z�賃�{
��|�����I �����)�ˌ�ي}\�/d]P+	��:�H��a��OG�W��r��A�ese|w�糲����n�׍^���w �~4�WSW�bt�	���aܕP�1����tw!	�å�x%���?fIM�e��n��ƦAu'}ME|�(װ��4G7�H��TM����W�eh66=��0�o�1�Ю���-�FBD��i����"���w�ќ�C?��(ȗ��^��)L��\�li�I䢱����=�%�W�dd�lF�q�j"�W�(����Q����I���쿹���r��`��V(��9L!�
� �f�m��5S`���L�%$�T1��6=׿0Q�lm̐?�5Ef����E�MY�~�G�hN.����k���>aJ*�Γw�����1���0�/X�h���{�U��Uu��^�����%���T9���n��'���2�D���s.u9�O"��ʸ��#��+�^��=G�'8��&�@$K�AO:�R�"^կj(� h��`�/�ۭ�^��hi���U��q��D��߄O;Y�u?��z�g&�,�S��{qJ&兗	�Gg
�쥠i���F��&��5UD�C�!�#R����������T����ć�!���c�uy�\���)�Gx���:��W�kP �<!���$�����B��&�9=E�q��2^���T]`%#��Kf��	�Җ�F�d5��۷���xe��������\��z�o�\s�'��[�(�*�:���p���@
�y��K��� �1�
Wvz���XR�a�OpQO��{��w{	L�̀�؇Ď_�J��ϟ��9��p4���|	)p1�Ic4�E����1���攢����m�J�Yo�gH~���Ʌ��	�Y�9.�cs��?E���|K��9��iZP;�f��������:J@�B�U����������H�veX��j��nط٤[\�R@՞�G+>�`vIzO���� =��pp.��R���Ԥp���zSt"���3��!�KB�.X}��sQ�d�&wϹ�M�1U�i���#'�Q@�_Si��t�4u���|�ΜYh���
p~[��K��Q��*�\4��c�R0]��L�]=���ݩy��.壁�Aذdw��v\JCI�}���	��"�e���A��e��l��K���@�"vƜ�����UB��e}.~S�$�Q�-���ͷ��r����2�2�P�k|�Z�z�M�O��"/@��r���v��(�]Ϯ����f� ���C��Z���@��>+���^g\[���A^��6�u�[Ac�� Βc��}G����P{L
YFٞ������si��� y�ú�΋�_Ek~���kaS"д"K)_�tٙ�ʼ�
��ݾoF�)V���ӣi}��"l I�9����a%8Tr"sw�ߚw8����\q}?\S�l�zL�ܸ
��k�6�[�����í(�� �%�^��>n	!��Ied��&X�>β�_�m�Y��r���zB!��ػ��,����J����IWt�F�1���4��`�u� �@��K�r)82��/:+
���,��g-k﵃��	���E�O;N~�ߦ㍢Z��C��P�bݘpI���T�j�l��-��](pr�]*�lU�h4
��6��GdtG*Ċ�Ԙ�a�mC	]W�@,cm�,S��э�w�lJ���ܫz|�TZ�{׾�X]���<,�2���B�s�2����Z�%��n��R�����o��)պh���(��њT=��s�z��[=���:j����>~~��<��~���ȝt�6�B*-����y�m������
w�@�!��#?w�{��?,o����;g�^���B}�G��b��B�e�"���6�d�n$�yj�QV���G���x�<2#���A��_�ܼ-�LL�ON`���Gtf��.�u䨹��Z��E���҃w��%��0��g:���ԡ�#�]�1�B��6��?����	��@x��D��0*j�~R�/��Ĭ4�:7r0�v~�И��f`
�n�$D,��%2���c�9�9�$��9p�RՋ=R�����q�/,}ƕ��Mwެ��Ђ|X0ϒ
�Qͨ��Z���UTxc�.�a�z�	���K������t$쿝#�K9����I�O/���J_No!��Z����B��[��E�Z ��h��^_��o̮��X���y�q����ιݧ�#���5���:�W����8������o�4�����F�.@�V׆=�o{'�TE�y�����y�t˶k���;)U� |��(�b�&��3���?��>�\��tQ�K�D�Jr_0|r2�Go9D��)�A�=�:����5I����_(�`m��ϳ����H��=��º�=�<��m�"��R�:�-�������yF��b�51a��4a��
�N�i��X��.�}�餥A�n��I���P�g�X']�.��;�#�Sk]���`+��*c�[���-�.\\�T�&ި���l����|z/�Vh`M�
���m�0��&)�~d���ڴX�Tr��Z;���,vw����M{��&�.�-�s���������5K��g��(�ߴ㊵��?��?D}�C�_���HwH��ҍ���Hw���%HK#0Bi�Q@@j����#~��}���ٹ��Ͻ����1�Qw*qV��T�WB����Gp��?S�6�hb,͝���.��[����}�Ƣ;�y�D��ey[K}��3^���Ӛxk�F�no�:�l��H�2]���������Z�{�����B���U�1u�ƅo� ��AQy=ܪ�
�;R��~�a���RtR�磳ŏ�:��A�h��â`+����ǻ��y(�Z��V��78?5��65�����[��8"4���%���9{�+c�h����~�����㪽Z�P���kV�h��46Ƶ$�Q�[�j��!L6빥jo��J�`7���*��'���������_�.�u_�}���gF�^�ٯ=[�K+g�!�I���R,;����ߣ�QJA�iU�J�
߃7ݛ:��1�n��	���f0�@4<��DW��X���,�i�F9���q/y��C�P�o	�d��&���
�b
��w~�ox:2~� 9����4�ڮ�Nת6�
�nJ�NdI�X�m��w=�˳���ݞ)7ܫiZg��2�>`ˇS�T�n�jl�J��n��#uQ`��T�k��&
t�=n���x+�!�iį��%���}�F�q�V��8��45�ڪѾئ���Q*(������_�9�Ȳ�7Q�!`�>0���a����r����WM�_#[�b���]w�͏mz�%�[x 4ި}��ǉ���k�A����Y�Xf=���S)��Y��~קPC���ˏ�N(�Oa|�r���_���GK[��+�au�jc�PN6��ܱ[�y�ޅ	�j�� ℏ>t���C��]��j�4�v��xo�T�B��=Z
6�J��)���Y��E
\p��P�V�����Afg��m�>[�$�9̓e�F��i]�2D ��m��S�S��ˏ ��-����,�Qn��|�}]��<w��p�#��U+~8QlY���*�?�h�o6�V?o�6Ҧ�a/�>�ϠA܀���+�D*�7oE�u�ju�y薿+�奛�8����e����G�#� ����^&�B�]9�R��A�o�מ%���G���j1��"@��o������.��F�΄A���~k6���1j' ��bK�ܕ���~���.��'���H��}J9��<�\�yw�J�Da�V��(�J��O���^J���*rfQ���x����D��D&1j�Q}���Z��iSK�'X͉���9A+�����-$AĵU����ϥq������<0�!�B���_�IKzp�Yj|ZMhNt�����-��v��1��f9�/�������O�F͸�dS�K�)&��d+N�b�J�G�b	�;�#��z�}_&X�l6�7~T+N��ia/x1�bлV�ld���v�]Q����x�BO�O�C��̑} �nB�;��뒞�t�ن��X��/����x�+����w���9%W�Iq�M�Ո��9pU���?b��ʷ��j������f���6H�X,[^C~9�j� �$Z�G^�����̼���EaW��Ȥ�+Q�:(	q������4��Xqv�}q$��m�ɣ���?�ܞ}~j����ϼ>��G�+Y���c��%�Y,�R]�L����*�d|$̬AO\�Ig>[H�6�hS���'WԌS��7F����}�|�E��Y�B��4���w"�H�L�r��e>�7�#h$��)���\�5Gl�c\�>w�,�F����KݗT7g����������?o��Z�ϴ޽���`TιR(���Hz��f3��� }}xݸ�>\�9�&P�U*��=V�S�xk^j��{.���!�@ۅ �O;			�n�W�>�&����
��ݭ`�d]	�L&l�����,��YZ�S����}������"�8�%�m��Q�D6V�z5m��vJ ���s�V)/Q�J�l�\0|W�MF�[)I<�����ّ8�o���OO�GĂߢ�m轷h3�x�_��%ާ�OYG���,Yxq��qJ���7�?�(���U��u<�e1��}�2����"k�]it�~�#h��'��x��tq!���/�K)��`����/��`WbA7��;I��=7�����h�� ����z�ېo��#|	1�C��o�b#R��|:�#�hM׷�S�K�X}<Ԇ�&.��4ӯyEog�M,a���[r�[�<��7�� �@�:�6�v]'iw���:��G�� �3p������]��j�Vm�ʻ�°9G��j�h���&ǚ��
!S��]���"ǎ����%p��W��_�d��!30����LB�n*�b����~��T���8r=�K���腀��x&e`�`Ni;߷v7�"i��v�	����U�Քi�7�y����1Ą<��|2G�+f2�ކz{������J�#M��^�6f�c�$�l�?��z�@�
���\��,GUb���Y�:E�����/LsD���Z2Q�/��bz�t�(�{�O���"O̶�>��|�f��;�����Q��\����T!gՎ�}s����4����V�'�y��a+�;���ʚ�g)���ge�X�H�zԠ��L��ˣY��7���L�]�;P��ޡ�9b*u)�9Z��%8��dLx=&�p9�x�+
��>m|a4Я����#-[vD�]+C�E�1�*V �%,��,
c!mm�N^LZ�kA�k��/6 �EE��Nڔ8һM�ǔ=� �%с�iv���҂;mQ	j�D����c/ϭ_U+>�}߶��^^���t���!�82?pw���[#�x�z�m�x<R�%wM[r��c>n���ͽU���[�9a�͝�ư��O�f��3�U�M�ir_?�MM!�����y����j����N��
�;|���%7?{N�E����Á�>h�v�tǺ������#�Y�� ,T���ɏS6�����`&�#x�ɒ�X�<D0��Hp,�3�sٶ'ku
���R���#�#�a���f�7���B����$���񫳰����F�8����q�{!�%���7��}��hDa���@ -A��Z����l��9d̟��n.�
ɷ���{��6Pu!����fh�dp[��f����޿q����s�"������� G!򻶙<�~��������2~=,�a�=!�k���?�|�B9 &�D���0�:������`�OF��'Е�H�þ��E�f�@�,b"�ύ�<8��Z���X^�J).Ր��M9���#��u�)���,�>��2����ɼWÄ䩂���b�3E4����y���b���n�tW��[��wx{N�4�q(86�X�%�f��#8|ʶ�&-� >�߫�%
��٪��Wj��4>�7L57^�.��-
� ���?��Q5��	d����4��v���$3�f�c@�_���24W"Ƅ��!Cw{���w������� Zt-y+^`L�+Ǽ�bɔ''��o��ױM��1U�͆,�-��\���v�Ǿ.:�jN�)ܜ�'g���έ�5���1@�9Ύ&��]�5����{�-���&�R�f��\�%�ꓩ�4���e@Ց���4�ܗ03r�.hp^��e���筣�[����!�(T��m��P�=i�EN���u4�$$�ǫ��p|��/�%�A��rv�n�������<�1K�?冹�ڊ�&��̚֎16Y����6*]ND#�^=� �2��Q3��v���cvӓ+8�Pg7{X��4�L��Ī�_���66�aݮ���K������Z�
�J�������3��S��C�GP.
����r�!��X>�骴��Eܰ��(���.m_I��\�W?�����MP���hc׭#�z[%��fDbO�~r�BAf��; �m�}���% ��7��m��TOL�*�+���t-o�o�;�
�Y2?��[�%��&uX����׾���~�YܘY�߹�մ�n�>R)q�=�����;�<!����]K�f���`�,?�����42٦�|��R�.�@�z�-�T����H37D�}�%����2����{�������5˂���f!r�����XU#��W��6��+�yH�gݳf�-�1/����9�g�_��-�Uඛ�D�;��ň.V�n�C1�oM�T>��|��o�<#V
�v��l��S����k0��K˒��n�T������rAx}��>"|��~1���^/�?<���L֫��Cͷ0P�{�ogQ�Q(D�όpe%������^���"3�#�S�^M�y��cnc���T=}l/@h̜Ou���L�$uϭ��1����:7Aˇ~�vLJ2�$Y"b\ԇNѳ��2����u^� �5y�.��`��H��F��(�`��l���6g��C(��fM3$Ǆ6�
1�+�wG_C�
�wA��.���8@=�(��� �÷�wUp�� ����i�s<X2#\0Ӻ]��8���W���6�-V`7!�i��v6��8�9y!�u�R�!\�g���#��&�/�NXӚ%��&��{�-�~��	��t���A4hgB��Q\)���c��!2N�N&� ��6�z�̩�Q\��F5�Z-�(ˠ��O�[�9�<��7K���r�7;�g�ΏDH�=3\�g���w���iIm�Y&�yq�^��\�������G���'����	�v�?(��F9m��F��>�}U�7O���(5�$(�gN�/��/_�֭���_3��<9�	1�kS��z1�>��6?%pz��]�B��ԷY��������h��Kp}�E*\���,%��رT�J��<���RI����4���P�L��a�>bŠ����8z �j[+�.|:e8+��o���ɴ��#���Uo!�g'-�bPy�g�^�w�<9?`�O��Dzh�4����J�l*��̦u��(�����M�%@C9i8
��Z2�u���{nI%���!۴W�0�yB���#Sґ�O�al��f�~�4H���H4�JP�����
CL�R<��1"�����V�3B�Ww�h=n�L`��8Wd��!�v~_��vJX+��e�� }d���Po�b����t��� '8��[�<��`��»ک�r08gAUHٻ�$�ܒQ�����u�c�9'�@�G�����M9{}m�.�WO-ѻ�V0Z�2瘘֐+)��L+ˎ�%l����yn�<�eXuuuEŸ��@���jV��ɠ�S�z���!�]z�E�2ס����%9�\��q�48�I��c�T�,�]�{�^̍���j�$>��T��t��/Tǃ�Q�D6�v�u>��h����h�._��.�oў�i%Ɖ��i&�B���w�v=��'��w�w���%�����Q�{
�M����g�݅�n�H�[�B�dw�ƾ��w]rfy����uகX��/B�W�7|���ܜ��;I�(�H�D��+�Τ��{N�&V������!�D���{�U��)��0T�b�W���(j���S�����8n.�.����Dp]����G�zM��5���Ds�mj�;�B-����s�嚠���b��A������̄KY-l,�·o�u
�����t:}���ת�W����T��~��,�>3��)�'�i�F���0fr�3���4k��4��ڵ1��<�,��Dr�1�v+�����N�;'sp��Y9�������œ��5�M(ߦ����Kt�i����n���3��W�.��su�e1�}��xh��j�����&x�~���-@���-�V)��L~�'+�4F��sę������}��qp�����VV�F���p�i�hO,DK#�Q"��>jQ���d�좓�E��C��l�j�0�-�o�e�r��Z�m��L��3rW"���q�kB	�G�1�%�%!��J,���<���g��l��<נ�B��A!�m���*Y��!|��̄������d�΍�M�:�Ĉ.>��B�n�v�+@�9��5�e��i_q$��>3v��C��l���������Nѝx-^O�&y�Me�������������Z�)�����Z.�g��2kb1���-���>�6�:�|��V�������W�ir���Se�������:��+Q���ȟ�;<����|{��g�e�嬹�%����7Rc5~mf%y$�xL��y���>�\/���<hjQ?��#`��}��p�>}��W��K蟄3��V��ޠP���"-��њ��C�ʾ硸���o3ǡlC�<�}Gg�cTϘ�l3�S�o�3��yvWbփ�������������W�
;�Ǟ�A����U����y�?`�7ʛ�8��c�J��錏���g+I0��}��[e���<�#�M���1Ο������,����t'��������qu�6�/�Aw�,�� ���>5<�f�� b����i9*��x�<2ʆ�\��N����B:��mx =�G ��%	"|}%C�7K�hޝ~�}�N�,(]��9.��C|�{#I
��b !��t���Õ���`��iB���p�����h`�,��w���K˒J�ar���7O�cnV0�ͪ�ի`�b�o����^c�#O?�S>�4�.�ߗF ���`�-KJ�	Y�i���]?s~>)�
�&�~���1�(�+�8n�x&�f4��)5a���6J�*�r-g?�b��	��nk��|����?��-yZ��LGi�(��>�}Pڽ��@PR�[����Ä4���e�z��;nYA_裷�#@�u^�/�',7B9
�T��A�}�S)sV��\x�6\�o��{u����ڵ�����]�H���o��Y�4�a�p��
���C�����g~ۇ��xt��u�ѬG�)k�	Θ�v]�zQ��8~���:���Vk(�S���q`���u��.���7IO����5���"��ݸ�i ����bK��#�\��D$�h�uz��>i���9jmo�Ӑ��3�C�C Va�Gɡ�c)�X,'l�_9���`���W$j��VŉK�:	�a>@1W?�y�+8�KY�^���tb�1�{�ڒ�;�n%�W�����j�l�n.�gۣ����˷s��tu�* ��>}R�kx3�0��U�Z�<]�&��y���j�-�R��"k[Y7��4����l6������q�B�'��3N����� ;�WCq,���ߡx�?��k����]�X���t��?9vq��\e��19����AB���?J'ۡ���n��U]���'��rK���B,�-+ZO�%Y;��A>����SM8�����o@�`��>u>z������-nP?��4:T���#-����,��d�J7���>�k�4�u�0$�=D#`y\�5\�V,x&1������5��Y\������0߼E�װ;<���R?�b�#z�/K�,�t�z8�'gNB�l��;�3)���5m|vfq�D�����YI�]"Kw�����Uɲ���qB|6�8rL�X�H%�|�������a�kn��yםe���;��5aj��~l��b+Xʵ�c*<8��=B��/��;���29`���[y����U�B�\�
�wF��N��w�Қ�n�Ar����J�A�:&83Zc�i����:�9���9!g���"<h=�>i�����_�V[uZ��Ja�PzctP��#Cu����>�vq�+K�}����.9��}'r���c�.�ߞ;v,��ڹ4,=n�����εa������qd��h�r�\Ġ�����`N[WW�O�?��w]��__J�X�
�elX����[ *�>�P�Z�	�$�׷z�̫ߣ���s백=K��(I.��cET�۾�7�?��Rj�T��g�m
Z�B\�ۣ�-db���p�߽~�6(�i��ҽ\�~�Ot��B��b Q\�A�ū^���]妒��>�WJVoS%:j� ��T�8p�x��a:g�)<p�啚,��©�CA��E����;3Ä���F-LM������=Q��ח~���ah�_L��)��u�,ٻ�w7����]�S�#�P���}φG�/��ϖ�/|�0��8�E���3�����vm�=1,��&7��ˇ���ȼ�{��q�����r�/ͮ+i�7�����&U6�cy>��M��wK����Ĳ�;~��%*u}��_3�����V�Ƚy^���FH��j�u�S� a|�掐�}��@_����y���l�ۦ1�jL`�v�s����4�2��6,C
��g,���C];��YS"��C+�qe9Ø(pR��%������O�Qӓ�%��-�x.Ó', ��]�Ӂ��7�˲~!C=�8W������!�SZW��"�|�/O��6�J�	 3<�C75Օ*�|K����6�[1[�l���C��tg���2��o�0���Y�:HuE�[R�;qoKp���R*��Y�����_�������[���C���]�YB. 6�_
n�tB�2�;�j*���H$�~�� ���<���5Gl���^�|�})1�͡*-�{`�v�S(D��v��9���y�a�) {fKt���NC�~뎝`t�uЍ#$���L,�;'� }��ٮ�{8r!Iu�dNq6
ܬ��)����Xܹ��C�ֺ���Yϐ�����c�?�'�Z[ˏ���߈�/��-�������6�^ط��	��M7?B���_��pgD�|�W V�\�V�đnX�pN�{����-����B�h��_t��g
?�n��Y�����_C,J��	���/�T�߮~�^X���/��S�ׂN����Y�x�<d���^^������鐫/M����/X�M�P.�=KL}��xu��a���la�Q�d}��i6&pٵq��7���?a~��㧷2���GR;7��f��>��'r���2.b=�UC<,�o�}��4��H�M��*�� �:��p���Ql��S��o�0	,��?��-)�Q��/{���9tv��D��4�P�|�0�{�rʧИ�#�O5u�˫�K�(t�8$�E�x�W�Y[/�Wm 8=��w�۱ b�R��!~�iV�<}V(щG&����!���I�Z�@/D�3M}��v��x�� ����
����]
���$�K���Ds/
g���US�~q�cOK��d�����QD�Í�D�k+[�3�R�Co(*l�t��]E7�@���g��%�'�f⮄caƇ�Z�+e�F6<g�Q�~?�(���o��\����憐$�\��ƌ*YO�g��8;�g�/}�@π@d�ߴ�i�)�:�g���!'>٬��=\��������2{̅:�;�,�<uZz�k�@���,yo+�a>�Z��0P>�h�8V�iI|�e�Vi���_��ϖ:�Y��Y�H.�>h<T>���ؗX��1 a�5��;V������]��D�B��ls��v7`���:�i�} ��p�{ܐР���u�J����x�����?u=�s�E͡�/�T�S<���7��^�7�9�!j�9�%�9���k%$�0I.y�3���ս׸���V��~��A��"�Y��sC�8qୢ�Nn��"	��l��0t��cV0�ur��6���m]	��
��p{`=`�X������?y`�<�K���^���tPx,l�/�&1�z�ǥ]~���X��^�|uv]��H�L�>t��r ��t͜����|��7��5��?����t����b�vJ���~��� ���z�"w�{����~$������0���ZY�»�8������*�x�ު�sd���_�s��(z���:N���L~��y��BYq��P���@ŁΓ�_�l�3�El.'�����{dԾL��:�W�"[�qZԕM��E��!�4�T���Q���yȕ_��3z!:,X�B���\x.SZ>�>�"��������r���X�>��
�NI�(�_4+��7���h�1�����M�`#օ����mc�X<����ٲP���1.{_+���|�JQt�[U�t���~��X��V�3��e�ud&Bǁ�L��0u�*��K��l9f�GKM���^cB���P/�>���N����A�s�X�]�Ma~�Qƅx{�^[;'ٗX<�yӾ�[����N�"�/K��4�	l?��J/�i�MЍi8�6��!�kq���x}��aX8���9��O�}��R��*P%�̤�����Ӂú"J[^I`�`*�����sD�M΁Zk�销dM�)��p):�
��.��@d��ϒTӔ���[�0l���u���)(��� OuS�5�d ���3��ІS��A
9�*�j^'G2	�t����4��ZeO7H��&����'^�E<;�����)�I'М�����=^�[x{��6��؁U^~~ϕ`7�s�[(�A�K���q��&� �u��c��#V���"���	�{�t0g�J�=R(�P��k�2O3�O}�M�d����]�#���Ɖ�/��r�1f�1�������ފ?��~�{�7��n��i/��ÿ�d=��"!)���V���?�I���j2�hB� ~u��YwG,*���A@��ר�V�5�0�P��_�΀�yT�,����I2\P�*�+�����T5��Y�uk2c�Hm�5D�ѝDL��u�
���-���
D��a��o��x!��Y%oK�a�6&c��~�{q�;���^O6�Հ[��(��y���Y��+�"]��36��p-������Q>��B6�H�\&f�8�t��Q��T���"77T�k񆾚��{�4��P�Z{����r���(G���Cj��2M��G�"D���Ͻ2{��;Z��R����Ƶ	&:��w�?أK�àa�8o&m����W�ZC�-���$+o��zT;M(T�2��!�����K�ӱ�Y��6�rڒeD���5���#ڪ��YU�h�e��~r�d��nQ}��^�?�u�d7��au�S̘��8�:��c��J�Vi��f(����΁�ņ!Q��Q&��B���?S�F��(��W�m�I���3Vp�oz�1�y�� �/^�]c
�
k�ϖ�f٣��~���٤�80R�?��]�&�4��ـ�j�Qb�@l	KǞ�r��K�Y��>�^�I�O솸�W�y�>(��ـf�%�r����V�+�3#�5��������%� 	��m<�YO<;���?�j��u��uP8�)��ږ�%�'�x2x���|N��(�l5�X�`�����7�yϣ���c�-ڨ��3��D
��{��c��q8a�6�ÔL1gR�䕊;7ߺm$��>�if����թO�������ԥ�"�.��Z�W"dl��	���e��3�Tt�:*�EC����m��u��\��ڣoBb�i݁��Th��&����q��/e����WP�{SryKBmۻi�&�"0�����xk�E�[x�z�ۈa��K�d�`�h:R���xv�B|�^^N2I���C[��X�߂W�(�ؼ���WI|���]�
ݾ�'��͐�N\z+Ι�Դ��X�x���� ��}c�񣆹�68{�jGF����F�*�yΣwg�I:�=FX� d◡|nH"�<�5��{3��R�>���E��4�T�v��+r�=F��ADσ��jR����OMU���:q��eҡAo!?]��<m�����G��W��آX��<YhD�G@+54�J�eL�%��,��-�Ӓ�*nֹ�TO��Z}���&���˿��E��p�r�����x�vZbY��
�
5�"���j��8���`����m��Z��F匆B��=����W�|@M�܎:�ÈO΁^Cee�ɗ��P��_�Q�nO}�bD� (t�A��ǘ0?��'{f	�&���Y8�i|��~�ʍ�H�y���)�W'�$�v���L�5�v�Ԛz��ć�K	Z���1��*n����iNX�D���}��ϞO�O5�
9��yզ�a��Z�����.�|S/v���Y Lv��t��+Z�>�������V�@ ��7.�%�!���-���|c��G8J��H�_��@��n����\����]�j�KS���=�	8"3���\r6�Z
|pcR۵���S�C�y힪�g(04��=�d}�=S->+���ͬn����~���{G���V1\5|7�O�i��!�\5�.!|rRGBJ�٥M4�I[Z�.X���M�p(��i����c��;|K���������Q!;�j�z�����pZ��X��x58�+�6+90x��r��t�&>����m����r���+�G�\����f~M�hw��/�N��,�,��w��D�Hz~�>�7��&�?+���0Mװ�a(�pS��+�ey}|CU�qI�km6gV���j�S��*����WP��hA��
�3�����e�g:&�g�@�ڃ��n�K뮖�,�8��*2�[>��$q�h#cr���\V�Nĳ��~���g���f���'Jϱu��M_��#�Wy=���v�Yy>���pɺ�S���.ol8tS�v���>��ES6ì�>f���`! J���<���y>���X ,��:�󕵜��Ǟi!��Ĩ*l�v:���q�,4!�/�i%��� 8�ִ5�I�>������'��d��=\�u��7pm�#*����k�n�$>Ko��!bԮ�f!���/C��j�*��-؇�@��H��N���]����GO�Og!N/���@���ֲg\�� k�a���H�:	��1y��k��e����g�c=��~��P��T�N�r����F���dE�n���dH�<�2���I�]��h�Ǫ�O�*�{/ķ��H�P�#>լl���[��䒄f��)A�Y�۬l��P����x�-1'�/]0�#�sT3nn=x��4�ͻ��L�f�t���W:�p�h���d镕�w��.�v����)�r̰_!����ׂ����nEWx_ߴ��PN����3���֐�����Sb�|@�x��W_��خ�'�j�䬵6��b�3��f��M\�-H�:�l��y��T9F�CH>L���p��w���> ������*:JK�*�n%��z�)�е���j9�s+0,��=SxZ5�S�����/�9qC���uH�=\$vY��΂�>j��AyP����Q����":��GxN��ŭ��5���3�I�i,g�\�ܻ�ar�&Y]���K�	��"�D�\rOs�ʵ?dIv-�X�cE<j�)x(�������!{�N��L���]`�1za��/��r�>s�`l�3��oU��R��Ѵ��~]�l�Y�緭��#d�9�M��.+�������.��J221�~�!�}ע�&�|�|^V��O�f�\+�ajQ� ���"��ߴ�d���W��j�����>�w_��a0ݧw�g5(۲���gO"w��/���~䳚\�Pf������'��F��*j�H��y�q������c0'
�m��rUw�8��M.��Ly�+��.[]�t�0o��6:�\�,ND����ij�˦�K���g]����.$uQ��?"�c&�mD�"���/�D���ơ���q�r1��m�4�����[B(���o�^���MS6��0)��am"��N*V�.A�9�'&��yO�5�&g�o� �����C���R��k���}e�\�"п����15%��,�r}#�(W�u:�o���6�H4$"�����Qp��'qS��8U��,�y�˹�q�t߉[[3�9#�I�Ͻ~,�(&��^1���ӡ"�%��+����%�Bl�6�|�v��`�@�@����7f�6P���c2��V�d
ѓ}�����A(m�&��c�4)�nN�Y��.ͺ85�{AQ������INn�,��B [^�c������VLYc��"�s�κ���s��2����I@d��}3�L1�"#���^��C���6��⑋��ㆄ�2`��9M��;�`-�Ǚ?	��+��3�ڎ�W��7�\\z�<�Ӹ�����&U/�����{	nå�ӊ5K�o��U�Eh������%`��\	�Uǔg'��|A�� 9A\u�%��x�J��s=o�(��ks<��;�O��!9\S��!L(}�C�����
0�\r܃H�������Y��:,IP��9�P]"9��+��M�ц n8v!�1�C\��pi���V��U� tv�k] B�
1�`�n��,�ۇE�����0B�v+-]J�s[�.�ej����i�3�IL:�dkh0:� �:��<��D������4�L��Ǒ����D��@���X[��*6��W'"8���Z?Z[?�R���4� ,��y\;�G̓D���XcTk��K�|y�ګǳ$/m��N�Κ�޷FL�!
�H�������#M���ew��E��
�Z��t[K�G���s��-ē#�ڀ��d�	(���7���-A{ySb&�ۥR�י��/	~hwuer����8^'WZ�A�9f�����V�9�@ d��O��8�	zT���^����9P�S����h�s,^n��>��F=��
��Z��j��2\=oY��wc)���;u0o����U����冱��5�r������m`�o�\a<���Bۂ����}J�JT�1�~J� X�R=�oa�|�ꖹ�W���������8��v��u�]��j����Eu ��Sjv�Q:��`\��8i��[3�*Y�W8���tי��� ��n$
syW³d/~h�,�m�H�aG�����g�a��Äd	��ܕc�Zv��|�ѯ���S({NO���?�+�%���oʝ�\�[V}��\-3m͏����w�ȃ39�d�~p=��(=���y��Xt�YN3.��9d@r�u^S	<��e�8�'�i��KZ~�t�|�8Q6.�F�37ҡt��a;3v�Ό���f]w:��%	l�ݦ��{`+!+�/�o�{��o�=K��J��@��tP�� E�p����x�=�.���<kX̕$�kd�B8�Yª��ȗ��pn��~D��i��|��M�����y����9����[�x#���apޡzk�p�B�q�䓘ʒxq�摙�II��y\��C-H"��~�I���]�P�QUK6���kh�������풛	v��&>T��|��tN�����)P/}�Sz���UB�h����(X��F!�C��?�ǔ�4����&��SI9{d�k���F�=2�g6.�fL���k���=��n�ۺf�� ����ʌ�+S7f,B�YB����m���f3(���F@ypch��� �?T?�۔8zm��Q"�����|����;,��,z��³���I�}�����%?�����!�x�2�c=��&=��fr7�E�3�P!p�]e���$	iX(�W{�x�$�M�^]2�oY`n(�X���l
�8|�Z�:�)n���e���2"1Wj$�ړ�ҜK䇅mh��!���"����r�lޡLh�)�շ�>s���8S��7���W"�3+L�<��;�����5��1�(9���riR�l3BW�e	���4*zęx�V����7�,�X���y?�*��>��^�;=}��M�,j\����갢�c�G���c����c�;~nl8��Rf���_��q�ة?��f7pә�0r�A�x�]���?��,}�ѪC�����$��;��:�/!��7��rk��y3�8E��%[z��b�1`1�}�9_LKb7��{Sݪ2p\�4�<0�ٮXF$�|>�����/��S����a�0����S�g�;=����p��\\j�+e�+_c��F�,ܪ�4�6<<�I ==��|��ٯ��W�o���Y�ԃu��S��w�����C��/%�l�3/�]�ѝ� �~Y@�#B6'�ȹb��PC<���s,�Q�q��w�(g��Z)��/#�~��+r���$	�+�Y�9OT�h�h���]m32�~#M&����"�U�HU!�g�uft��SD.��/OpIHH�Z �v*ߒ�U6�~�W;x,?bOU �&����(���H���!�qx�P��bš,n�(�h���c���
�(Q����\h�����G!��3pH�o)�X}V�>{l?���z��dB7c ��A��AG���/ j�:̩ng��-tf�p��Bx?K��K�Z ���
�ރ����q�1�`�cd���?�.y�ϴÙe������ ���6U�s���b�tx�ҥ�..� ��7�xO��=4]^��ObX����2q��mp����J����o�)/=-����f�~�?ȃ�/d\��h� �ӱ�Ojv��&�ȑ?�UCW�Źn�i<T0X�������w��X��sag�t,�ΐ��t�����u�uXj�5t�N)�XB�mB�
�eY�IU
��tz��v}�������GC\��ĭ���\*y�����?�����9~T�g��̖H7.���4A�`�b#7�4"
�`��p^�Ҽ�p������x����kgK�Gvv
��٣��+�ڛkK�!3�{^���&{^\�^Ž�������~�����<�3��u�Ё �.Ej���y&r)s��_�w�Ȼ_�I}���g�� |@p�m���}�ƞ!�9�=�ܚgu�M���w��i�/���b��F�܃8-���?���5-A�̷��w=Rz?տ��c�!��IoVP<��ޟ����Ūb���{q�"X�R����6�f=]�f���uTi��yCq�POZ�1����/���	�q�۬2�K[k��W~|�(y�I��������p�>E$u��vJ!D�o�猅	_��?vEw����[sgb�2
��֝��̭%��݂�4�\�Gy�AIOXM(E=$j�-�$�w�4�����Kj���;�^�P�۱�R�����e�Ֆ!g$�~���^�`�K�[��
��S�|��'e�3߲���T�:r�>Rm��iyG=�.]x�R0$���e�������ڂ����X�Nֿ+�JIN.l��aD�E���g���N��֣�ݖ�ɂ�G�o�+����]>��AF�2� 1�ެ��oF��������]�Ѕ�)���8���5'CM�x����\���Af�v�tY�s��[��F�ɪ�B��O�.$g����C$Hp�ő��R������(�6Q�9�Y)�����-uk��jg�l�ܿ�P��Vyg��3x����y`�Iv.��=���AJ�Cj�j/r��JĦ��c\�ε�bjdԸ��m�wcǺBLZN����]�,��[�?�<��~��J�V:�sR���{e�? �G������p���!���j�����V2�߰C91(����;1�̂���y6
,w=锔|(��!=Z��{e��@�O��6���AӇC�l�ec��ם8�
 P�s"$��I��F-��#��2��~j<�q__�V�{�:]Q�Ś?�����i�y���7���?��6ȕ�|_v-T7U}ٕ���������eO��,���<?��e��G?����%��G4a|ҘHԓ��>$�x��vaۍ���4k	��/;�m�����؏��^��)������j��=ٵ`�59�����"^���i��$o?�[���X[s�5;�Z�f.��/Pe�La�\��x0�\c���8\�15oM XR"�U!�/����0�+m�Z?�~����udtƥ�у��Q�\&�!��i�{���t;Jˑ���Ia�tҝ碘�>M6n�g1����L�&���l�m�b2Go�WH���֦��/@�z��O�&N�)��J�dHj����Z���hs�:����v[��t�uN�i��W�� Q�4����;�>��z��w:_��:���?�2��*Q
�er�c�*��;�~\���%���ҝ�
��2���:D�dk$��6������[zX�"���GּD����pt�5/7����5b1�~=��C�C}e.]��6��sɘۛc]QZ��k��=�(����MHM�i.OT-�^����>�O�QE��=�@�wd���H�^!�&=*�]�
�\�ꡒ� ��\�YB*�	�];�H�m6S�:��܌Z�SLt�/0n�n�g4_��Vs`?�w+����	۰��%���J/�~�s��` �{9ó�,ϴ��FJu����d�w�|TG����7>8��f�]��%��tD0
�lJ�q�����g0����!/nnO�mj�N���L?�t�ŀZ���utuVwa���k�w��=�5안����xl^Vd�<	�"���e�󖖵�,��Qv7�m1�щ��-b8�5
5��O�OB�Bv5�ɾ�务��Zd��	ɟ���!2��������))ZW�T���1���Mؽfb���G�'Yr��v9��ݭ���/?��;3FѸpg�j��5"4Bv1fC��c��)�?��\�!����y���6,�u+��y��� ,�f��Rǽ(��N��UD.�I�:��)_��a���(�;2}�6�A,eٳ&s��Vh����`�A�|���(I��j�~y��E�\�[<��k3]?�E�<Œ�B^�����k�T�tp��	3����+H���ױ˫�v�*@�E�/-`2E�5����h�ǈ5�і$����Xk���}�V>P���D`ȋ�"Y��[���/��	^�:QhRA�l/�B��Ƣ+��~A;	��T�yt�"��g6E��9����*Sx�+/N�)i��@�� �9�Z���� ߐc��%�eW�m����,����ڗ�b�!)��QI���#�ѷrccDF�����G
4+B!�&�*I����*��k�~���-�'���rVƝ�O�]��\�8��)%���������]�U�� �tv6�U��)H���o�#6� 7��Ⱂe0�X�2�s�zR���Hf�]��+\W~l��N���?ՒS�	�|w�����`�]۵Ӏ�Vh~��@#d�#�ʘ[آK�����t�Re�'/(�hƭe����<5�>1�y��%n��s��ڽe�|?���&R|T����S�B���#]��C����$�~Cܱ�B�2�	�7������nv����&QT�=?���{��I���s�0�Ȣ�2y���|�w+ �*��#�'�K;��wٶ�A:�AZ���Zr���AJ�q��A��_�z4%�Ys���VR�ְ{�T����9��K޷ɜD4kN��Mb�$ݶ�<�B�W�G�g[�VUQ�ܓ����J�d&G�WǸx�a�6Al��=�d=*{���G0��F��ܰd����������}�U� ^*���XBj璁����'�/���n��^��M����t2j��J��G���j��_Fm�ej�)
��@�>&Ў~�#m�u�WgR�{s~���G�	��b��켿7 ���?}D����7b�N��vI=���Ҟ*j%cR�-�6
��d�P{a��Ǵu����1H��cE2�m���_S�zU��Tu�زa������
�j���А�	����T��ct���k|J�����#�R;��ޣ�B@7
���lz�A��K�\L~.��^kx8-V
��n���0�F����0��%1�,
7&��i-C^P2W2C��:HV����1�)9P�-���Ù�}T�LVC�[V�Z�X�}�a��/̇&�U%qߋ������ݠH���6���)8t���թ>* ���u3j���e�m�!Y���%�;m�A^�.aS�Dig����_e�#�ƅ��@������_:L7d��~��D��O���s�iä���a��"���X߬�=J���Y̤٥?���I��!W��|�
 ��C�u�/e���4.���R2�~D�S���0��e�m�>�zd�uX����,4��k��<ّ�����=���L��T>P��L'0��P	�RZMԩ��q�%��%> ͪl:X;��*&����!�D�sA|{�k�9�J�d�7���7�����-E��m�Io0�����"����G ݜ����
�S_�W�� K��k��E���.1��_Ǹ��<�u����O�QQ�O��,�U=>�E_>��n��W!�v�OgF�2�����b�����А:+�v(���#[[���
uq�j�:&��e����#���j$#q#k�lG�1��Y���]�N�2!;;{w��U��~��]a�G����A�DN���4thl�J(�o�������\��,B��a}�<���ч�DXT�>J��C&�K${>���g�V���&�$�K�o;f9�N+��0��r����T��Xfy��h�X� w/�I��_�'���/��K222S"���cL)=�<�l��7���o]^�'K
͊�g��Q`j�����X{h��p#��G�i��5����H����C�ב�;�h��v�C۵ٙ��I�C���Y���>��-�r���)#�����-���F=�����r}��
e]Z������C����BN�S


:�$����	a�{������'Fa�Mu�G���7p����Q.���D2����#�#TxM-g�״?�&=~���%�A�k�i�ܲ�h���Q��VB��l�O2N^��E^+��>��D(���i�OXJ���`���@����~O�n[�G�a��K_��"w�������WO���;]�� �+�v����;�T�A�+�9�^=:k$R���UOl?��IP�� ��w��Ժj�D�;i��>�˰�LKQ�`�0O�i¢�`�� ��R�M�gɞ�M��m��W�/jʲD�o��Ny&��H<8%Zl��6�|a���,��������j@�0����<?��KD�C��w��/�GM���T��t��?os�=�"_��ĳ����S�!�����D��(ԥ4�K���o7�� �k�"�Y�Y�Ģz�pN�[�ޝ�Y
P>ftG����}�ݨ�l4�{E��:> e��T����dT&��c>�U��`��{ޏN��
��T5<� \27MM�☀Mϣ'�����������B�z�S���l�A|Ǒ�`�z~�
Q���
l�ހ�[�+7��'��l���B���DN������4�0ݽآ_.p{���+�;�ϛ�끕��1�'��d��eg�뙚hI��cG]N���ͯ)G�A�����p��:��كҋ���P"N��/6�L�C5���s�oIO�X�.~��+�j��� D�ġ$-2��Z�Ws5��Ni,-�>���lIҭ#��w<������rz#�$6% �M.C�xSs�r�ݩ�AZB�%f�N��4�.P��8�A���!/����sx���-�[�4��XV<W�u�`���n�KΌ\�!PX6���՗�.���.F�	�\�\�[u���|��`�4�^k"��Co�,����د�,}���|o����.2H�j,quoϹyh��?@�'r*�6�����-���P�7<���/����ˈ�o�~"q��EB��;��(V�;]���z�S�M���w;\�F�*������B}fu^p�# Q߿}�,��Sqe��n���@�̞<~H���~H�c;%d�R������`��\Rўd�h��j��|��N�UVg���@a������c�3���!�c`kck�ʺv�����2dN��hW���"�F6���<�'��\����������Bb&��������G�-(��[���RXʐ�#�����0Dsٹ���& H=q �ek�;'j?}�ob�u�5��:��A���q�#>�� .�����@��IY�� �Hz�f�m���I�E�%��Į������� Q�+��9���%S� ��A��:%��!n�F6f�� �ϡ����K��T��5����8���_!M�#�>�;�����eT��%�G��fX0�J�?CNJ>5&��HL��@%=NG�7�=H������yH�>��I4�ݽ�`�YJ{
��l��>��2���N}7� <���h��![��Ģ`���S`��t|<V�F�ܕ������V���a��x�90�%M�Z�7���v���=;��x!L?`��>�y��i�?��C���P������2Q�{���[�.��dN�q�I2��{�C�_nw�Di3���_����hj|]4��3z�V�a���i�\�Z��߸%������}��=�9ee�}�'sK�1���sP��|>�^j.!˵�7o,�����/���6��A�v����O{�� �U"���U_>��~��@�n����>����-E��ep��!_K����r��M]�ʁ~��T�{U}Q�3M�^��;	w�t'�߀�y�y�|7��F������C�x9��������>���vl[5-�N>�*�+���p"w��9)l������6�{mY�Vq��Qߙ$HqB���o�^��+���]��Kl��ݐ@�����Z<�Z7�X}{!��]G��fxY&TR�J�K>�G9���+Z�b\ۻhIC��� �,�R�)�S�����@�9�D ��R�a�!J]&�4�l�w*H=5pg���S3��h��D̗<T� ��ΞS��%�4�����
�$} �H�����d����)�l(O�Ċ,C\av�7�GϏ�v,��g��cP��>���"�!�M�7Ӻ��r@!�̳[/R=BB
��JO��{=l�>�C�ͩ��eC9�M�ϬF�ZicB��pT�ˡ����%�����o�%����[MM����a�A���l��F
hm��֠�h*r�4Q�I���F8�3TFF�1�|���W�P��鮕G��͊�L˝�D�V-��J�HIn��Ǵq-�J�����h�i��,����k��S0���@
��݃ƪ� �P��Y��U��1���ӼG$�1���,:��V�\>���BWr�g�F -�{K�M{_Q��.�:%��utP��p��G��9XG6DxEة-��Tk��xIrY�&�d�Qnڧ�|�٧n���|���N%�/ޠ�e=_�RnR������Y�����#q�͆�Y�_��_��Jt=���Hy�=�b�r��yv{-���w�i��[0)�7K���5B1�1���7ba��9�۲L�%��F5�AJA;�2<��^%%%<���w� ���'agi��9ڰ�e_~�?<���APT&�k��Ml:N�#_�+�脭3ğ�-��Z�cv>�?z�ȶ�ް�?p��fJ-���������T�\*N��Tݷz�U�m��J=r��]�-�Bg~��'H�,qR�Cg(���_=��������5������u�)�v��5o�4db���m�������ùx���J~\�U��!�-C�����+���'��䠩׫6�RV��T0��S�31�d� >����S�!����;;U_�E���C�>`��f�z�t/+٥W��&񵓹���-��%41#4�{Myi�`ڙ��ECS�漸p��;���IN����B�"��q��+e�a�����@��� �!g9��qQ�+Ԃ��<��pz>�L�z˕��7o�#���v{W�4����U�Y����\��#UD��g弟'a�U���9XrR<;��6~W�7�Mx��p�E��<�>-dTܺ8Nh�Ĳ��h�&�E���+sT�.`�g���K!�͢;p�(Dg��W���L:b/ĖG� `�W���#)�.-nk6=���Zj1�4��EN{E�s0·1�P�E��]�oSd��z@4Q(�Z"�ص���'Z}ĺMѓ�k��ſ��b�$qL�u+m��[*b�6��T�}�s\'�uF,��D�N$����Is��[��H�qS��i"	�h��m�G2R�oK#b��|�%��k{���x����yNz$mS.��3����ݮ��X����M��!I��I�F���K��lA,��X��K�4�w-传��Ԟ�C����2�}�Y��=b��Z|Z�J�[��@���LU�2�hyl_Uh.1y�Υ�:K@
r�8e~a!�
E��ǒ��P�` @�Tte.=�V�-7a}ҿ�\��ǒ�'�o\30��r��Hn|���C���I%�k��jN�V�G�����Uﳇ¬�{}��`��m������>�����A{�8=8;�!�z��݄��r�x'<m��&l���VI��U#p/�9X�▘� ߨe��}!`������b�l�8hL����1�f��(6rt�S͌f�+�i��^k��i_�b�7��]6�@��@ͧ��ӧ��l����;�������	�KI��iY۶����:���]?�.�v���oiyRG��S��NPw>��F3�B��#`>���
��b�4�@ �f��n^AT"1������3�n$j�4�#�~������N|�?�E�7-E�5�fG��4���=$����ܾ�6�54�'�˖kiݥM������l��ƅ���T���y�!^��7zc.�!�.�Z�-���.ʔJ�ST��jʅ3tl���R؎`��"������G ��=�ݲs�Q>�UA�U�Z̶�^��m�^<o�{�H��೉���l�����폎i��h�.49�O3r*0��m�v�k����\#2�W2و��b��/T)��v��Z�?s��v�X�X�1���G�÷biZY����}į���X,� -���q��jr�j<��ߩ9��ޝ[z��T�ݽ7��E��`�HM�
=A�b��rp�q�ω���>�Z茻*#h��p�XU'h��y;�2�t9��������Y���;��V��E0)s�[�����B��Ǿ/i�BOZ��3�%yAp��Ϊ+��p�;�׻��'H
��Hp�eg����G�g��$J�u�+��k�^K�˧]�l��~� qE�̢��5����װ~�ϟ��¸�C�%�FH�6�r'h�z��{m�JJwW�Tك��{n�O������i��46S b	-�;V{��!�nK"1ʱ8pL^�5�\�B��	�#|�h>�;�8 -/���9^+A_'IZ�߀SI'��ML�-׍���bZ�z�^Hp� �9�ɲd����Aߥ��~�Y(��6�T��N��`�^���#E��R!�Mn'7k�=(?�P1_{v39���o�&�,*[🗔��%�m��MCČ�F<������:�F,�*���"1�J!�=��l{b���0��09@���y�9�Ka�A���.�d��/T�f��� ��R�j�
M9>�ҝ��:w�ו_��`|"1ߵ�6w���8��sn��R��pӅ���4�۝���	�\>xg���f[x�L6�p��|ͧ4��A5�i��]ʹ�y4w�Im�y(��>�by��K���Z4 v`��(i��܏�ʆ*~P,IF_����wfe��S��jp����j����a��`���:��Ҿ����nd��M_��]M5�F���<p¡K�Y�M��Lyej�}�p8x�[���yl�{j%��l*��냤55���C��}7C�k~��\XѼ�6�6r��翞�h]g�se�n5d�� `<i�{��(���2,7��6������J"�Ώ FcKޙ�H��� Q�͒�T	0�Րa�~�wu�[JI��3�W=|F� k�I:TC��Am����γ ��f�끞�����><T�#��L���I=o����_�8#ڴ��ـ+GaU�x��2o��ґ��SqNn%��6Eu�\�G5�_-}�_Y��L������e��v����� �6� ` ̔b�;�+�A����U@\:z�@Gװ��q��r8^7��#y_zX�i$�W9�-�������T��K飒��m˕1��Hhu`$P�&[}ҪX����Y]�p��u��VoѼ���I`�-�ݮ��`	�����w�*��X~� b�n���K��f��RCHeg�%o p>E7����m�����$��V��bv��ݢ����]��}C���0��V+h�OYn2m� �_�1-W��&-�a<*;�2~����H�����ۑ0��\�5ǖ��y�ھ��.�嬶w+-�ۅ���r����L����*-DN)G�#��oВ�A#�����u��^�L����FB�ru]t��ww�nߎ��o��8�����6ޖ���!�nM�[�s#���*�D-<KML�s�P�4���~�;[�
�t��$����F؇=��؞���kԣ���o�҆��z�~O��C켟�]��o�$z&�Ǩ�}+"�Z����7,�,��4�ߗ��|k�V������>���΁��\ᾎْ�]��Mƙ#Щ��_۴w,v�"�(����l��Ӱ<�F&�����y/��/~�[�_� 󗴥/
��M�?=��Q��kt�5F̩����NE<��]�@����,#|��ȱ�fm^�K�U��%J���(V�?��y�ȩzmՎfG&��r��R}��ITt~�$"�bz$�$}��'+*<��e�i� l�{��L6xq(v�Y3�ش��;�|KC�e�㛪{ľ�\e\�_�ݣ�T/�@��[��3��>�/~��VA�����93k7Z�h��l�kx2}�ưkG�ĽGjg�9��`Y��uG�L��!FZ���֚��ޭy���z�e��f��Y\1(=��)ȃ��#a.V�r��>�$g�(��ة�� tzn�d���;?OgW>]J���jD���3���#~A�wD�u����W���E{S��e���[�y�N{��/��Z�q2�=2�� ǔ�:ܽR�Ihdb�ii�0�xE���	��mִ�.⸥0{���f���;([�)����������1��[*��1v.	�6�H��)�hg���9��}�N���^�`�������9�č?�ZːͽL�T��X��ϳ�}F�-
�ONo����r�dj�֙�LWgmJH^�	��|�m�����Q�������e7IZ�k�]և9HGiH��}=�b��-5��_��YP�	yC	�D��0�-���rI�ݲ u(*����S(J���͍����W�nf7��71��ٝ�)7s��ןp�gBhNNWծ��RБXK��}
U�C2�����VI��Ƚ_��|1�����Nv�*ŗT�a�:�'�
I��p��灕�<�"Ku�OL�E����� �-Ub��Сz���X$6�ml�EF���ޒ��j�2��������[O�flom���Zm;~5̛�d������?��6`��l�M�Y���%8��s\�:%Z���<#\�߇ޒ,���ڎuuZ��ߍ@wr�9����s^y?_��i��#��G��8NR��?J�L�v�,�b�Re�*_��a�M���5نr�����%W�B
hB���"5�D��C|n*��l:���BYSY8>�_T��i't�8����)0������>��e��A-���f0A���5g�z���h	Ks>$z�ey���f��+�ɮ����}"�d��B@b�9#cgA�39�{���Kͼ��L�s.a�9�Q!��������@GF�΂��2hn����<]�0w�'����&�-�	o���l��**�<��ⲡ����ZɁ��5l���t��H����/R�Kj�9.�/���Y�����2�p��>��
�8k���*'.n�~~�RU9�K��KO{0�6P
.p�R�Y��{�5[�l9Tc�8|H����}��G�_YRWy�ߙ�B �R��*B��|��Z?���vn��KU�r��2�Mvh�P��Ѷ�T��"I�߾[���x^����zȇ�ծ�5	��u�G���*�нy�n؋�H\���E�5��H "=���l�7� ����B��+I�f��8�.�$^��Qy��b.zW�O�};��d��'�P��܆E�i�E_?�� �+X˿��(>w>Z�E9�P�V�����(
��r������ ���0�!u8s-9��N��+]	Lg:{F�RT��va�s��&!0�_j��O�&�DDiZ��5u��u��=K�<̏��n��� +�ܼ�ڑU�?]��*Ds^5��:�r�j,�ibŵE��'m�.vn�~7u� �i?wL2��Er�/M������(�k�P�9�Gj���|rT�ms����`p�S�%�լ��?d��^|��d��fds��u��(�Цw��k����x�Nw��d��=u�2P&�
u�󡙴���W;�ş��J�}�&���Ѝ�c�V�z�-��\]��:���؈LT���}`o�"�����Q�+Q�ҫ�	ټ����q���N P�R���n�����(2$?^��ۛ���#� ��xs3^be�Ƒ�Lg}�Q�(���S�X�n9�\�vԨ\*T�j`���r�"/�~8�f�N�f"����LN��������=�d�����b��`*��d
"n��BaC����Ԗ�H�w&��t���<i��Z�Z
�(V�"�*�ퟘ�sBSRR�����6�%AG�s��%v��cv6����@o��^f���>��B�
��z0���\�� xtW06����n�]�u����pwpy�5?pJjB͖~<��d�i�4��?��1�{=cC�����wX u&W�ұ�q%|2��_�q��8�-EaZ~�O[���E��Ēs�x����v��ز���E�g�����X%+�euY2!ĂCW�~+Hl3���̯|ev���A8���ٯ�.�}=	�* [jH͆��2w�PrH�=��o٤�����ƱWCuC�������&~�+jٸ���H�TI�'�d-ͿTK)_W��)�WE}�:�Gb5G���W%H{�jK���0���k�{Q���+���	3y�cz�y���D8zV��Rn��Pn�ҧ\���K�j�+�R����&*&W�B^�ɒ�Qr�)䥁߂���W��_�Ħ��;���'�|OEE��{��nwJ�~�),�n�V/R��%���;���o�.��?{�p*���.��/��B?�u�̎�D\�_}�J�dU�����N��+��B��'@Q3)��5u�c��\�r��6o{hI3�PN�e2��>8�촳�s���
�/Y«�*|]]l�9t�Pܨ�'3�Њi7�F#���^�į�KKf��'�h@�$��yG6���VNP��}-Ԁ�n��\X�^����s�ph!"�2~�۝�d`�Fݎ�<kw�w���1# �p��M�O}1�GF�A�Q��VuϿ�/��+�)f�t/�����kӺ�������~_bWv�v�:�����^O�~�_m�_Ҳ"��!{�� f��-��mB	���5��|q����~��x��}%�Y?a��33����Y=ys��9�ސ4O�t�S�G%A_���U��� �@ʘ�ћZ�������������0�� 2����� ~1|Vh:��T�*M�Q�S�7��M����k���K̈KW�䪒.Kr���t���O����6����Yw����><�#V�	�J���<{ndj#�.א���q��jK`���Qt���n�7�T���3�[�E�
�X#�~�z[� �()M�@U-�����[�XUD�ER̂�!]r���w�l�Cݯ6o���
^�����ǈF70�"����P ��?{H����fn��N�d,���{0��ji�N�������$��BikW��|���C��4��]��.�����5C��{Y��)�0-*�M'џ�Itm���J8�݇�v����i�PRy���KW���B�V�u-�8:�`mf�f��_=6GI(J�bv�8��z?��׋[������C��Eo�IZ�����pͯb�e��Vf�_���HJ3������Uj�0��6~X�z
o��]Е7Q7R{Ɲ\��G@�D����]�{�^@f�/�o�k#�r9��cI|����E��oȯ�6�Lq����kҤ����\m�E�R9�@�j�͸$+Ѓ|cΊ�)�L{S���|��V%͚k����{+��Pw\6��6z/j�i���,vѼׇb�;�Gn�s%�c]�S���7�趖 �GD�	jNF���F�dO�N�g|wVN�~��|��H�
Ġ ���!N��l٨����� �s5U,�d+R��Q������A�X���2�f���o���l���`����hM����'p�e=z���\��k��k^�k�CA�A��+�^�{>���M����f�0%�uWK�ȿ�(�UR"x��N����DJM�
r0:SaU���:��a^�(�W`��_����/����A[�N	o��-|���~��P��moq�I:���4�|�/���w�J�s�z��tW/q�H~���_��2�`T��m`�fs�;�*&�tMÑ���Ĕ�I���
����_¯��A!���w�m�:�����ڿ�.Re�t����wD?Ɗ�.��ӳ��9� {���13��G�٘	������5��x�F�����T�"�M�,�i�O�o��y�9�����J;k��7~fT�5JGa�Ե��uB�߭�T��w��/�+�'Q>v������e?t!��U��Ok.۫��Ҩ��5J ՙ��>�<cp槜�"��z�n�)�1P�\��Ҁ����m�Gt��E��|M�{��*8����V�Bz܉�/pxH�d:��� M*��uD���8�̓��� N�ƆR�"N�L����;z�-i��ŔEI�{�N��l.H;�D<�\�}k/�hi�a�ۜ5_1���yw�N��h;Ţ�zܜ�
�xQ<�}l>x��^tK�[J9������a�lT�+�����.���'_��.�F��/s��Ϛ_�y��c��X��f��FD���)	�ŭH>�T/`o�y9ڗ!lfh�g�~@顯c��U�m�䫽�������*y�;&!	/�m��-l�rľ��:���_q���H_�r��Q�%k�Eާ	݇��D��������pQ2�;Ý�&��I0V[u���}(�L��޶�
�N�ɬژ�O%?˓�
mӒ�܌� +L�wg���|$z2�g�ø�$��J��.��&���p"�(^�^Ψ�Lf�Z�9\�����M�B�F& �\�=�"�X;�)��:�f��2�YB���ފ�4�m��V�D2S��.��7,!o�;}��������l
!�
s�:�?6�٭�/�;�5u��J�%��#�?��e�]�uH�$ecs�5ÅmFk��"-�����_x$B:���Z��6�.D0WE�Y�,M�M�H��4�+���g��c��NDMja�����8��(���ှX�����^(X8E5��D��v�*�?��{������t�s�~cqzg7��Gc�@���!���ʈ�N�@6K�	%f���{ۢ�i=�A/iZ��SA���0���>����K\X1rأd�[��0$��S=w+c�����䏥<�Op���_F�p}M-cf�˕���ϻS��r���F��Ү�z���;o�,+��.@�*��(QRP�=�3Y��`�\�hy�H����>��ԲZ�S?;W�D���MTk����rC����������Y�	�����8h!��mG+_"�,R��<T@�������鵹?A0J��|E���B�%��h)Ym/&��z�~�¼?d�Fz`g��%F�#�wg�E%�[$�(7׹
5�)�t�ɜ�O)�6}��T��e��*��E��ܽ�]N�Ubx�P�[j�y�g{��J�0+2�r���c;ع(�#�r#N�u[&ȡ�UzC)~d�	~��SL���\�_Ͳ�9���N7���i����T2�]w�bj[G/�/�'���E�������� 6�0���߽u�X����1�����H�Tʄ�vf�v�=���u��Jo
��~9n"�l��^^W���StoG���R�KU9K�PN��ʣM�+�FY_���yȞpi֝J�a �llX����
ꬅ!��R�ր���[�}ZTm���jؑU2$ǻ��[1@�=�K��� �n����Z��ї��)@w�����;��7��lȵ9)�V�,���h��Z�7����ߛ���	��������?�l;g�Z����3D���so{�2�1�ƈ^��o��+<���KOO���HsxdB�v�mrhЃ.�ͯ��lE;�9�J|�u�V
;��?�\��G������)B\,'�T	�{b���U��PR��_�u��X���:%e@7܃q�W��{+Py�R���O.z(a#q�o��l��a5raX�UxP륖xP"�)s���:��m�E0��gA�jg_��[I����o��iԔD��H/�DP���^�pK������|�d
˚�&���@��N+2Ōi�v��>gj��c�v�N|H�X���J�p��\��?�����!��d�4����}k1a�����r��X����ͦN���6(�n�Q����}�)�i����g���熐���ʌfu��wΖ�wȚg|;��}jbz���ڜ�.�O����Y1��7��c_A�,0Uͮ�f�h�E`\<��z<zo��qa�'����]��W{C�\|�K>�o��t��C@FO�l���^wAs�!U0?��:�*x�1����c�ڽ����!c��>K1�Ξ1=���oul���!D����� �fԣ9Pj٥{����8�0O�6�J���� 7[Q�C�v�&�������;)��T�j�<�"����V�6����w9�>��>WT��y��),�=��
J���
�%'_��Yw�).��y�q�6N�OS�8���!��rt3�/�\j�GKV����-vg.́�K��p�FC��e�&�'�<�t6K�G�v�0�[�9��������"�6�W������4-�T �J�G��Ά�6��>��e���/���vdٙh�)а�v��d��y�L�U��z4�q�_S:sK��\��É<��\��WWjc�����0=t]��x��e�VEi���0�q�c������y���F�����Ұʏ=M���Ģs���|c*�)o�rL�(����'�X㸿��?��g �D�CTm�J�4(�0 � H72��� -]ҍCKHݢ��1tw8t�C�}�s�_���j�{�[��t.�0���u�hc��\���CW�EJ��!!'��t��Cf�Zk���S���z���aZ�b����c�4��qA����8���/�G2�I]f"^�	�q�}EL�� E�f����W����T�Ӽi�	=�������,�S��/���=�'7�O���Q��*4W؉���ӊ�ʻ/�ء}S�o�n�\5]�*��f�-�F?�5
y��#^=���������	ŋ[��5SP)�F��1���7���<���T��ؤ�|jm����󂨁���f,��Z�_���>�l(�i��'Q9�p�i�嫠y�Vc({D�+�OA~nhQ��|qhR�^�P��˲eiTߚ����3Ґ����� /B��C{Re�:��vGUBޠ�}Ǿ���z��7a��>�(��WL��E���*$-
������=i7��u��[�]���^��ڣFU�1�u���kdς["g1��ϗ�;e�ή	�贒Q���p%�u�̥aP1}%a�6Cl1ðSr8�*�%��	�Ǥ��N.�M$�߿����l�.~�j|s|�U�m�<�s�o�^Kф<�;�'�LX)v���/�tٮK�F0Vx+���v�]s�dk��,��bm�i���R��������TS��P$i��{4�Y�X�}Tj0��m��|��Im^`sxS��]8Yg�鎯��>k�o�=~���8��k'i�ʷ�]��L��~��ޯ|L���a�+�"ȱ�:�ފ~��X���X��Rˏ"}�Z�h�0}{�v�I�ȃ��R�=Ks'R�����)LK{5��?�~J���?� JX�٧�G�����ړ&�<N4�,���,���9k��|�Oc�߬g�x������,���<ਅ�Ϧv�qF�!���������	&/��3���:&u���}|�\���3���R>���N�"�wV7^�Q��"K?�Z	~w^�;�{
Bd�$������s=<4�"'����@���P�n�&*�B�k��y�;JV�b�c��������
��ҌE����Py�A�W����w���+�}	p����	^_OX>+9j�w̻�܈�v�eH��t�q;�磅�S�O��M��
�qys�ss}��d3�o�]j�л3U� �Nї��xo��(U���g��}j)7n'�=>G���+**6��:��h%���{���I2�۔ٜ��-Vi[��<��p0�u�K-�X�Y��
�"�!F�O�叇Ȝ���uX�Zt��T!D�.t�4���-�p>��U�F<49Ibb��]T����*�9�_����?� ���[�F�y�ġ������(��N��s������ݜ0,uO,p�?��&qh��k�K|e�G�#r8���oL���Z�k��9���4��2��d�����Ԯ숚hmR����������(���o8���Դ��4�bj����~X�쇷��^��)�}m�����Ϫs�4;��:�2�.��*��3��}..�A�=0�}�}���]�?	ԏ�e�+����>F��	���y�BZ�kvh\@N?+Z���Sn)�V�-��ä�\t�Γ�M��|Hy�}+s�5�g=/=)G�`�<�s㷌��`,����3�g�!����n���>6v��]~��;:�c~p�'�ebv�>�(M�c�2�b���~�A.s�5��z#r�l�`a}�ZK�|�Z��G5w-#��K���Q�����>��>/��j{����O����&����e����Eh�Q;�I\*��שR�qq�,�6j���0���6�!W�p[�����P�.�2E$�Vr?ٗ�åv�fL;�>;���R����Ȝ�ƆJ5���Ƞܛ�؃�p��ʛ�4�X*����@��::����C����k�؞ާ���]��*AG� g�<"�F�_{��r�|���HJ+��a�߭�=*^�����C�t�ܯ���9��_�d��V�[�Dt��!P���b�+��}��ϼW�I����ZsYg=g�]+�Kh�N�S���n��}��$��b��_Ln�2���9�Py��T�L�-���\�gu��N�ο����rr��ި.�G�9����o��{�r`@��4:e)I*3�����+EѸ�dw}ï��p�-��l�w�6��&:�r7F���4�ִb�g�:GrJ^��)�5�1��
��2yVD����=���e7)a]F�`SD9`��L�Js�dW��N�����9Ɏ*p}�a�����!8ي��������*��{�k�K�B7���`�諍����)�ic� �݃gm����z<[snq�54����/I�_��ˑ?�>N�}8:���]���uK������َ�u;a\�2N��Gdx���O���ʂ��>┚�+���D�G��ז��� ���|'�����g"��Dzc�g]�e��L�nK׹od�*��T�|<�kҩk+า i|�f��8�i�-H��=��2����E�U�#�*�FH֨�ɣ4��b���}�ӏ�������|�U]�fSC�c�+v���c9�@��>T_�1v�:<���,D���ƔG��z�ʆ���=aP��Y�l�le�
o$���>�N�N?�N~p��*O|�@�@��_�����=124��Z@}�p��R���_C�g��M���OJ���E�5�>�O���Ƙ3)���VvM����<���7��DE�v}ڵ�i�$m�C��RG�4�R�����*�u���/���PY�:��"_�Y������?���-�[!:^�f�����ArH@ ��l@�g�X��U$
viA�/Lm+L�S>u$�W3ֿ&�Y�otf� ];�]�����_Qnx~����;�ո����I�ܜ�Z�p���w�y��wp��|�pI%E0��\o+?)_�gZ��w$�0Ɂ*��z�������z��N�'� ��8���~�/���Pd��G�i�d��$6�]Yul�����f�j��v}nӴ*�, fuKP�i���4�W�w�����2v��[��A�B���w��2�".x�B�Lݹ�>�jiC��ࡸw��~�ˢY��̝.��C�eY�����ZS,������'*�Ƀ�`�;�Ư�IB
��8��34��w�M�>Ф����ٵ;�\�u������+��C�Q �|�oe��Ðy&��#_�����4��R��ݑ^+sW,�$��W�K��&��/x\L��찂\�̍-քX$�����L��F�ꐊQ3DW����/��{>2� ?���_q�N�G��U�NA�$��a��}e�ri�o�3���g�I<��&\��ëY�?Guj�(�4�����w&���z;7U�DlT��a���Be���mk)��׋;R�N./	�t������X��hNg?�a7�9M�g-RTf�?�����V��l�>��ĵ�Tҗ�)�6EǛ�6�'!(�)RyϠ�̚��?�� �	1�s$��ir�
~|t	�e4���
��c�	�&�l&�D���*	BV��4�x>.�]�8��p��4�!YW�l��3�L���E��,��;�Kb]�g��,�#���ـ��h#=Z��rSԦk�輁�n��['[Bƭ����sDf�ܫ�G(���7��W.��sf��&��e��~�*#n���uD&g�'����!U�4ý}w9���ڨ�v��b�쥫�m����`��a��:m��l�Iѝ��lR��Zī��,߼e3�w1��jmK���$c�!�sV�7�_FIcʘ��l�~�$��	E<�`C}�;�Έ������.�R�/���"��r� ���m�oJ�Zl$�+���[f�x�>QJ��?��<l/.�<����:� 3S7:�>�`�(�5�d�Tx�a���UZ��w"�����x��(3e����ەdbT/Qԇ������v��i~��&˹�~��m�Hϸ������D����J��T������2���T9r��[ʪV����8Ȳ���v��&������Z��2hO���Zm�*,,}��{%s���������.`�,���y��@�ʮ+l�~�5�x��Ĩ��E�fE�2�D���g��[���9R�gN�8�j�
�D�������^�Ã�}T��΀�#���ؽ1����Ƚx����q�Oޓ��,���n�
,���Ŭ{<�}����r�+w�ێ�m�(��4Ɏ�$h��(��Q�'�t��Ö�yQ:W��~q+�P���O�����֞��L�'�+:�Ώ���f�
W����j�^����x��LFM�URqZ�i2IG�{Z��|��<f�6����[�}d	q�,g�> �C�h�$�@��RH�}�%�=V�p��9�j�&���A~타�|D)F��D_�#�Q��7��5����;Ij�s���ēu��U��T=����T����� V��b#�+Iki/'O)��/�^�s�b{7����� �͖mE�1�N������w�_�)��k��V 7��}�$�܀�q\��Wo��U 4�HZُ_ue�;W�,ԋD��_�к���jϜmO���]n�{�3�������,���n;�mÛ�#8�R_�$�v�soF6%(h����6
��7�n��lb6� ����a�
+���,�;c��;2����ˈ	hԟ��*F@��&�,���90N9�+���_�=#
/�ؒ��%G*@xh$K��٠|�4�+Ƹ����K��}�� �L�F��K��f6�VPD�v�nջ�p��e9�15���Mqv>x_c7�s��j�"��(����J����Btѳh��.z�x5vW|���;s�DT��b�3��/�2Pf��HK���g�Ҙ2I$y>L�r��~����C,���YL��r��)ݚ���+�AY�X,��2�[�g�g�C�@���l6ߎR�OB���{��QO����M��{�/f..>>�ƙ�
�2�5	�V2�J�d������<�����dZ$J����,�`y��l2�޴��\a$b�&� :k`�ި��~<����b���F��}>��/�����~�
	��'�LS���n�˗�$e��JM	��9�z�/��c2���>���
�I3���ǉ?LrԦ�1�<�z� 򆳇��&B����JMq[f�zl��	��u���q\?'�� D6�m�q���A���|��x����Ww��-A�D��3l��>�=�[�@�� �vXX�??`iA6[z��\,�p��B�YX��֣�ny	L�}�R��U�O̻���X����a���Q��tw��5�}�K��yx�:�g�*e���/�f��6��2_49��/t��R�6*�f�1/�v�}�Qԋq�?����o�"4~x5�Yg(�dF@YA�K]���?�*�������	rZ��ֳ-��;v��:}9�m��R�jշJQ�C���mݬ�܌5�l�h���V��Y�����+d7!�+�ytcg٥�ɥ$��㵅{���f�����
D�Yk�/�S��S� ��Y:|h�|X�K�5_�M�h!���0�I���Eޮf��� ]�q;�u��c��FGŪi��l:���~�����]�]�s�=���(#n��Q��")A��(5$�JPm��(B����fg�i���"���/9X��<ရ\?Ⲋ��/��ǋsӇ�ph����$v�[SG�O�̅j��l���u��J,�^�L�6�� =���c��Rߑ[p��z|��߻�|��~K${�g�?�:��l����h�H�y )~��Uj.nǥO&jqꉔ�j�#z
g1.O����<�I�o�������J��>��]�%k��AW뀀%֦G�'Qgw�S{�����q+������<41\��Nn�BW�[^&�X�pG�Q|**|�lk�ҶB�nq�R�=/,��qGM�RO�CK��8���L��7��&���lt6��ζ}������w�����Dz�\cҟ?��g��vߘ��޺��:U�cP��:�"��r��~t�H%�P�.�|VOK�bJ3�-��EN/��L�T����,�qo�0d���b��-F���;�"�����ӳ�0��7�I4���b�U�Յ�%V���-=�:�/Q��x2�,!5��d�/1Sqd�D���z��dPN�6�/	'�d�bg;�OUTRxk��d�ñ4�ݷ�A�R�22��� '7]��?R�}q��`�|�H&"il�[�k������B
��h����B��Y�l�p'�CZ1�Nn���7��w���d͟M��A�����,����'ߌ��6�`|�h�^n�d�ǻ߾��^CdZ;R�f(�q�Oha�̓��M)<�4�v`vC�g-ֻ}��ﻓ�b���QJ'H�GC���(�\��	�G��$h;���]��X�G�W��*'l�_ [m�Z�D��h���4J���PK� ~3R�
tV���6O󌾶���j���CZ��y#�7/�r�)��p 7���[�yEB������e]+{Q������|OJ&�B ��٫W��<�~�L�]�l�0�uq7?�S�S0��2.�z���O؂��aaԐ�H'8c��������ޑ�&*nLΦ�g�OZ��^���J,�S+g:t����H�'u5,��'w舷P�cD4\ݼ]�S5�ҐSz��;���1kF��s��/L`�� ��ݪ<�-�G%h���=u����;�%�������+���7���7z��S�|�~V>aƾ:P}E�J�ə-1�I�z�=�*S����`����3����*P$�D9�\~���ܜge{�������"��xI)'���3��}`v��V����mU�����,Z��hWJ6��)T)�<�N���4��b�"�,E- ��;�d!C1�������y
�"!�����)���&��7�S�� �(�J��\��*�?<PS�>.O�;Y�#&Jv#n�VX�lw��?�,�x�/�k0��|>x�3O��X	M�y����Qm��a<I��mZ#2�ngw���=���?ٲ��	�=�O@ȢH�hv5��`�q~�\]]���u�^&�"""bze[��!�Z��T��X[z'\���~���ׯ��=�u- ���Y��_���lDٻ���p��2|������'�(y� QP)��^+�g������&���o��8�ǾD�c�{$[>�/�j�Yh2n���̠@BY�s��TZ�m���' �<%οW(�>������#t��p�sɿ/�m���-\)CΎ�B��:��x��E�f)g�+ƳN�P;������Lt�2�31��e}?1�����Y@B�S��;Ap�@�;&���1��g�=aL���[���F"sx�?[p�1*�7H�H�$�PF1c�II��KW�n8z@��"9� ��^DQ�?�	�i�%tk�lte�Ir�ݢHaO=F�ac���{ɟ�VPQ�0T��"��Ճ&wd�cu�X$��Im��ΉS�n���q8��1@����Zi�wG^:έ���$<y<������"�P3�_�]�Rd]�U�I)w�|]�Q���lB�6��I���|�Ģt���a�.i�o)��w�p�Y�Q����SL~�<�#Lh!���s�0̦r�De{;�@�6d-�5Zya��Ӯ���:]#v	�;E}L�X��)Қˆ0��%�Q�)��~�GC�������%gM�5E�[�}
��W�S>�{�1ո+nx��i��>�K�
�J������.~���g����-/����Ơ0�_3��U�]�l<�?Z)�j򁻋qT�V����1�A��5��i���v�w0N[����R��x6�x/@"�/��6�M>�3�|��*���My�V��*%�4$�g;���^��Ӹj_E�V��			�� (�C-<�0�#5��X�V�X�^�����q�{8L[<�N����W�^�(�6�<��9��6�H�o��a���w$��M�=�y��Ag��v4�Z�]�x��s��bT\p���[�=s�$���O'G1�)TN�tZ�m��U1�z�4ǒ�\��v��]���[��mCA�����("�m��(��"Z�;�.��{|�.\n����CW�;�j@��#ֻH|�����N�<�o������Z����\L�w2�����gP�M?�[l����>]X��Ƿ��t�P��:��y�\���v~�f�vb9F3�c�sP>F�<�ٯ{�9��OB��.ͯ<#Ge��GK��U�6o�X�?g�dV=��Q�߻OEɗ���h�Ѣ��:�C;	2Ol��F���.JJ�q�n�7I%�h��1c��iGU����m_��Hʜ�wC���O��뾁G鿾���5�����i݁�p�ڠ��H�zEg�W�[��\t�bcB'n*{��^x�*V���p~�g=D.�h�·%'s��n��}SS�nl����!�m�6�9��8Rz�4����I	c䥠��h�����[�KU��0��.A��4"ZFX��>�CW��6�(`Wh�v'�"WL��XH����~���M�<�'�z�<��L';C���^�����qz��Ҟ;����e<���S�xv�b�8�K�e%U��B.^��iy)wr��I�iў��da����O1�N6#G�����N����u'�ؕ�Q�?�I��l�%�v73Kcҏ�����~jX�&_дk�?�_] ��W0�m��K-T�Ë���
dE:���,��*�1�t����Q�^j��|�_����D6���o�agwq���RQ�ź��X��n�ezm�.�C�1p5���<���5}��pJԠ!��T˛=ش��
���K��Fbsr�*�Ì )�n�
�\c-���A�֨�$���'����@tUp��2*ȏS�m��BT�}`��(b��xAs�;(��;��uk���O���%kԿV�I��w�*���I���]M���L��3M�k����)���=�0� ?�(�C�U��I����ֶ���;}z
�P�V�˳*��6)��5	2�W2�P�ݔ�2��7�&��������YOt�Ms9��C�H�7'm��!�Q�����������Hh��g���L�(u���YG�b����;Ȫ�,Ɗ�i���ס9�a����D3�4���^5i��ަ.�L��@���_Y���i+g���U��_��J/��}B~���֊�@� �g�J����U���Un*��¸\5��p�lH��w*jsq�!�8FDU�D#��ʶ�B�-,���bI�'��X�#��s2�IC�|����Z���&��%f�܌?"~a0����'!.��J�(�����]Zv���ȇ��ts����k}~�ÇF�5�W�$��G�}�/w�ҊZX�Mw��P���o6��{�Tq���Ӧ����ܮ����3�"@���N��]\毾�2*TGR����f(!y��;P5G<:Cƙ�K�$�A�?*CnҲ�ԭ�;+�'��]������β�bS��.�\�|��<�l@G�o�T �	X9)�Hߏ�Χv��O���r>'�Aְ�i��cp7+�������&"�`0����*?��;��X���~R�U�I�~&�.������!ߤ
�^6�����Oy��/��'o>!.�-�D�9�һ�����8���4�	.Տ/����g��{����G���Ҷ>�ӔN��ׯ�+��9EYRqS`L�El�?hkZ�t�p5�Z���$-���Dq�ݛ(eX[� �YfX�vFg��q�f���X��	��aawqE���'�+��P�nT�k�8p(�/z-��e��oyU����W	\�����9b�P2bus�R|� �}�˄>͌��p���G�\�2N�c���/8��9[Fq$K��XZ7U�-Х�3�L�Y�0"cx6d'��j�̞���u�<^��>�*���@*
�~�׺XB�R?M�腡�S~;��RhO娂?B�blo��%%��t�~����餕��i��S�"�	�]v.��"�w��^�Gs4�	��~5Ճmë��C�uy�� �����?k);e�������)c������(\���TZ�K5�����W~���&��N��8���q���W-O�)�^V/���3A;�M��5��#,z��*�?E^��,�N��) ��[A�4P��f�(Ai��䯅��P<_�Rhb�R��j����+�ߙ�׸ڍ�<b�\����U�����y��I��[~Lr�����Q*V��N�g ��3ݹTS��{��O~�P����OQI���p:��K�i�I���ic�b��4���q��5�:��:|p�v�����@�Z="��5�&�3`�!�<"X��]J������$ (�"=�w_��(�#&yu� ����h�Y-~c�\����^b�q	�R=!J����p���ջ�T�%�v_� ��7^���7��{F������Ld�`�o`��kl��p2%��vLE�9Z�A����LFDG¦�>���mq�{#s)i�DP9+��d�����G�l���i�2���&`�
��Cư��m����'��G!��֏^�L��|���R�J�<}XY�^�j�1�¤g0����X���ϋr�����ҡ���Zjy5�t"��.�r`P�15|!���9�𻆙FF}@t��V��^z{��fW�ۜbKD�O��,�߇��K���;�y��u�-�k�����D`'<�%@���.e]xz}��f`9g��2:W��Oc��s�]\'������Y/Tv5��o.!��F��ܤ(!-q��ܳ\����%ꛊ��p��̫�h[�/�uMi���v�5L��Ŷ�l�=� ���;d�G*�$5�}�[�픨��^�9a���	��y�n06�O��5�����bN����*�^
zrY�Q.�,�ۘbQn��
P��b�\��4A�2/�%�J�.��^S��Mvj$�zS�M*�B��fՌ\A-=�9��K�W^B#7F�~���[G��� ��^�����̓v'���>�6J�|���Bsu�_����XQ�❍��!*�^������2�B|�$"R����FM����~u%W�g4G2��,/����:�8yu��ۊΚ���IyA�^��u�$�U=�Z�ɩj���S�B��(d2��
sD��R�e���A=��[8䢙�5py��k�t�9!G�H��9V�nʀ+���<���\r{�c�'i�	�50�j�Lx��ԋ�$|>#�T����+
�����~�Dx�L�B���1*zb>���(������^���~Z��D��������(:�~�Cn���$}�=iXg�WF	1�T�Ű6��"v�~fo�6z_�'XY$�S���,���ʾ�1�D��i4�����yD��J�ly�4��%�-U�p�����+�[���p�����d�$Pn�[���PLŐ��_���`םN�,V��#�3�Rw����L�!^�<u�)�/�h�Oo<��`ųR(�ӡ`��8��F�_�O�w�o9�!ׯ��� 9��lP�������T>����4�۶��.p�O�tZ�]��s��dOGP�c���g(�����35�V��>x��K����ǰu9�����0���%l���K� H!���TP��p���:�]v� 8��$
� �!�����g׀�� �0�@�zg����Ǟ@�)����z��14�ґV�S��>�VV�+'����?#[Zp(��V������=��I 6�TثF��T!Y����"�9�L�f'yhnVN����p��m��7��lx��1u�/�ьe\�̾��ǆ�:�p��l�����1���iV�p��h$�Z��T�B4��=�.^�Q���R��n	���FKw���yU�J[W���1j��Ž�e`3V����'���)(��^��i����r��9XMMM��o	����(�"��/��$GL�+��Q�6���jj�7g0i��m͡!�^x!/[{Y��/L��(|V�N�}�'�FLR#zP=�D4�����V�o�Fv&a!��St��89Y銯YM�*--�v����*�Q�._L�!F�+`-�e�C\1����J[f�j(��̺o�,ԩ���NP��N,�����քq�E�1Ο��?	�SƻYr���/N��í�/*".��8lC"����7#W��q�4�!e�K���1���+X�'o�CQ4G�E�SN%/|}���-�)��_��&�s��e����O�� {n��1xC*-�CS�ͻ⢊��;s`�$�G>
ӏ��.N;�sP�V<-R����b҇��$�=��V={�0��d;�f_:9�3�$u9m̓�B�ܤm����_P�n�-��_��~e�ovʨ��U�(�C7��U�ߚ[��/�|t�`#ds��H�h��t�C�%�nD!68�CV"��m�C�KJ,���J���S��l�*9��SC��7C�nR�⴪�٤��u �>�/¸�۟�/OD� �ߨ�I���ͷ�Z�j�=��� �Թ-䬷B����7��Q�`{_��w��\���^��@p&��p���e����������I�x���-�@��x/ہK�㖃T���~1��)J���?���;�<�amd�:�5�@�\�T)��jU?u��8��� .�#�y��}�O���{RULAW�����
k�%H�����d�8k�������W
�ŝx�F�k�8Ĺ`�S��&�F��*�ɐ*��_�E�r�W���-#@[M�N�-� ���B��;6]"  �y�՚��F_z���Ig�������u	�������vR�Gj
�c�9�`��k�	���LY���r,D���Ku�ֳ(�Iı�0 ���y����r�͟'���bX�w~��t�-�~�T3�h<X����P���f³�� |� ��E9�C�dk�\թ�����a\7�6JgѱJ��سȤ��D�c\�_����<bM��kT�,�?\����Z��W�J� ^�p�JaP�5����+��3.��'��Z2?�<k�p�����b�f	��j�:k����?�~�6��Ȉ��/����G�F	�Y[�'�э�t���)X� �)��_O�����wM�����L {m�g�r�)M���sa�jKk�T�HE�%��׾��ݝn#Pn#���*��bZK/���G�s7;��X��	����G 3��W�'�����;]+����諔ߍ��X�f��4p���l��*�Nx�S,FSkt�+��C����/���|L��1급"wKv+4�KYͽi���>���ve�p>�X��:,��S2�V����D<���B&O���e�䃃��\��Ӫ`���6�n��$��v��v�Ϟ�;}�a�$m������������K�����.�~��Z�N�F�v��棊��F�����L`g4�ۑ�
s)�Z�%�2QY,e��j4�IkJ��o+_!B��%�G[�� m̳��h�������	�b^�8Kkي����<\����a�3��3O7��FN�/�1W������>�c�<��{���z�����q��G���~��%ʰ��|�21"ɉ����s��d趨:q��P���dw/^�D(��n��g�o,V7��W�\�]R��5f���6%�D&�^�!V�;8C�r�r�?Jy뱉B�F^�ie�'��غ����SL�y��jp��öao/w.�՘����*0�4ǧO�y�<M<ߦ��R�o���~��@3��Ւ(a��R,9�gB4�n��yU�q�h:w�gh��I@���R�~I��q�o[��%�rP�s�@���v�G�M����eۖ��-I\P�j��l�W�+oC����(�HYu錳��A,��0��E	<�/&g�t�7����]$=�bsnwiXֿ��������a����e�az��>Z�AA�J+�m&�cY�z�Ғ!1� ��\_@���^h�Ĵd�Q]3O]6r�G���:6
ߘ^1,jH�	�p���y�m(i ��w��P��;LA�7J�bm�����;����V����E��xBn~^��<T�ߺս4�p�x����Sݜ��Mqq}��x��I�����{����� ��5�|���ɭ�/Ռv�s7�s�U�)���+x�h�}"��X����9��ө�~�ڢ�jkH���;���M�	#��G5(�4Z�p�&�w5z�p`3����n�m[��x_�~�9O�V[J+�����cZ6�]V.ʘ}[u�3��2/}O�B�Ot6��cv<���GA�|�$6`ύ�r˻�k0�6�h��,C��K�7�ٻ���ؤ/�a�k_�cg�(_����3���j;�l�z����4%�4'y�F����L�I��_,��O� �:B��uh�xǌ�a�ܠN��|6����]�ݩv��S��G�n$r#�r�;�2��m���:�JKO���d��ݞF$�o'}��$1(Y����^��%�o�y��?ŉ��ߗnV�	��bE�;:S50Uxj�7-�Lh"�~F�ױU��[d����h]���G�����c��`��0�8��ײBv���J)�QvV_9\9v��ʗ�A��/��~'�*�*��G�aW�P�@j"�/#�"�{���]�������I��}M,�@ڢM��X�7oHUzw!C�pV�UJ
"�
�*'N����k� r��i3���%��n�L�c�%}��-�6���?tnO��Oh����m�O&ـ�v��$K�hZ&��z�pEO8X=��ޡ�GM�b�Hg��X���OZK�r �j�Ҙ�4^�kQg�A��x{|�z�9Z�������	G��m5Qw�B�$�<�L~�zA;�.�?��8�N�//88������w#�b�z���:/�v[��A^`�;�6uo�&���#tԠd�x�����Da���!���®_1mY�Ɂ4�͆s�1ڪ��S�/hB�=�6N�:S7��j'��RXX��D�{���J�eX�"����x)[l��Xv0�$*��o���8.j[]�ш=�����C�jW�j�(Bղޢ'��$�;T��+�z�1��$��h���F�ڛk����;�;��kK,`���"X|Kdp|A��Co�\��姚%�{q�ۧ��I_�f�2j�6W@��'ؖ������xE��6b�̘�G�]�)���D6���1N<\�U$9[��Tks�i�F���7����ģ����q�|��)����0��mÁ28V�Br�e-��Q ;����|@IP*z�>qM�N����O"�OSg)PR�;�5������"]b��I.d�����KR ��ab��1��ܩ/>�����j���S�lXTZ**v��c�C���|�z��pΥQIKt���Fy^�0�߲Qc�fT��},c�R������a�놇��T1�
��_Ъ���$"X�Na�p������Ru�9�K9mG�^oJ�u}>��v~^���4������K.�	y����a����B^7wi]*Pl�L�>�٪�.�D&t 6MG9�#������uG~6T��=��k'�T����o=���oC1�k��N�TC<{mfÄjrK�C��>�:o�"��mVQ���Z����*�]��rd�Z���\j,�csLZ�x{&�Z���p�:��xP�h�ݻ�uQ1�fGX�Q �x'o�
Q���L��S�5�d�#�GN����j)s�Z
~m�y�̖�����t�0�;ZQS���b��>��x�z�*-|��R�h1K�-I�Y���H�j>�*��/�SHk?@��r�F�g�	�W�Ge�#�lq8�- 2&�z��bR�0 ^j�(�*���2�]�\�����`c��
�|�Z�(ұgS�Q���h��pn��_��6 `���e��	<��ɒH'݊ŋNx�R�u��/k�;z�G���r��]9�G��?*��	L1	�8E��_�C�C����<�i?���fK'�o���?"���9���/XA��3�-,�HO>�̘�㌂P��#�um�e	��
Q���>�}��߶*��0~3����:�҅�׏\z�˼�`����M{�\�7�`X�G
+��p���a�;fp�!FPC$���WSH��>S���Ɛ���>�J@��_�6 ��UQ�m3���LK �*d�����ו+�@�U�l'HH.�s��̔M</+�OZ�,���6Y�}T`b�`������6�g7���AOfcå�&~���#�b�'^��������濝����5q�j���?M%�ھ5{`��FBAٰ���-�{j�R�����=��3;�"`nZ���K �밑v^ǟ����	�k�vVӑFgdӢ��Y5ݯ��$��$��q)�y�m��,.X<є�.�M���������k��	�M�qi_�:ۜ������s��Ś�(��(�@�3�OP�ET���c)��#��>�1�/n����*�?�,>���R��XJ�~?���0��qM�q�I�p4H�42RAAA��Q�0R�A�AJJ���9R�F�����y^�����s���_{a���i[K�0��B��P���Z�,��@M�s���5	_��cXǌ��j��o{�{� ��x�-'�s]�sv6�/]���ܸ���&�)��䌟l�bkРt̖b�t�G�X�
�50�4��k ~��$�6J���/g�I��3�����=c�Z������l3������]͇JQ@��I����%�ά:�~*L����U�"���A�F�8�W����*�K;?,�ˊ�%����R�ݏ�ؗ3~U�t�+�Y���}q���X]c��YdB�*-0�֢	���: j,{W+�S[�?��uM�C���`�Wo�(Ұ�I��`V7s���x�q;�WVJ�Ў����F'���7!8~g�u��!$��*��RLTA�c����ߣ�]^Ɣ�l?i���isp>d�Q_�_�0�C�wO2����$��3�Z�o��C�*:�Uͣ!�p�D'���t���5����M�7�j���Ab�'C�z�b���6�6k��g�U���NO�a�����*ς�ϒ���PR/���o����6�n�h���Qj�%/�8���l �6I�ԏ�W����#�|cG�7���g���_�)�CYg%Y��i3�jȍ�s�N��3�����J%	���u��B�.Fj���(���
������|�yM��غ=i^�6���@��T&��9 �jZe����"���g)�Oc���¿��tF8U��V_�c��0��y��5��g�F_��7`Et�׶��I���1��G�Agx�-��g�zZ���	��P�k3��玷V����Ϸ��x��!�,��S�c�Ƭ�R��(���Sp���H`*�>�qږ���&aEH�8�+��H�%�JYg�Ivu��L\���y(�o-����<{�$�-���1�&/�$|	(5��޹��s��ɺ�j39cā�M�g��ś:�:Ҳc�F���*1'��^M��=E��E���q��`�*���#��Z#�,o�_S����)q���K�]%�U�Ok�5)7|;:�Ď*PZ�B�V���2߲\�c�����uL�A��#|F�ό%�؟�K8���)Cm�^Z�R[*@��z])���n���}-�>y�!;��ĳ�}7�f;����w��4�PK)&��5����*~K��JmM�2.�$�>.�}��\[΄��&7	�a5��{F�Dc���²D~�1�C!�࿔� h$o�L�T����%�p������0�ܚ��:�:}u�!�n���L�
��/-��xIo��'�6+^5N��b�{���UL�h�(���,�QB&P�T.?�0kC҆�d���EzH�oM�5���~]##S�����x��pۓ/�	��7ٜڜ���Nm��/yB�M������r�2Z}W�,TJ�u�©�D�f���K�$i�+�m���?EUO��ĭ��}j�i�*�g7��݅�|����x�5�՗qR�\g]6[�29O݅�v�<���>�ߕ���M���k�Z虁�2�s�|,5t�w�)o�T�T*r�mG
n��۾��A� �>�}�MF��
b���q��v�R�y�G���8����zN��jP�aa:��<�]�K�5wB���A=)4�'�%�WN]��׌ct	I	Λ;]�j$TT{�Ӗ�e�H��[b�"Z��lu2��yNmկ���0��9r��Rp@]��ll��s�����Cm�1R����1&�HbwK?�í��W�Y��p�Y��$���T ���hۦmm�V�8E2���)�q��3#���~xk`{b��r���P�ۼW٨�HL�3}��rR��m6&Kbl���0�թ�p��wֹ��y��߲��F�ͻV�x���7�����
�5*��]@�SR����8=�4�}�$���3���l����*o�sx��Yź�LV����R-�K�=�Pk��^�UC��\R#�=��$�_���q��Y'M:���%�g��|����O۠�����%��I;_��vЖ&�S`$X�1;�W�`�L�?����l���K��zh��S�)'�ck����dKo���kG龥�B��a���4��e�*�\b��0��EN^��/r�IZ�-q6�i����ȼ	c\�=w0��N��q��G8% �}8~��-�g�a�
sˍ���J�(���3u���.:W.�|�Â��d<tMa�gTx��N3L��ǝE��	����I��MŸL������b�l����5����뺗���^�3�S�^�-a�(��Aa;Q�r[�
���)�˚�����a_��	�i��Ӝ(��+��A��J0g�`��X�h��6�[+
���O����"��G,j�*e��L7q�UR�E�HI��5���&�)��QzZ��l�Mq���|�sK��_��4�)"���$9��u�Au��
'�;�rܠfj��Gr�?����]��U}�]�*� ��l磈���\��ҿY�?��P��/ͺc�+���+Xf b�l_�P\J�O�U�e�UӴ�x��c*�7��)W� ����tO��,�� ��MY���#���i�+��++dm�����ѽ������Z��a=#^%i�j��g)��v����,|5���0����V(��p�7l	�6�Z޿�x߀�E��ƿ��*�C�o�q9�R��`�'�����+���x�ka���[WvN���3y�Lޛo*4A~E�s��q�g���*Rk*��C�`X����*?kd	������s{w�'��+�ӍC�TH��+U��\��s���*��A��p_�1��㬽����SU�-r銍g`D��ՙ��p�Tx�3��0e��[�����R�|V��%��ƍQ)���<�Q�:'�/�8��MEnKG�j5���A�(2Lh�4Y�X|�.)[?�ߟ	�,̌Q�N���u��@%h�H��5!|�e7q8\
��-;�%���ޔo�������]G� ��;���Om���QI(����c��a���GRUK�z�1L���_��L��M%�[�މ�O�3��}����d!L�p���6��/\�%塙L%�ڣ�i6��L���E��[�,?��8v/�R��=ݔ4��_�jd'6a����_�iT',''�5��5^8ED�#�t��"��9�u�]�^GUUL�}gO��&�N� 7;92��?�Z~0,mv5��72_�e?�Y�.BE�E�p\�]���iX��->���:S��fM�`}"%{PoOk~��e�U`u�ű=2=�U*P9`W�ct�z<��"}�i*Z�N�����\����由n��5�7y-���!��3��
i'oɬn=�΄7z�R���6��!�&?�lzMد�F=qie�ntɿ�2E?I��y����69̼�I/���ȝfMh���`�J�g�+��"ȳ�o@����i�?u����]T+���"��s�̐M�:!<1#�'.�s��C� �v��k����ѴE������֚� kڗ�7q7�X�����J�,��TL:lU� w*7%'+�集ć@��%9kgx-IJ��w;;�TZ��CnͼZ{��`������Ak�5^t�����R�����W��aW�06��3�φV	+���T�YC���J�,&;��|&�Jh��oĵ����äȤ�6��W�1
6��z����6�D8׻���~�7�Pr��$����<�L5�Z�M�k��>��cZo���*�J��;S��-����߉x��\����&�>��-��b?9~?՛|�������r5����� v��Z�s�q��˼X�P�?N�a�3����d\��A�+�̡���� y)
'�͒0&��O�LP��9� }��Cb�U�$�C�J
�r6��4�����7Y���,�u�^<�'�n-\����������O�HD^�&������@Uo�查���`�i,��e�Bj���g�tfmZ�f:��}!zbiG�_{^��V�أDĿ�:ZW��ӫ�'}��1����m��kx{W?Ȯb��03���sRs[�M���"�(�Ǻ�O���0-
���w�2��j�j_G J�����*P��Ҧ�}�NN�׻�'�1h͔��?��6��ӯ3�g��a���:���r���dra�J�
"ll�߫�>7�0��6�ɮ��GCKk �"����s��IO�)�9Qf�7e$yQ��x�<�3G��R��-h�C6UZ?q�y���~J���쐓(�1��z��㪧\N��h���Vb�(���e�$2�=�5Cˠ� �l�����j���b����a-^3f6Q�|�/�=�
n�n[>#�����:ӺW�'�q�;*E��f;�����Hmj�[�.3� B�ŝ�&9e���]К�D_��(��t�!� �A�o���۽c�b$�~����f��N�/�X��~r�=*0SF�����l~V�щm�inpoָɐ��T�9�q��3��>>����c�;$��	��\!���fFƁls�J�Z�& 8�P�ڗ������5l��~t�-��T����\�Wzd�R���RN�n&���%��U�W�wt�#&�D1!>�?��8=M���GN��nWh�K��b�Ơya{%�%z*v�K�M�8� z��U���L/�?����N=i(�OZ}�b!����`���<L?��О���լ;�L�!\J��/P�V�����ظ6�x�Q��D�ۧ-H&�M�ƙϘH+�iJ�(��5|�c�9�u/�ٰ�-V� �J��_����r{\�"n�'ߘm�P�r��}�D���?�8[���A�(i߹\��N{��ƌo�-�&�W;�ђ���{�vbR�&��犮R�3q�9F_!ҿs&�o�e�(�V����%�Ȍ:<$Π�	��K�[�,q|�y��LOw�2��v3o��`���:J�Ÿ2���` ��,�]m{L�����]�vOļVe���늕N��v���2d7uI�)��8���0���Q57������4˺&��u�;>�w b��V�4��I�;�lf�v^�!��n�0�0�@�����,)�Xb:�N�>h�����o'���v=b!3� �4�d�C�$>qvP+l���<c�W��Bj��֊��\ƅ�=�����R�+>�-���Z""/��Sd� m�<_��T���r��)��{��",��5��3�̬�S�"n)�04�ӧ�n��ejfC�]�Qw��p��w�0:w�i$����=� *�7������ǌ<9���@VO4�쯪����ͱ�����3\nҚ��bR�UNQ3��x?��0���F�^(+�P�������J,�"��/ �����������F/Ud�$��σ
��u?�뱉��k]�\`te����)����9ۄ$:6H�v��y����=]}�/1�{��[�G���0'K�A�s��>t{�Qo�n��t�M�Nf0y�l���~/�[Q1'%QprvBe� �C��hqՒ:�I|��)�B�}��T�)��ja�r� 5���o���53�6^����klkzٯ��Ь��:\�
*ՕP
�yoC�]Ra߿�1��~Ur@�z�|��w�%�wƟ��p�d��	��j�ߣk�-ß���Zk����l�����R/-H��W�*au�ӭimEMq`D:|���Q-k�c�:Q�蘇�ī����9��GK�a���0{T�K�-�)J�3-�5�Z5x��G���e�,<�7�@˳�����D�9c�~l=fܱ���{�
�?
�*j��2}���z�[N�ʥ�9e�%��a�����a[A5��O:l��t4,'U��G"���ÛYA-��+g���S�饾`B*���w�~��n6�y���_�L�����;�������T�`=,>�9�\|U��2}���U����^6�I�-Pfm�,���W�����#��!��������W��i!��=�J;�V�G�@������b�1�M��7t��#{;^���Eg ��I$9�M���/���zJ�౻��>2k��r��ُ��R^���L��i=�И�w����x��b&���ŷ y�s9׎��6�W+�=�����2Z�k�T%?EI��>�|�����ǌl]���B|��2$�����A�o�Ɖ���pU	A <���	��^�����x�.�K%v��%/�O��fr�B���>�|tx,�/��Œz�I�&��W��F�=�ծ�F�]�*k��i�_�6�������< �Hj)��&Ɋ�N�/��	�.1E^^�����0���j���9q�S�����V*��I�_����l�ك��(x��įa*X {����Wi�V������x��@Zӕ59��d�u�;(5��iJ�*�Qs�-��$9y+];N3l�����}�[�8�$���֚Pk�I�/h�Ǌk�2s.ˮ8{��il�c޷ϔ��W�y/��um#���#�Q����"<�#�~�y��d�)�f����j�	
>���eabs�׺�6��>��<y[��������,�i��<[�l]�m� �J�����^�#�S�n��*���W�q��B+f�S��3+�C���KmTJ��3���T��h�����z:�o�҈뎞����}��$�4���/ 1�n2)�m���0�\N���tM�y@�g�8'ƵMf�m�l��r����ĉ^+	l�)t����Dv̥E����R׶�%t��XYZ� P]���z��ɩp�S�ɻY��1�X�+B��E��u�o*�Z�*��}���@�<�o�V"��M�&⌇y��	O�~�A	M�Ҵ�2�l]� ?�2�B�Zc�Ŀt��*<�Nko<-y:�r�2꟤[��{�)���Y�D$�`T���v*�]8�#w�O��@BDfm(߈�噫b��HYT@ʰ�%Ve��$��c%�}�&���wx#�*y5�3u�>�L�eYo�M���0@|;PK�,�I�7V�"#����lp�b��2$�����d�P*��תojh"̥�Jd�锄n��Oq=�O�b��ӱ(�Q3���޵HO���Sb��)�
P�tO�; �JEy���}�m���Gr�su'�\	�t5g밣�{x9�fHD�r�[�rrkJ����};��94N=�?)3=�\���9UN���	�տmˬ�h�sc!�.)&5�f�郠�姢����jS=O|c!Q?��?p��+�6a�O�p�QS��_P�З�7h~(�y�D���` A�t	ܲ!��]G3�P(7����Y�pF��wc=a�iX��JG�c��|��|S1n��,UjO��B��`�w,b�r��yRo~�aVk��U��-��3��G���<�1-��E��������'�����Y�Wiĳ,�5??��A���/���g�)�9"��(n��)�˗�������JFF�_ �x(�p	�I�x:�LՏm��=�L*A�X^g�:��^����ۀ^��>WP�e�Q����T����Tf��cp��pQjq�3#J�ŷ�����Ax���ui�k��^SVr����|ɂ�5a�Ȁ��w�6�K@&�-i�뮣yy�u���ó℺c�h.��	��'���<��s%�s����a��ɤ>D�\߮�8͘��c�;�yh�gj�&]��O��A�7��m��>�ҿ����egg��ܪ�|����+tg�I�a�?����ԫm��bI�v=#�jf�d0_W��[Ї��ʬϞ��0�W?h!�N�9�$�YƲ�o�L�+���IF1"8�bޠDo���v�o��MA��@�
L�>s�E O��1��W�����bk5r�>2��c��\Ƌ���=��:m�e�n�R����5�k��r�7$k���醕�t!������r13��(����v�z�Є��9��=���Iċ�ByV�V�?��{EP�-�5󛊸�@�/��U��v�����ѳ.��D��k���~X��[j�>[*_��go�e	fp�l�'��	A�0pGUHk[�91IV��S��S�$҃TZ��dg��	���ȺR�i����軞������=��G�ko{��Jż��b�eH���'����?�� '�v���܏�+?������,dg_�mM��d�������r�]W��y���Cʪ�ʾ)�z�� {<iբmԿ�)��c��Y諪u�$���f%흟%�g�d��ax�?�8W�W{�O���(-"�0W+�j�������S��BC�7���-чݙ,��U����Z�Ϻi�J�WcW��=ok���U[?0bJ��7�h+�G5}�zSK0��a���V�z�������/�/f���h�mI�)	fI�E�\;�@��
s�B�dk�z�_U�>v���T)Z�j�0�߶���vBJ������@=bJƮ�ts8ʴ��GEJv�#~?��R��MJ���Rijk2W�cm�wޢҚ_�j�u�ĝ�SEǼHv������Nu^��q�8SsQ9���)�h3?�|�y�wt��c�.RC���y@'�����o������r{O&�t��R�M�˴���L�=�����1��-��R��*&pP�b`k�SM�i�XOU4Z�7M�S	e�������9l��U�43ad�]s(hW����L<ۼ@�aSh� ��M:wOX��M�U��v�:�c{r�y�5��j� ��9�ZU�TkB��y���9國ܢ?}B�(l�K)�����IĦ���*ٗ�ehw�I}_��i3�����~��5���RB��x����������]�y�C��Bbɷ���[�9�9=�=B�HL�^�^��1e<��p���Y�Wb?�c7��Ŭl�e2/�mߺz���p7x{���o9������$���5-�Xg�"#�>L�Z�]
;�".F���f��,�
?��K�i#��V<���Qx"�{�M�����/�m1[{az���#k0iP�S�āw�T��M^6�����l��'���c����� 2U5U4���S*�fA�>[�u���\� �|����^y���R�t��Κ���FQ1]�wC.>���d�и2)�ٸx�}�9��2��%=vo�ظ�S�U�2�G����eY��Y��@sf�^*���T�#�]�M��[�q�Ƚ��ͫ��k�"��Q:"�ދҧ��TE�5i�AM@A�>������������8,/�sb����R��Fz����8Qhi�i����A�&�� �Pg��DRu��;�����J�po!�j�vꞫʏ /|6�vݶ�!E��J�9nR�7/d�`�݈۠=�^7�Y�q^Ʊ�����S%`�ɆO�� ײ��+~�m�Qn�S
��a%��S��}�T�EJm�3�8}��|Q�aW@�l�����ܠ�q�_�l*��9�<8gѭ�){�#�"�0Z6 L���
�%�����Y|f_�[L�'��)�^�9=�J����a��	�Gx��۰q!�P�/���h��s�Sܸ}?y鿷�v��^�H��W���W��Jv#@�#��+��@}���g�ٞ����	�%��ê}U��[q�:��&@��PS�
�,��D%ˊ�:���˓����qW���ZT�$g�����d@�?|kk�!9��8+�/�:���٠�-���M1�=�Hzá������9dNl��Eq�*��:�ľ�������5t�h�O���ܜ����4�$!�~��.�\�nkJ����	"���O�W�-?e�&r��O����\�t�~Z�����,932 -����켶� ��՜�K�@fjv���aTZ鼆���-6T���e*" 4?�2�!���$ K�N�k�����������4:!T���i�J�ϣ�j16hf����κ���T»|�gk�j�w��@��s��P�Ҽ�s5jYݱ��WљT�����}��>�|T5�TV��Q�-c�����:cBn����[�+q5�me��N����+	l����aʈ!!쉰����)�u_0�"�1�U"�BpU�j�������Z%�	�y��� Z=#�v��Ob[ͳ�( @���(��c3d�} -���?�2"� �<��8}��Y����$g�*Û)�6'��b��,�-��F��¦	z�|b���&�����U�a����
k�����m�T��ۓ�owwq�%�T�)
4,Lᾖ�r���
��T���J��k�c�b��!|o��qR�[�m $�������f>Q��ј|��$Q�J�&��S\�������yP�Q���g>P��.�Iq���ʞ	.�b&1o�N�l�ܼ��PV��Ӊc(CV��3��p �h�p@�ԣ���'s�?#�DkuH�2ȽQ��׺����U��������{���?���%�`����`;��(��:t߬b{�)Y���K�[�4��(�h
�lGME�OZyHx��\��fLet�5a���v����;�b���Ey��fu�]݀êS�ћ]��jh&�?�:I��y���Ϸɦ���./(���,@�3�,әz�0�v��ɉXd�^�ٸ��7����N�d��n��fR��{ey��x��#�dwU=F������eC�dt�����\_ �ɚ�拳�;ۉ�6�뎵,V�.�٩�T�Oe��VK��?�M{������iv8m�a\��n�]v�?ͦ���[���<,)ꩩW���n�ӷDüR�c���>h�H40�R �� �+�w���N�"7�x�K8]������V��t+q�}��S���;��`��%f^�M��������Xd�r��BX�:kc����Tڵ��;bϾ��?���z�=y���qKV��C��<L���b=�J�S_�b�C�~m�T�4;è�^�uvx��;W*�����mM$hA->�m����;�W�npF0��=�t���˲�4�n��T��>��f)J�����1���]�B���#MH�{��L��Et�#`�ά��;6�Cx6��ϙ���vqkU�$���guв��̞r��i �8>��F9���O� �[9nW��o�¡U4�ʀ���4�ۻ΄N���&4�/>��i���Q���b ʫ�Id��:m�\O�Q�̬ٻ��W�:n̡<Ǟs�niZx��$�ޭ��m�G����.=�daǾz�MOج�x~�Ҥ
Q@��4�K*Gi]�J$NJ"��0�FP��/��+}�w��K͚��)�pUe�aB��}e�7W�]ښ��5C���av��� l��!;|F��$u�ĸnv+aQ���>ݦ����N�vx>@�[���}�5�M�\]*H�A!�� B��@da��%�;���V6��>�f��h	b1�NX,��6� Y9��$|P�VT������y�����{�Z|�%<!��k��Q@��16�`Mc��g6R�W�Y�dnɎ��JVf��%�GqQ�h(�լ�w�^�C1y��ڑ쒉t��v?%n�̋�<�Ƣ��Q{�:��� ٝ�=}���-۽YU���c�O��$��u���'��c�৚8�m�?w\�miWt��l~M�S{c�W�+ Oi�Yw�(�R�j)�h�q�5�\Loa8��i��[��e�x�}�J�w[�r�a�U�L�r�a���ׂ�����ֽ��Y
 ����4�x�[��������(��me��y�/���D��a�@$�`$L5����_���'ӑ��Q��!ela��c� 8�Xn�X���Ӿ�+T�/41.�F���?6q�,e��#����-���%GT}��I�)���bI��M�Z��'�I�$�6n<x�L�PЛ�[w]���;�8�ӽÍW���>�P8�]z�ѧ�?x9P�V���i9�~�[@�|���[$� ���l�,i�]���AI,�J�	����L{V\��[�&?����p������Qƛ�e��o��t����M.��Q6�[x�-���@�KW�e�ܹ��3 �gޓ+P���OW$P�Ж��Y�Db~�Dǿ�K�
w���{$=��cl*5K	�����9�\cOy��vܷo*�irm,
�tdg�����B;���|��Y����A�Q��^�}�#Ȧ��"LV�O��n�}�	Բ;�Vm�ޓ/>�`��$��Ex�M=�[��+Kẇ��1;��縴E�M1��w/(�T�(�]�9S5(�c{l]Y��w�Od���tc4;�fV�k�"�ne��O!��*Uf;,+�<�?��W����۞����/��d+3�e�]a=/��yӺ!�3��o��^���KHS�L2�d�>�{5>iA����m��F�*�nI��_~O��;&��	ܬ�fU�U��nb���0_C�糒j�S�^Y��#9�''/&���}*Y*!��ŴBX�����~�D.;5�����4��D_o�rb�ݮ�!����<��m�=�{���I�O���l��S���H�������Ux��J��m㣋O ���_3�������n��I��,t�X���a#��n��X��H�zL�:.D{��eW�I�!{
5���ux��۫�/�~U�d���B	��C�xU��Z]"�g��!����M�"U�,TC���&��d������\]q���J���
T������-���?�FN�S�͔�=5�;��ZT�x���t�_�f�4�����ۨ׭��%<@�Z�+��9;�Ε���s#|�.W��,�:�|�o��.�nI ��0	
�(���;C��˃Ia�'�"���?��\*�h�ď�����ߝ�����������p�k���~��>7�F$��ҩ�۳n)A�&�H�u2���o�E�y�+����	��fo!ӆ�`|9+eWO�h�%����
�ﴷM$�q�k�7&�ohSj�r�4���(ekIBd��M=�42@���v�h@�����R�	�L��tND�sפ�E��Y�L�o�o<��R�<J�6��.=��wC�\-{�?�S�P욹媩��X���H�����|��n���n��җ�vq�{m+����34I±>1�+ɟ�b-O{��K�mha��'��@����o��T=��'������A��X� )43!�?%nϚ4� 0T�ļ7�D�"��®q�]��-��j&�z���R���3�P�aS�YЩ��^�D�զ)#�Gϓ�!;N��Z�2G��r>6�A|W�y��IQ���-�o�/��ny��[Jl�y�H��f�������P�B���!1Z&���'`fn+F��wA�� VV�<%l�:Ԥ����ٜ����A�����@
^\�8��c� �5�2��*6�<V�� -{s�z�Y$��#è�hLR��#�U'Z*U��.����K� �o�����3Uq��5A�����O�0+�I�2|>���;�ձ�3�y�}����A��ŦM�#)Ԃ����t������Ǝr��ޝ�"�> b�kQ]�NC�� ����ȱ"9=y��8���HuN�u/�Oj8}-�fS�V]0'��3��꼆�ӱ���9SQ]��e�s�gO`>тr�߿T:���G�3&��t+8�\{�O����Ck�>�2�ꐞswTW�����0$�0��M�)�9�p���h�}��噯p���f٫�[��@����SxC���V%���PS���a�X`p�D	F�af�#8nt�"��B}��Uy�I���d ��`^������2��Fa�BͣiUy\���w��2PU/^W��Ϫ���)x����Ҿ ���`T{�@��+C�,s>�<$�4�j֢�ѐ]�s{	C���oWl.%B�8Բ�*����l��b��{ܠ��f,�0?=���5��6�$r�n�F�o\˦ꊋBy��D�F�zk���?�P�VFi�!B	`�y�/��6wQD�p������β:(|��(�f�6���Mu0��.�{��p�n#�3e7��w�������:�T\=qڂ��t�E��s޹tb)c��W��8?���`1u�B]wz� ,��k�9<��3��'{z��ݕ�n�Q��Ϻy)ț��I�����!6rI����Kkujy{�[8��aNy#m����~�}	���0�e�5��H�������C.�fW�D���|^�k�o����� �V,��a����ɫyD�ew���"[�)'��g=��-�ϱ�n�)N�`[,<E�3-LC�}���F����ɨ�IC���T���;n�>=u�Z��wt*���I����gX�O�/7ި�N�=K�����H7���pտ8�}��5E�y�h��E�5���2�@�|�8��n)��x:5���-�������3Ц�mu[�~T��
�ލ���^$7n)����h�s��~�9�r`A����_�Cz&ϧ+4>��ֶ�Ks�oi�d:��k�ҶE&�<����=�B���{�Ő�]���G�,���܌�l?����� ܸ���­<<�Y�∧�Q�#�, U��V^��� �9v��-���{�O�#�Zg�;�����C��nK�(7k�{����K)�_�!"Z��G�T��%#�� 6�C������BiqG\�Dj�u����e�{kU�ƭ�An�}e�������9kYm?���\�E�1�Fb᤹#R��SZ��ѻr$w�Cg�A8�u/k� T�9��U�<�n�<=����'N�$�k�DZ�m���hn�aQO�g�We��@\���4���Ux�}Ĝ� �F�I��"a��u��ۃ{�l#@zF/I����^c�9~>v>��J�$�`$ֺxg�x;X�]����|�*
'EC��/��{)C� ����Rv���k���x#����_�=����[�;��*;�u�; Ⱥ�,�	J˱5�\�\��9�NV�3N�� ^<}�O��}��i��/	g����NF��W�$�A�/��^x�S�֍']b���X �5�i��+�]1��+��Ŷ��H|O��*����cSO���t2��O5�᦭g��v֋��![sq�}S�2ڽ�.��T�qֱ���cT��	�`�|���v��2�bf�����<$�*�ɠ��H٬#&�dq��C�bj��e3�N{�L���3�6�tc($��iB���Z��z�7]�^X����^E�6}zD�y���j��sMT*g���,���
���A�Da!zh͋�������&�xeT�"�8��Tȯߏ*`���f>`Z�(Jץ(Xr2x^�*�!�ڠ�j���j�C����vN9�������|~m���5���h3�v��%t:0��N^�b���W��P�7|�?��wL��� �����}C���o9�6)�urZ�r\n�DD�� 12 ��/=��ګ�w� �ۮ�
�y^���N�����fu�k�Id�ܼ-`ӂ��9��:�3�x�ͩ�i��$ز&���x-6_d�ߢ�N8/S8�k덏�*.h�G�_�flD�aXޮm�sn�n�Ӂߡ�>[�u.���;=�?���
6�t�������v��a�9?���#�	)r}-�U�䝂�]EP�ww�>��A�o��3��ǳ��J�4�0ΔYJ[ĽX�HYfiɠ]�`ga}�gܜ4V�9�?���d�༞���X'8K;3@V�%��:"�w޺�؆����)IZ��ݻ�պ��쎨�y�N�ȳ���>H+"&r��O�͙��e���{D4�a�5D�����lAˢ��z�Mڽ����;���B�?~ך������@K�+�}�](��~��w�<��7P��j�ok�8�Q����&.�>h�M��Sm^M��ȫ�Oϴ �GL��l�J5@�{/��#����ў���ǟ�oPKڇ_C�)R��0�+1��@ԍ��=�����/�f4�߸�2�b�m����=�	����7
�0���op�]Gj(Xݵ�^��4P
F�{�Z�+��p�']�����8J���!�j]��/��f�g�A�ݴ'}u6��>��R	�Y�������eҤ��뉞�k�b>�tcL� b��G���m���G�f˙�i��ꚯ?���6�6�zq����~�ڴ�e�kE\� �_`#�ųj�ܠ�긻3@�ӽ�v���X:���'�~��P����pQ���S#h�o�c8��	`�������䙏4�V�NKBF����2[B3����&�'��(*�܁�����w��i�H����07.�n��N�&��(��"�\i,�mj�*7�vOV^IF�u:����ȈC�~�=�0w�
��"/���^A�S#��0�Ï
�o'������ϧ�^c��<����[m��a �-��s.���=�VLa3�Ą�	P{]��Z&�wbuG;r=q�����4,���9�w��f�m��{<Rk&� ^U�P㮣2#�,���U�3�M��F���B;MF˚��}���]m]	=V9[�}���4�{k��*��O���V�ܿ*{���4�m�9#��Ye��K�A���)a���b%��I�<F���kƳ���)�W�u������-��j���P��ܵxKphq�
�(�w���Bqh�Hq� ��C�����}���+ɑ��̬Y��Ι�?��6�1�?�k,�]G=f��1�0� DI�7��u"IO��tBӦԚ��;�+�ߕ�oE��m��ݚgt:je�W��!��/;�h4ߢ�j�g��n��7���b<��ɑ�eş�I,�B�'�2G�������cp<���5�^h���� ��F�X�V�YE�Ѭj1o/2��p�6�d�~D:D��mX���+^;x?Ecr5H5�o>��ݢ^���|'n�h�=�Ck_�w�w�'�@t�o���"��_����PN�1z��*����D�m�s$�M���e^��yŴ�4���Ü׌�`��t�a"6� �`;+mS��8J��`�єM�J$YnA0��&R�۠�o�֓Y5�ni�0_,""�� ��}z���ē�@D�@lg��x,�.�Љ�m���VK$��f�Ǧ�Gͻ�pQ7���m�)��63fS�!3XK8]�ν�F1E���O�|$�B���Vw�}#�6^|�Y$Vd��Y"L�ǝ7���2��A�6�;��iu���� �e� ��h)��j���.���0��;n~��f�3���� �yӮg������X��Vb�5��N�W��g`t���˗��Y:A{j�/��\��NL�����c��-��+f� ��	Jv�,/-��hY���>b���!����T�C�q�+�;��|���
P�E�=||�e���x��}�1�]��>�	E>��	�E{�I4k�O������^޾������$�Ȅ�S��,#�Sz�Ƨd������>�����i�9���t#�Di'�KSE*\r��eA�}Ҟ7%����$:�����ن��S�t�g�i����S�[z������I{B�gg4�E4 ��y���]-،��SP�_&�n�dB�i�W�-�V�pb�����ŒX��2��+��]�DfVgz����B.@ct���6$�˙fI5�1%��⽘�?�[g�)�'���5�:��i������:����9�J�3�RUPJA�����L��_�`�6]Y]Q݈!b�÷8֦�ē�2B�y<%_8S�56��;�='��"�կ:�{.0��s\�3I,Py�
���g?���_QC0�$-F��	����W����-������c���ߨ��b�T��i@�Wu�*��~����(z�=6@��an>�1H�s�h|D@1�a��$�a6�<^��p9{qBc:�3�&R}n]����͇E}=�L���٘����T�Ң7'�Ct�}d�P������R��B/G�:�-��7-�S�M������Z,죩i�3�c��i�+V��Z�O��)K��:��1�.Ǐ�п�P,O�*��I3a⡝ʉ��w�"�}�*$]��+�L>�^��>�E̻��^^��^��x*x��Jh���cɒ}k�v4T~�x�]�d� X��������H_�Q�Eϲ�o5 ��f�u.�e�r
�
̾M���M�Q�;�v�2/��`'"�
�Mv�;v�#�-��?����cSl�pZb-Z���Y��B�Ζy�BjN˂�b*>e����\:�\ �W�c��FŒŰ@�A�٫�[��P���y�[�c<5�(���wHâW�y�Ns��$�5˂ت
ii��'�,Y��<�{�6�d�U%��V(���  �)�����=\� x�=�UB| ��L��׆��"�A@ t�3ϲ��r�e%��EQ��z�$��M��l�}��A�S�f>�ʦo��p6-2kp�7�s��i�����+�k���O���(�5��5�s���Éi?��ҙ^���Ȍ�댾Ǔ�?��m�y]j&�#x�ʠ�\�C���l����4[ S'd������x��u��y�K0M}�W�
��ON!��˼�����7r_���K��G˷��(6�p,U
�ү�&ė�"��5��W��  6{V�x���ݳn�U��K����?b����@��\ �)���*l��f�xQ�l�q����Zj����Gbh�I:bZ����S�N�Я�1�/�!�=��^h��Ӳ]S�%�O��\�o��>w�Nw�c\�;L�L��ed��
��.��̋���X��* ���o��>���V��������<(�B�8H��!���[��P{��cP��.:�� ���|%t
��v����ӏo��:���M�����̓��+o����;�m��t퐛d�e��݋��KE���bA����1�\�i��+��|,��c�jwsci�N?=��Q�����L�=��IW�A�{U�ϔ�16�5��m���5����%t=7�
���}_�pDTE3�P�P�t��m���'�3��@~n؉�c�6e�����'��/��ы�]��.73�������>Sm�Dq&Y��S����{����W������iR�z>�+�Ǘb@����26�H��Ps�G�~I��K.��0z��O'nl��9�u��t/���2?=m�ȁW[WgPH��ֳ�w� ���Dj~>���m|�Z�8�	u<�Rg��A���m~����Xx���5�&��Z+ܩ-V*�iŅ�|��=�GLi�2�Z
���jJm
�e���zDl����*`�n��5�8�)5��T!hɪ���T������X�fC�c�������EK��IR�w#�F���b:l����?}�o7��N,�:��+$[��,����E`ҌYr��qP�k>��
GV�<N���� !�y�J���h����B����E�a�����ۗi�����5#L���h$��2��CM)L��T6jRꖱ�+euW��FmS���K�AI}PԨ(_�l>��g�E�}\���`{��5����)��c4
���.�y�aG��> �xSVf�C`�)�x ��G�Փ��8}�da��bk�VLh���6czc|���\�[>A0��SRx�w&�	����wzuy0G��sp�����/���?a�M��ɃZ��tӠ���:⋥f�����pde��)���l�A=�A[�bjy	��gy%��ؒ�0����8��ɤ��)Y�j^;\�_3J��,�u�&�/�j��#_�7��������Q����l+������#���ܣuN��˦��O%�t��=�[�诨�$ȃZ̸Nw;�ݿzl �.G��gQ���,�$��.������y�/��ݙ郁��`��$O��9����Lղ��P�j8�� ���L�w
�W��yN�_~,��~߸ו�����g�����j?~}��P�lA ��ͥ׃������'>x�}4�1�ZWC����!覞��in��Z�(8Dj���T�/$�����T'�R46�����*�,n$���/��z�@Z��"KE��X�l��<�Q�^����O�	�kr�Ѿ�TtG{[9�j�d��(w`snw8���Q���@jt>��$�F�~i*v�<w�mO�@ĺ(��ICd��h�*���L���G��K5F,�×�t�׶H����o��N��
U���.��UK�����b����<�b1�k�����JǼ($L*�_��{�n@]�"�^�1z\#���L�zy���0�^4�k�*�-�P8���W�SV���Dt5Z6�:~��!�q�I�*���>�:?0o�s�:�O������yFA5�ޗpS!�R+%B����l���N2�J���U�!����.K&�*R���- j�x1��sҮO��e��9�5�P�������Q�%�`a�������XXC�1��|�2y�d͂�ŧ-���'?z(Y̓s�9��8~��	�H�:�,�q\�� 3�3}.'SeۊZU�;�v-��r�7�u(_�{�v	�9]�Л��V�z^N�.&3����^�: �v0E>�N�4�Ib���h?l����<�z�L��(uw,��[=�R����aI���k�@��x[F��N�j��$Lq5�%D���|Kt����_��.R?2Ro^Y�ِ�l�Cz�úӀ������C�ӂ�>R���!���R�b]S7�m]�'�3;�����ߦAڼ��?CY�.G�3FI�E.N��3]7����e]��l��~�n፪�����ab)��Z�T2H̫��p#(�ozi�O+���^^\e c�ad�N���˗�ܡ�4c����+�Z(�� ǭ�8d�d��W?�	���L��|M���_kqF�̊�� AXS���`cc��jI6�vrf�*�_�)6؟�+0l�q�}��v�Bd��x���NY�j�]���D8�zT�4���U�:�ѯd�sԎ�C��=R���ZX�[�յ��"�un+�w3������ ��Z�7�@���X��i%=n
���_�w�=#Y�	�S����$�A	�šfK7H�9���- 憗L0�D�W�F��t�3忚A[�E;�>�R�o�p������pj^�������~Sm�s5Ɔn�U
�Y�D���.0R>�e�tk�|n{�K�S��9��(o�2�ܤG�ԅ�Ut��$�{��;��<R����,I/��/8�N.��[~7��8RW�'Z��o ]�n4���}M���p�\���� �@0��K�nu��?�(Ppf{�6q9W)��:���WzJN��5Ceф�~�;�v*1m�9kR�A�IMv��:� Vt,�
�3��oȹ�N+X�*�h���۝��X3�H:����V�����MrXXH�V�9[���@���n8I�q�sU��|�,Iq�Gk��ۣ
7��0�����~t�=w[B�zf{��u���I�c t�����L�N�2�*y#�ɲ1��o(5e�(w��>�W_i��_yk�r�H���m���J��\�����MY��wM���h�g�Md_�.��g�/�h<��9, e���)C`6as�k)��T���a�&��~޹f�lo�� E�����m�=����Qq����bZ�.�e��K'�b����5�.��. $b���T��xn�廡�#5/�YJ�1krN�X͡O��5�_G9g������UF9.^��5����y~;+sܲ=�ԕ��v��4�m����T�[ˀ���ʕ߫n��ߗvh=�̖�X�2ꄬ�[jPE�c�!�]#h�W���ydr��d<��{���^��\�=�s�{� Q��7g�V:w�h�U^4�;g���9<*�D#×	��KO��]�&+E�*4���T�z�:B#�Og�v�xVbR��r�ڭ�O$����!��C�d�d���b!^�׸�Nf.��EB �b!�9��۽����GZ;�hF��b�k�ރV����/T�[fgm�w�]t*�Ơ	�E/�KrSG��t-oIÚ�Ʋ
�Q<4n�Ñ�gk�	�?�n���̞��ʚGTO�e���u���MaZͿ6�����r�'���켿�:n��a)���%�{��0.v��3C1�pS���[���PJ�e�[�T�����ͱml�4X�Up��c�%�4��Ȏ�u�|ws.��G?���z����
�6� ��5�-��n"���7ί�>.�1b����������o,i����syHh����:��-4]9��=�%	���F8gK�yx����W�N�(]U�1���h��$甞���m<��>n�"��	,��/���pާP���I���7�S�R���g���������=������_/����\Z����r�׃�P�>l�Df�>�K��P>��}�l�����P��P���g��]����YĠ���@�U_�IYM��N����JX\�R�NaX��ڝ֛����|�uw�m~ޫHفΨ��+a�L���(������!����~�'W6���K͖����i����Z��	KM4�
7�G�D�ew�26cT��\6�K?>_6�&�=8w3zh��\�{�w`dD0؆૮-���6��Jx\���SM��TH�׬�t(mp��pK��I���I<�觺��}Z&����x2]�2A���h���'�t�����2U��ƑP�Cb�q������%���Qz�s�$f���$-�]$���l��D�f@��ćotS�:G{ۺz1v���"x�o�GhMU��in{��Pj�Zix���v!56������f��;b�6G<:�ם����{B��C�.�Me�U�i�������7o厁&_;)!ƈ�p7���]Q8�A�`�<DIz���tu~�bzZ�0�Q� ��
Gׁ�4������봥�bs�����s�]Ł?�F��ݝ.,ؾ
�،q�k�PG���۪_�����{�̝Vl�{�)0Y��'+w<��]
�+��E_.�4r�\�v�MJ��xS�4c���ކ�k-HM���ߛ�>�ě�~�0�7���"��>@[[OF�D!��r�[�1�{��b�P,HF��s~vA\�ip��)��	ye��xv���{��⫑�3��TF,w�f�*m+�����"�/�Pנ^N�m��:�p���ܫ����o�ح����ha�t�����6�H��<����s�x���C��EV_+f �C*��o�o,/�	�7�� 0%��ɾ���~�1���c�@��]���wK-ƳM��_�/S��N��Wn��G�5��@t	/�=ͭ�����U��u:T���p�+b�S��7E��7��L�R�Hn���{�0�I�.�vL�1�p���b���fܾ��~@P4Q�0U��ޥ��N^>O��#�%����+_Y�����5tL�S����z�q� ��ֹ���jcd��O�������!��-l��Q��^ �n�ٗo��aJ��)F�C�+��Ge�1 �t]�O�y�0+'w��/1n�:�K��u7��3���ͭb,|-���[��?ٮ4���|&ﵘh��Hc�1����IF8�������#�� >�����<v@��̸Pt}[-�����Ͳ�AAX��ld#yS[K#��>�V��ުXV�;�J�e���n�
�r�qʨv�;����d5���}���aw74�}��Q��\vGFǊ!�; ]��!�+����"�[��}� �*��f�x���Z�5l���F"�� $�K��Ձ!,r�,X��S��Jl��f&2a�3�xiA�c�~׼�r� ��M#������\���܎����I$�����2�C�O,������^;������dFY>��q\��*]��(��gq�i�E��x�LM�J�=�l���s����px&j?|wԂ���##�`����7g��p@�9��$�K�/�`�^k��>un��~���<Q$Xl��OV��V<���P��7��խk���?Pv�`�M��|Ym��$���n-wIQϝ02/����`A����c����Ư�%aR�&t���l��-R�Kls�������5���p?��hC坢�]��k[_�Fs<5���w�Em�+/�e	{A��[˲�V�w�>^�͂e!�y�vyw�U����4�������o�����^�CElP�@ym���i���3�wy��:����n�>Ƞ��	 �
6Xhd��q�B:�����X�u)�YԾR���(�_y�[��G�דW��-#���̒4�4��-�i��m7�e`��Jh���%B}x�T/�}ꍚ�ki�W�ӕz󛝢�k�}��!�z���ƙ��̪��ï_:�-TO[az����m��۪�D�	�O����>k.BE�l'�;�9g��4�V��b�sf��!���7��l B��T����ӷ������"�k8K.�(�|���X��w*۟# v���E��:Y���}^�Za�_h��k9��ТQ$�3F�X_r�:��︂6YEV+9
��"��*��b�����M��|�	�%��&�q{�~ݧ����<�O�s,/��x$5�\�ޕ�w�q�}��	^���-��{m�I�w�>}��
c��� 7_]!�����-|��)��7{-�Q���������Z(z��LWQ��`�?~�d�,�2���qy��h��W��q�<8<�VX}��Ï��#�u�4��x&
�=5��d�	DN�!O�ƟDs�p���j�?��;���b��޼I�����%���C��.?��R ��u�k�Ś����$�1�:��=��d^�O�{�f�G���'�Mg��I��Aݻ5O�ߛ-��4���L�A��,׋�8� f��X�ަ!Qˋ7�z���l�Hm;����'�#M�¿Z|�C�eW��V������5��g��A��?�&�g�M�����n �}��z��(q�b �YRZ��<�I��B]�w���b��K�O	U���kJen����Ԍ��K�דhd�Y{�*�?h�O�-_���>�d7g2_F��˶E����[eG�]@�
X<��/�9KJ��J�T��ޏ��/)o����
T��u�����cM*^,�"	�����T���GH����`a?f!�6^m�ƂrJ��Q���!�m^w�3~W�[��V��0��Q�;��ث��4���r?;�&���������!3���Q\�v���	j��i���s{9��ɉ&���%�{!��0�Z�ˌ���,@���2��t򷞳���a�h��t��4���Tb�	������g�����搢�?m>4�8p��}GuNv\c*H!W�I�敕D�L��>l����J���7����q��������t�n��ؖ/�)1�E��{_��0p�)P���ݘ���9�Ve&O1��>P��`�>���찬��ỹ+}u^^S���^�T���'���oo[�τ�
������ݬ�=�x���[�o���@3fO^T��,y�hn)Ё����uP��DL���������JUx&���U0����2��b�w�t�%��|�Ks����PB��`���߂�v�ek'q ���a�j񕊒C~=л2�ϋ���u��'�JbO�jFn��x8�ES�x�*��<q����=�wH�Y��5[Fr�ƨY2�����q��թ����æD�G��@��y���a~�4*��>� �>H��}���z������GL�WS��ҁ���"X�����R���3�M�i�.��\����G�?ZI�S� ���i8�׸�h���{Q\�sݢ���8�ʇ�2���]�����oE�%��I�rp�*��g�蛅�봎17b�U��S���.��k.¶b��{s�*w�R�����ֺ4�	[9g���y��:�V3f�B�Q�*���R�������ߙ�ߡ���cK�'�����i��U�/N�|l�l��f���e4���:����k��Y/ m�&wQ��=�Ш����0�ɧ{�׫�CJ>�䣣�?��G��=T�r�����Jע��H��<x��Z�2����M��"oZ�}sc�+�Jx�7ФeX���/�F����"�P�~7KKun~S���}6v�.v�C�,/��i4҇��&X���|�|5���0����V&��vr�}�ИWZl��O�;�{lN��?v�khr��S���g~,U�2��0D2�2��p;h��D�D�!��r#7h`0���f�׃ʳP��+}��l��f�E\��SS��`��_��&B	�E�et���d�Z7���|K^.Z�c$�K�(�ј k�t�;��<E�s��i���9�W��,�RT�)1Y}7�Z<N]�%l�ت��gP���Ā���춋��ţ���g�̛����;G�Ed���_r��(�a'�/�>��G�'�ݎ  �!= /��;U�%���x�m�b]�S�	nݒ��}�b�z�;2;3���z�r����-2�g�Č`n�	h������P���,�����^XN��Nh��	˛�<�c�G�|a��|ݏ����w�@��*o��0IK�J�h����ȓ���Pvar5)��}_���Lo����U��`�J���֍��7����*�,/G}�Wi��߻��f��K���hm���G��u4���SL�Nзi:�ܬ�Z{�n�����3˃� �̠z�;�g�=�0_ˇ���CkО9 d2�抆�j�n,x�``�И\N���ډ"�����'P�+�����~�����P�����|zt�C����߻ߧ|D�I��!6=�l;�!A@���o�v�T�{D��Ӻ~�gw������L���f$��vK S�b=*����w[o�:Y�A낌5�=\F;FL�N�eወS��Q���u]m&���ʳ99[��z�?]m�9���k:@��f+�	Ӥ�k&�W2�ɎxK�<��p�'��s�u���ݱ��mt�XQU���Tpl�ݗH����"jb�V��-R֎����Sy*�.F"�<O2� ���S�!f��7�%��7������?�����6�n�0�
�چ���S�mI|(S�I�����<@'�A puu�70�}0
E3��{������9�2�5	��%�&�#��0Q�(�-d*��{�c����PhW1��h��E�rP�
��������Uy�D�up} �xį���!��`�]���Dat���z1�=���,��
Y������Y��H⟢�A�t4=?���!�7�ʱ�E���&v�+u���p[6aŧ��������L��*j�f�qK=ɗ�{�ds)ɺS*�W�����`Z*Cp3������{ ��X�98Q� ��������;��^�HX	�t˧��ҫ�N��fgCHU�T��K�|�ɼ��t�A^����8B��BC6q.ݣC� b5�ě��� ���U�#�mW$U��C��_M��e�o�
ֽ�����c�ű��P���9����U�O��͔d�u,�-�4]'�|��ġg5�߶�ADC��m���Y�?b�=i�F,�G���>[F�X�$n�]���a�F�TY!܄���-0�H�fd��>��p�E���'˲-.�SEbT���Y�:���cL�R��Do�9�&ՇƐa�����g�?�7�ػ����d����;_�Si�܍��4�5��8��"���
��-':g`��;�*�B�.t4AP¹7���5=����/0�`���X�����Q?[�RK��R~�d#�|�6KM�B��0�F��Bu��d�Y5uh=U���o�Y��b��5�Y���6���%�k��R�U�[s1��(l[mC8����u�B#����p��9��D�Y����v��AR� �UQ�d��:�O0���M�]sd3-ݝ9}<��7���o��	C��8�8ct\ϋl�\_���p�4��߂_>���ZW��o�M�2Ds ��Sh�ީ������鏔�k5P�X��p�%b��&'V�$C�|Ñ����qf-��kɼ�"#�C��J~tylv&����ڰ{y#k�[��O%����6�,���b�9�tI��5TȨ]��Dm㈓�o�lZU���܈���"�����W�\��9�Un��Ɨ)�a�SF�Bq��Y�[P�S�u�_y��]�w/�3���&���m�Ҋ�	�ࠍ7*�i�|Uq�y�2x$�xbc�,�S�W���K�*:���V�T�ٹ��F����D�Up���1V��8��ږć���=�IÆ�9V�B���9���|���%4��G7U����9\x���L�M�� �Dp�R3ڱh��D��EzEt�A&���/���ſ��^��Kv���g����t�J�ov�Z&��rt�w��x���������*
�$��0��:��&�k/���,�����������"0��C*7�Ep���c���3����\2��-�@�Q���������)�U�
����{�v0���:2��H�B�luM~�)�~&{�qF@��scȥ��+D.?�'�E��\[n7}�1?�k����Ə��S�q�I�hI�/�*�E$�]�V<�ЬXFS�x������X_J��̛��$�\
�*c��~��>�㠋47����8�GLG�%?�	дE;B�K4%��y��J���-��:��n���ƋT�5 ��5�@��%��c�AM��f��_��d3�|� �GJ����z%�<E�zLY���x���b_��XY��vj�V�ߕ�hs9�LL�X_��K������(��b�v��o���(���R���B)X/��1��`���LE��}2\8�Ħ�f�1�y�KVa߆�_:����:15C_y*oE�K�Iy$.���'|3Y�c}^�F���U�?+����/W��8NDGC�N�w`����S��f�9����~1ń��?��ܳ �<as$W9έ[��ά��9�;��!'�xk�X�"�V\&�R������ƔW�	�� Q����_|��p�Ń�8jA�&�)�թ�
-�Xq'i�Oq�2u63N�vm&�5�:��ˑ��Td�,>ûb���Xw\����W����1�!Ǘ���?R3^���k ?��jKݐ>�.$LY��^:�f��  �os\D�S"[@p�-`Z"gC��������g�j�@�5=$�û()��_d�4���QΟe�Df�XUZ��U�a���˼K������ �eW�W�$�0.6t��v��]�u����wN�}G)���ڃ#�N�4�C+�RR�IL��kݥ#��첊{yu�ZΥ��^�Ե��Q���u'?=�"�ehCכ��S
��yD:�6�J	�Ή�@;��9��ߜ�3�A��� ����VOL����0 �+�Az��R�F������DY �Qj��.�(�;�y֪��������(r����}����<ֈ�z0<���I,���<-�;�D.Il�\��,����xsq�߽��5mv@>�#�>����+��e��
g��U��vUb�L�s�%�b7����{�S��e���eW/�Q�PBz@;�vq����GTK�?�����c� ���Fޥ�����&� ���Y%I��V��,L9,�Y�������y��.�/m�C�����(.i�VEGT�E���.���F�8(�tB�>�d�n���5�M��)w����y���h�Ӱ&���*���C;
�W�3㋕q�p"����ZX':Ct��l�;�3X�e|�	�޷�J�������2���s���(���2�{��G��: ����	7�.���eЄ#��(���t��B�ǣ���\��vFj!�w�u:��Jc���,�bTFJH���S��;�^ه�W*�3r�����K,��/2��0~�S����ǇQ&�iYt�+�
�D�sIM��h��h.^���JfZ��"Ub�0QR�~8��5V9�����_�b����",�#����9������E�����Y�r��,�����l}\M�&�R��8��$Sگ5@��?�����#hG�p�g_T�Rn�u�˃�?�fI/�oX�����IW��jܪ���4�����'�����L6����L����n��]�� uxO���F3A���e�57L����SHN2o���Ʋ��]�\D#���y=xB}���l/#�4�UG,�}����%m���$Y�q�c�.-4��)K�]I&W���ơK��%b�o���)���-��0-��}w����'F��M-���_�Nn�2oQ&uZٚ��,�˂m�nT��fN��W������ G�O�ؤB,��dh�UR�~]T>��
R��l[&���8J�L�3|Ӏ�x�;��Y�K�����T��>$����w3��^���r�����C�o�H:cBp�uZMR�m�>�ĭ���^��Cq& n��y��@���$�ނIj��΄����C���m�
�gM2p�<bA"��\A@,����N{�8�����e�p����ws�#�g�uL��=��YBLSkh�3����p�g±���W��������>�ud��(W������N8 ��9�pݴ��;���Q0fK	J�up.�����"��E�l/�*T����5�zˠI�TK��h[�~�H3jr����Ӭ�޽��!$�T��Xy����2��+C+�}1�k��X6�;׼�E��;�DG 6b�ɰq�WhF��w��	>��7t����=E]�I�_���8�O��"���j�b�u��}����u����A��\y%�p�+��HA��8h�/��y~��J�b�q�,�`C|��;�WvE�nI�#Sگ�-��d,��J�EBf�A6d�GTYz"̖"a�T]��g��w�ea} v+($C��J�1ި4��<�;D%o�]���E=�ƖGg� #���5�1��Jxp롷Ǎ����l1ǈ
��0����C��"f�4z�aq��ԛBf��� N̒+K9����>��rRrQy��R�g��EM&3�Фw�:J_��Q��(�Z�WB�I�@��DK_7;����?y0�m8���C��κP�Xv� M�|͕�l�7w	r��6�M��N�B/���U�\�ʎH�a�_��\�9�]���S�H�,_��z�LT�z~���������¿�7z"�]�b�O�~�ۧw�>���V{�: ��I����`Z6h���{����%߫�W&D�X6��cT:��M��a��Uƨ?�K��N`�ȯ҉��U!�����Jdo�@���)s�f�2�՞Q������a��#4m�a�(4�A�K%a��Q7S2�-2��V����9/-RNC����nrC���4q�($絬K��=�+$#z@�1y+wg��UKh�m��{�HA���S��\������{R��=@���-?Y���W���t����4wqwdWy����#5��/1�c�<�7��\��I����v�8/ƕ����8mfs�^��}

�L&�>�D6͉���,K����	LV3�"�[�/��o�'�WDG�������;a�i-*� ��lV6�t�w�lj����=�P�׫�+a�bΗY�1	߆1Y�i�����7�ԅ��obxjβX���$�����^��iE�oP����߾!W�l;X\G���<����S��L���3 �/��j���͕g�ki&�Q�&11����ݤ�F��,��=�����R�T�]_��>Qe�;����w�	s�N橁����l[�c������csYVS�|cZ�]�I,�`��]�ŗ�2�Ֆ�٩=����tTj�jS�����}��ڒbl5�QT�I��*���P��;�b�xw}#���~��_zW��x�T؀b����`Q�5,�V�0+��w�@�7�"#v@����g�<��m�qk������H��*/%��X-�\�䃢剶G伬D����%�ݾ[0��/qL_�0٫���2"�|	���H�䅲ĉ�(�e�R�N\&��fpM3��,:陖�P����ѲU�C�M=j{a�mcN���?Zث��=��������c�"�gKt�M��u��n`�1�qQ�@�p�45���_��U{oh��g3�wOΙ_j'r�}3l�r�k���п�V�0�z��;l�:������!���i

�#,�&}�R���q���J�a�������t4l<��lA>��d�k �Nu���/�:�͆&O[��X6�F̜��*I@���E�бJ\	YIH���ᴩ
���P���y
QQ��
�)yt����v�)}(%��-�5�I�t��]�.�v]��k�!w+1bX�"�v"nЦ5]��I�k�^!i�O�I��a���5��r���v��]Lf�_��om�T���mqk��JW(!��32+~�����z�18n�=�B_��ԗj?�)A��8Ѣ��}C��ZyN����(�))��v����g���cI�䶙h�u�yZ|�nim�o�ϲ�B=/'�ʴt'Q9��5/iH�?t����5�wH���y�iC�ȧZ��?�no�$'mG��*�������Q�#�h��܃�/D�aO��6|���a����5����y7�6z�P=�����[���tQl�B~Яw|�;�{HV��\�qwO��]9L�X�����i�t���X���3���8�$fVQYyf)��F.�#Ə.��1�%�O
�I8S���h�#�iN/���w%����{��D#�EЄi����}��.0ǸW�l�&��J2g���LSL��)���V�љK?�m��e�~q�fl��\ژc k�-ך�F��KA��:�����!�rfӼB��M�'�г�c�w�-a'˛PΔ�$?��ɣX��A*��K���G3���ft<��,�O�� ��E�j���0�ϴ�/B��c�m�6|/��T�P�VT;�Ǚ��;��T�՞Y�����a���>�<�\�����Jxܸ+�]M�b˻Ro��>�I�F'����y�i�ٖ��ݻ/ڝ��uq=�(��[r�%YG�i�e��fݔul�>ĕQ��j�Q��n:��>�/�ơ�;!h�Vy���4�h��C��Z��趝�df����M�=Gx�����b^�7=�/m,P��7��x4N�-�A���Q�ȑ@'[���^�Cb��>.ug����w��}����2�msYˮ�e-۶�p��ZƲOZ>�e�v-k�������}]�}=t��yf�����W�J�Z����Ș8��J�ڜt؍v������k�"jҬ J�1D4��'H�|O�<��V���ј��ɯ-f-4�|]yr-�.�n�NF�^����џ��1�t"JI"��ry��&�fQ�BDR���c�ې�@H�Y�g�_��Y����=�Qz��>��r �5י-N�;=#���Ab�l�Ma�'u�+sͦ�9uo$�/�=+��<�-nf�=�E��qVu�S��7w��P��2����bŀ߻$�����_�\碑�0z�7�(K��9�K"���Z@Jz�$��7`�f
,?9gLq[ �1�=?F-i<�N
�0����*D�!K�P����K S��x�(��-�x� l	z����B:��6�hGp�I���\�6�*�t�ŋWؼp�0����p����V#[�����~����w�#���V.M�i�+n��'g�T?v���!H ����-��~��e��n��Z?m{}9�[�X�J
P��"cc�&7��+���U�3*���=�Yi�a�bQ���HːK��i�e_o���ab[�+����H�j�hX�
Zת|7��9�����'N;Fb�.�ї�١:�|�?o��R,\;��#l��/|=��e\ڀ6Ji����Bv�1�1��x�J�����X
��!��W���ڗW�0mG�i���d��Qn�J1��Oo/}�[3���c~�� g��v�l��T������677��ӕV[d:�w��Q,'9��#+FFJ��Ł��v���)��4������֘ؓn@gJ������n�fD�@�ąO-R��w�F�f�)t�~^,&�9{�gi���*�z{�$��	�Y9�`�^.����6)�Γ����/��6�bY���*2�<�M)����A��9��_�,��
�[���*j�HC�8�
�e��ʪє���&8u����w�nnǬ�2=��Q�젘���! ��������4qe���
��JS%Ry���٠�n�	M�E-N^E*��&��9YH� KO�\�5[�dFo��]w;�>W@�`�*�F,� �[/_Z��U���&�b�}P8q����|黂M�t�uK�0�-Z��|��Dg�� P~���pC0��e!j���R"СOW�q9n���,XG����%9����%y�!O�`ȧ.=Y�uߥFB�T���͢][���~��
���v%P��c��F���)zs!�J3b;��/:�����^���|6�i�Q�] Vu^C��v����w�^���v.���\��j-�i"��9�8(��kn� =�p�zE���!yo�7�=3�'z��dm1�I�9Zm맅�����!���%b �5��سf�=�*N�n�B�p�(��з��h����9��goP��&���*I}n������r`��~��r�!��?��¬�G�r��Q,��xɣ���U����FOm�Sȷ˳���N%փ�b���;�����&B��7S��=]DL1#
c,1
�6Ϥ$qc	�/�7�씾������������ڲLkf��������ʈl�'�u�UK;ᤦV�1�3���� |q�!���>§Ί�����j�j��}.�v�g�P%��b��$��nȗA��gE[򋺋�>,�9f���T�����Z��1���?�~+�=���|CL�������'�3�cATIcq��\�vDR�m$������p�KI�!~S-�"��r�G4ם����jiL�^��<ۼA񹸑Y��d�%���C��.g�W�2>����ǢP���lቌE_�g��*>�?�QWJ�"����u�-��|FY�p�I�΄��(����_���]�N�U�<�Hh8�HJ��{�餟�1^�p�:�L1�)���~O�ǁ����h@�:r��|骃~�� �Q\� �� 閽�si�Z./bP&#�">b��U��e�o"�JIΈ�SE�	��+�=&"����eOF�sQ垈�S�:y�9;�ritc:4;{���L���&������[�q\����z��(�;���V|�գG�L������1�sa!	�YAdl�ƍ7�+�䭡����SKm��� ^���T*!˂�����ѓ�r��#���f�&>EذE9�%M�ɕX�<��Y���Gܾ���K�B��+�tH����e�p���:\�
[L ��Q����Z���Nr�h*!&��2��!�u�H�O��ݎ�=���1ߧĞ��P��+��K�	y�3�U6��r���@���������eI�]U�8iւ~������O���[Xw潇`����j���zS���w�h`�aA�X# !;�o�tW�����o��|�J5�J�X��ţ�V�� ��͍�;��\��������@�e�c`>�t���,�:h"��kOQ&�sb��Bv��<\[����|�s����b2xH�O��� $_�!��f�z&�9�%�CՑ�=����*�U�D�X�y�̶I��D��ܲ��<(C�m�ru{����&�z��Y�Z n�M"��-?�F}0�	*���;��m��jk�e�2zu��m���1�'��dLF�$�k��iw�>v���>(����le�(�����N�W�I:�a��}�Zw_����ǳߨ���zզ	Ī��D���&�������i�*���SdL���\6]X3�Y0���:n\�7��Ϩ������=��bׅ�TC��:ji��P�H���lb���� *Ɵ���)уb?&�(E���|x��^�OG���LZYHsl�VBD�P2��|V���[��ǒr�G�M�R8M�$���\�P
�����v�K�}K�-�Hn�NFcGϚ�J�V���37���~��O��N�;�����.5$�+��c!C�BrT&�97��\��iw?DJ�ݨ��>)A��U��+I:E�i��;FH4�&��E��0E��;��[D9�`���T�5�oD��YT�Gq�jM����,�F-%�7bj�+�%ʼ=�ۤ~ޙ���j�_�Y�_�\�	���;��t�P���mἂ0��T��#�\�����GZ�H/��S��!���'�R���1�⻳��������pX��Yk�R�㟗���P�%Ԑ9eM�l���
,� }��N��/���$t]
Bwi��H�~���Ty˼���[���v�B�C��{W���T���X�
[�7f�B�7���3T�d���l M�&�%�gs�UR_8o�Gz}V��]־��$o()��O"��j�-,���yƵR?V�CA�95NgW����D�eک��{_Ʋ��3���#�����kp���ӣ�������+#:5ӓ5ߡ�K�\�T�z���券��X�ɉ����h,����e@��|٧���\�)����2�^Ey��"[�tP�Ӕ�Yt��.T���HT�t_y�U�A�H+��zN�%�^Wy�h��k���],+��N��@GIt��,��m��Q2���cz���i���[��U��ӏ��?�~;�NZ�|q�r���q��	8]# �J�Q��cY��g�������X)'�;���
���Z����b�$��w�hL�)"]k�6������i	D�\I�L:�����1�Tq[� �m��Qc��Z�t!�^�+7��(j3�aU� �ijBK�ŝ���s����1И��C�}��L )+.e�����=,���ji��������\���H�X��r
]8-�u����$�۝��d��,�F<HS����/ͭ�t<��f"��v�^ V-w)�~y$'0WFp��~����0���}k#�ۃ�>��f;��r+��z�i� `�O�|'�(��ff�	�(Ѝ�yjBT^�#: v8Bb�b�;����ʡ���z�)T��Q�?e�H�.��=�$�$u�44|4"zw��!A�.�UeQnRkml]b�`��|M�/��}�
YP�X�#�����c	7-��a��bc}To�����ē��.��� �JUf���s�K���^���X'}�%���w�Ͼ6/�Cs%Q�/ڱ�e�eH��1E(N�m��>��������e��|m�w������xo�o��8/�-띰���4��ÿvo �?�d���VJ�6���t���x.5H�"�@`	�?o�1%���.;5{@�.�L�C�<]E�>'���I8�ޛ� ��%N�P�.M75���[�-|(� �Fؖ�J
,���P���Y�݆���a�f
Q�-��q�����QC���x�1�Z��x9y���~� �Y��F)Em�y��f�QS�ѥO��Ǣ6�7J���u��&f˺��§�;(��g��a+��M�fYwx|���mT�)܅�@F\�B�W�O߈�;�>Z�J���;�a/��R盝�D�T��������Ƒ5޷���'�R��=WA;C��<� R��j�Q�������8#�1�
J�^���!X���n�gtʳ��|NK��mS{�[j>�Jў��`��9�Nn�з��ל����^��X�oԣf�"ڡ0T���� ����A�I1�X_nY��օ�����JX?��dQȕEq(�j���;�d֡�#5�#��*]�&�Ί��iӔ���Tr/�&;�5��L�2=a@�T|Dd5��d��ݼ�����D�%	q���؈~`U��^n)I;�����g��6�R��w��p�3�¨�;��h��7�̈p
���]H�lN/�syy���U����[Ma�@�7R�*�ewZ��yd�~	����������1��X�y��GQr����Z4ָE,�҂����H�p.S���%��@y��ᑨG@5{�d��V��ƴ)R�?M�94��r��u<[��L.�N9!@i���D�#�8n8� �n�T����D�Q�z���??[��R���[~蕩��V#�d�4�6�l����</{Z��"�2Z:N�blB�$l�O�欖�!�MQ�;�u�>$ ��ǳL<��d��'��?=wK����]�[9#��b�a�����p���C�al����\��A�!s�uqD�n���s���͓
��S���n���@�P�#RT�*��dw�3�?�ǈ�p��ׂ���_/�C�-q� �~���'�b�'��C��W��v��n����7'K8\Oi�a@$"�����BaS@V�!������+���s�	`��e���j�|�&o-��5����Ú�Z����^!�G����V��ĸ�����8�{P+{z�K����s���Ŏj���f�G��-��?b�}�Do �Q�v��Q�n��|є1�q� ՛�����X�`�;�ލ����[AKC�(�j���5��K�Bj�~x�j�"}NF[�'KM���<���3��;�.��b�����p�2�ְKP���K�Z'��bI�m7fme�UH�Ylk�4	�S�$#:��m�d�;�aDg�^�SU��fJ�"X��˴ 4���ۛ�D(;��o���#[u�c�(+��K���V?ʈ{!��W#�z���q�)�]�ҥ�(���kt�m�׏ ���M?u�oP<�'��g�
eWg?]�_+1�a?���D�R�Xw���0��	[��2�����q8���_X��2A
�}��%������0ۃZ��U=-�����t��j���v��7�l��K(��reOE���z*�Ez~��E�$����
����c�d�6Y����(�W��q�o��oƿw��y+�o/�pS�X�l�u���(�T*��[�{KW�$��?��8���6�Գpp�T;"YۗJ"�xc�N8Ҳ���L��(��k����_p�cjس�E'�������`���.���ş��TfQ�Z��7�IT�e�k�R���nF	�!��ླ��;�bg6 !��6�>�52��AVa"cMQ�Ѯ�`�D ��I$��9��3�!��Ԕ'�|�=�a�����S��G?��e,M�C�kv���rfA�,]��q�c+Ŋ�+�*h�c�]�#C*<`"�����="DO�?>0��F;QM��2�lP��X�#U�]�W�h�=�Q?���^uf��	-��VGt�r]������򹃨,db�>�J!$G�����e��<��HyS�Όh��Փ��T������i�[͗����?.�����{�Y-��(� p������+Ǘn����L�7y�1t�-y�2 ?"���"��M�
�&e5ŝbqe�5�	�ҩsl<HO�Fq)D���cf������<��#Y�
8�dx�ŝaA��oX�]�e����h�J��zᬒ��.?n�-5{���$�^mݖ30�6)ߛpa����ʀ�L���k�U� J��9#{�I�%�H<�9"��R��=��g�d��S� 7�O(\d�h��D��[�#Y6z3��H��^
��;�vuq4{ߝ2&�RZ�m�"8���i��j���i$5�l.Gq;���0IY�����H�=��H���?^�L�t�r[9��V�AA�I���s�J�i<�P�ԧ��?Bl����^|� j6�F��t_�E��P��|f[�M�H�����wD�-�8�c���i�;n�@�܏-��b���bd^MM��Ld\�1OX5�B��%6�a~^7�H�,z�CN.���dB�.�^�]zVL�w���r���=��vNռ̚�	�t=���B;�X�Ք��! �c��y�S�f��MG`kx�cz�H���L�D��fȵä
%wq�ϵ �˳����mH_s� ���� �9kh9ZQ�"wC�/q �1��/c˜�!�V�����O�ߘ&Wh���u����>bQ�Q�q�]�����dl�#)�AM��v���D�[��Rډ��Z���#ԣ�lc�nw�_��t~�s}[,���x�_����đ�ѻ^�Uő+D��6�'��1���}N痔}�{�܄�;���!^}���cKMv�Έ�)�����L����=L������:Yb��ZT�A�9B������q����	]7���=&T�ޑ>����>�ؔ�[�^�il �K�#�٬�%NF��fA=���[��`����@���{N�n�V�Q�ݶ5㢯�q�\*� �/L0Z	R�F�zoV9��n��ok�M�Z��w�Z"k���F
�N"�����m�<����N\�tr>���=��[�Br.�
��=��L�g$���b��ى��L��a�3�%n��6]�vqA�� S�&Qx��jD
�һeA|�,�;�R�:�j����zJuU�Ka#�	��J�*Upt9'esȸE�}a�Q���t��{[���<��� 1%���A�185�Ǣq���|�o齖g�7��/+�x�-��j磈��'5&�c\��ɗ����E�&I���M�P\�,�M[�����|�cݓ��[뫮� D��T̢h���y}lc�+́�#?��I6�GvW�������&'/�tv=9�K��ueڨ���"�����O��UT����j�$�V�������A�H��u|���� �h��<(:^JO�(��= ���x�M=+�ɿ+j�<;\�P>���e���A�[����:),��fiQ�J������-a
q���#%o	�>쿖75
��0dȍ�$�>HMs���<!4~_L��	���]�ļ�I��p�KS�(�mSp����BM�s�0�����k�/
-xofr��,� S?����G���7g�w�*�i+�����1�`=bJ�۾ۨ�ǧuՐu��+�.��C���z���ZUYkX��,��5����o��Aw�-�i��!�����D�WW�0;�{��Z�W�Rk��.�8�	-��N 	��~&���e!1�Γ�kz5@6C���R�]w�o/krl�q�pB!�W��y�p�oc��1��C�n���n�"�Z���HE�b_����i�!#��f�G!�r��7[���ʀ��ܢ�Gi�o��`2���k�91� ^eok���ܸ�Cb�	}R��~;8t��ø�k�N����œ}����J;#+�>�����.��߻��q����A���2��K�^/\��*%�t9[ٗ ܚ�_���J��=��h�?IOdT�bG���
en�M�	j����\�0vN{�>S�>���~�h�l�O��	X`���s���5^WW�ajs��=���{���o��� �!��Q�ɷ��Y&���Y�BM%O��8��<�3��+[n�`F�+�RF�ȭ�����$�������P��&N�}R�����a��J��]�|s�K�a-�}���T��-ff�!��������;�*2�ߓ�Lo�l��{�F\�0���-���36�N�R&��h?$'�mj�
����X�*�0,��HT��ؕu+N��B&���|�M�s,�}�.5i��cfxD��4_A{���&L����dg�ٓl9{1�{�?�w�(�e���К3�����(<F?�E��B��;Ɲj���-QP�}���8�	B�[�J�?�,���+�3���T�5�E�"8G�B��$PDq,>�=j��w�	�F}9�����'3WȏL�w�!�M���8���y����������z^kN9,�]�[�0hTB4����[������8�:xY�yt���Y'���y�8�ϹU&�4�6��GD��D1�խX�}��BPg;�[znҕ��8�;#������%}��L$���&ڧ"��V�Qi����9t/�T���%#=�Pp{��j��M�x�]9�j�႑����z��̩�M�Rmr� k5G��o4�+#G�fԫ]�X�p.,;4��`�`;�V)lq>#"��@D/� �ܺͧd�c�Z�g`/1F�d��۟��=I}�:L���r-��	��pF��������JH���iƴ鯃�:����72�_��tʯ�c.��*;���T%za�lF��8��j�f����ʽ������[q���h ����S�M�
V{�7*B'Oj/�A�ڙy	Kvc���:B��)	�t����5k��f5oi�r��ߐ�2��\5�Z��UŵO�d�~��\�HY1[���v��4ХrV-H�eB�A�Z��p�,�s5��h[�ї$s�reU.�)����W/��];��YŻ����������m�8��,;M�G�h��2��j�\um\Ȅ�AW"A�^0O;5��^a�"!Pԩ'���-'�OF�
&Ѻ���si�I�$+�z8#|�LB��rٛGϚ�p��G���K�<��3/��l�R�~�/�v��˚�5r2&�ķ}Z`�c�mr�$���;�8FXC<���B�� ���48	�1���pn�\4�@'I'�:�xm���
�I��5�����fE���Pn��VĪ�+Js���NRY2l�{��Q8��1�������(������9+tE��e��t��������g��2��,��_�$¤��".wA1�c1�3����3	S����M<ӭM��ܖ9�E��	�y���j�FP.���׻�Yf�n�y�b�@���,S���&������)'�vW^^���F�Qi�?����� Cf��'�w��%_���w	2�<��*�c	)�qU��mLL�}����N�w:��.�� ��<l���
�q�~��
�0��KY�5c�}o��掆��	;�ߐ��_���U ����X.���pro�vb���*"��f�-�`*��\�"U���I��,H�J���t<b�[#&cSu�>'��8��馐�H�hyqK�4ب�C�r��V����F�֍k�.3��1�\�[l���cL�<����dM~,�;��^&�x�q�Q���_�����	����_x�0�������.�DE��-N��e��
����4&c0�B:W�sm&�c?�	��+9*�C���]I�����y�@ktqW���"�#x��4�Ƞ��Z3]
�{�	���ht7�����:._�jpis0�J|ǥ���?�PӐD1�N�؉��w"���i��v�����\yv���Uf#��K�H�Q|*�B�D#��x��[;n> I��l�c�Q�b����7v�u� o�d8�) HEE��-�S[[]XH��綡+�p
����зJym����-�v�澱I���BG��+a�۝��ݘ�ܧF�*I�u���S5�f�->��wIf��Y{Uu|��	 8��<��/��B��;�ҏ��~�>$2+�O!C�BF�)�g1rƉm[�x���G\�6���Ѿ_^��a����߬��2�$]1g��2,hU�ad�%G4�f'����&��>ߟ̰Q�R�0%Ԃd'��m�����UgpsI-���w�q�v�+���Ƀ�&�X,o���~Zˣ�h��B�Ѭ��;-��4܄~	i�t�ӇEԹ�_�9>QbNj���v��n>x�u1a��hD��"}�_�U�F�]=�o�4X(���
{�e:J���O ޯ��<0uEK	���F�ݥ�;���6�!�����L���.�M!fL�p�/S�@�q_z��E�?��J�-B�HaJe��oe�.�>z1��a�#zNT��$�@C�hlb����i�D��AmCX�MV��1H��9���Ba��<0s�e2�0E�V�$/�[���c/������A�)���V�w��$�|��6�'��Sy���0)�|�����/:#6�~�����{��|<;��>*4�H�=d�#�;i�����~��U2�4(M��d���>!������Io�4=F#�V��٘�bZ3Y=����a�ph�.e܇bu'��cmm�#U���%Z���"�p(V���Ru�.��KٝΜ)�ƅkD%��V׺M�饤�o��<=љ���o/���8�L���k�K�"�rV(��U����1��L�ٷ1��Kvp�}�K	k��3v�~��b<.ɷ�NKɮ�ɝr�� �:��y��R����=��������_�cL�7w_��=$b�<z*�ۘ�w�>`J5�*�k�y 
N�a/A|q�Fu~���4���7�)��!/��(r>b- �"�θ�M~��"�m�5��n��&�$�F�F�/��5���*K*lD�m��Ѹd��n��X�y�� +����'ȴ��%�(@��SM�ᣟ~%Ѷ�@�	�e��@���4Jr�T�����sǜ��@�R.� ��l\.O"6�[��!sy��(�f!�B��2�u��\�Ax_��=7��G`Ō�.�C���~��ˑ~�Ϝ���PZ�����g�֒SDΪp����$O��/ z���D�>*���@�M!E/7X�A03�(���P&q�5%n?��-��#�����U�$��<��U0;Wʙ�q�n %�z�3��e�B�TZc��n��4����B0Y��
��*��A�#��	K�U_ �c�e����J������a*\��&h��ţu�Ҋh�/�����m����)��_U��'����H�?Fe5�a3�&sUE�Ap�"X�H<
,ä��Ǹ�B�㔛�TL����Q��;�2M��I��f47"��w�&:$r)ߜ�Ps�]���[�=Č~�-�h�[�C!f�O[�WI��������d������R�̘�6�;f�ؾ��]����68�W3�qW��+�������D�̏��>nn�A%�ܪ�j�!E/�+����г:D����J���?���Ύ��N;������[\�%g�K�[�S		g8���#�@��&�m�w�����5�	G�R	����ͲiX���n��xF۬e9ն-뀃�!\�3�<%�!c]�I����(A7D+l� k�����g�F�bE�!��zņl�kk�TpC��d3�odY�	a-6?��>��(q����Yn^EvnU���$9c�q���y���id ��l11�6��e�ǯ ��+}��~s�Q\�'���*�fF��5c�����6��B�0<�0���ި&����MA�,7�0`:���˸t f
�	J���I'�I�_i�/u�?�X�O�_hL	�&�H�~Ԡʝ�s�V�� q�<F�(�;��S�)]P?&ΐ}��?��R}S����嚝X�b��}��
�ȂVP�vO ����@'ogaѹ����A�f`%�(nx2u=��L��R� ���vo�gЯ��ҋKA�E��Υ�C235��m	�*G���Z���W|��j��h�9$��ؒ7xH����CT��F:_���J'ibp$ns�{���Κ�\P6R#�*�XT����R�X�ܟiO_}�0P�i�X珣�\r��'1D�W����2�0t�ԑ8���i#&� ���4�%��1�U�4����-���
z5>ڔ�jJ%c�Y/gR�d˱F���������%��)�\�6�'����2i=�*��G����ȧf?������dz�X�j�İt$�Wia���1��l�|���4+�]e��
�lE"ω���ߤ�[��c�%��B�L�Gk��A4g,�f�9���O���[���,R(t�,���zHlDj��4CYVΙ|��T4>,&�<�jKa�˫J>gG��GDֈd�X���;�)�#��{�%:�F�CP���]�g �~�e�\�y&�PB��&���B�[U�1c1�ڌ2#ԃ�Z�ow�I�z�Ɯ3��,T	�w��O�-�L7��h��,R-2"�>��Ȅ9���
=�*oT�K��찒:c��k�5��SN�w��o{���;��
z<�u�k���(T+���<���]H��:��+�p�C�C����>�c��c͇E��9�y0��P�{�[�.>޸CK���X�]Vf��i�ߠ�3]H�rO�ˈ�t:�z�5衡��E��z�|�.s��w�6�p�	b�i9*���
97u076��P=��qի�c�e�I<z=Y=��'N�t��]�v���N���e����xf$jH�<�yVA�碛*O�����ǻ.^�*�7`x��$r��铧��2b�&O����Mm���Q���tV���
=u#���-é��N¹̇�D�����_yՀ*!�6�������Cz�[�������k�$Vi�+�|��f޼vO<[�ѹq��`���`��i<~5���%]�����������2�b�
d5^�.���l����ľ02;�A�������[���L$Q�+<�+�?n���6�I�d�+����$r�{j!;�~W��v��#�֒��Y �x�F�G�f�O�d#"s'�ޘ�-.��A_P@}����.��O ,��l�v��2�T��J G�Kj�����H� u��Fne�y�e�dj#����^�n���;�.쩮���/3�@�Hm�Z��p�E�?x�4-)�l�4@�$�Q2�H�WT�j�+<j�[��@%aڲ��m��b��c�Ϣ�k�s�9�z�^jE�P��R�c����1>�d�u�I�Gj���Խ��_�e�^>�%�kD<��iA�EJ^����xP:8𳲓`yc�A����1o�q���zC�Jm��� �[r��Tl~D���3�oS�[AG�_�2->(��0/o����B� �a�*QT�ϓB�R?Rr&�x	��B�d���@���.��è��G�p���V��.��r %�0*T���.W�^C�����jEݒ�Ks�+�C�m18����{���;��-H?�ڕ���߳�%/e�x����E��a$���=���k�Ҭ�V�ԄO�����}U����l�<�}Y}�'��*&�*�O��>80(v�^����@T?�L�����c !��sQ�tJ4|����jc` ͑q��K�arwmƒ��§�K]8��k�.��MC��?|%{#Z�������GVV��h�T��|������!I���w$�^o�K�:�˽�a���ɝ<i�c-��q1�ë£��9z�WB�7S�&��H����G	[y
py�8�N�c�	e�7�&N:bӖ�'N�@}G���\);:�_?yW�pr�ǤH9E�K?�Z^]�\}��͋MT�&)��U�2���x�Apۯ��?7#y���������k��7��Xf���O=L�J%�S�w�Ȕ����*��O��U@RZ�t�
M�L����*\=��d��c�t��K�v'Y]��u�PЕ��1c2jR����8Q���6��l��N��H���)�I���s���Yʵ�<9����݄c5AUq~��5{Q�(	���Ec['.�hI�S븓\���=b�-�9�F�ũz��h�
���{q˖Ė�1�hF�����k��2�Yw��vݎ�����@Wu��̹dlk�r=�=��nV$��c<��˝�Q��\�]	tF:�E���[�yS�2�?*��K)���%n�%�'N-��|�����-X����M�"���RQ(������|-��[�s� 6������j�����"�>���^��+_�T-;p�"B'=2S\�Xl�U���x�X��>b��jQ�4b���B�1���$�3C�c�ͮ2{�'e���N������2^,�?��B���y�p,�Ԁe.{TiIN_6�W��cW^��OWo���}�'���nMߞ5Cւ�|(|�{H��� �^^;�tqxA�Z�|*�D�*1x�u��L�xf!d��\�OKע9ހ���襂��\�+l��Qf�`�䃋���~��-��Xo�9�>���4�o+g�]�<F�G��U00d���i&#�����\�@��p� ��n�U=>�Q7}��K���\}�rO�<B�#4��*�/�Bsq٩�: H�R>��#Kաxc�� ��p�2�tk����F�8WU*N�M����>���eFw��������i2�=��W�F@�g)��V|zl.[�I��aL:$S[�=)��*�3�j47��|{��)�49 xtfm�S��p�K �<VC
y��O������"�*d���9�mR�$L���?tYdj�����g\�N�v���P{f�<hkF�,�[�}~>4y�o'��G	�d��������9?`K�ч]��Zr1�*�1$�p/u�� H�HK�ިǀ��H��1o��.�P}��W���y��k0�,썿M��k�ݮ��r��C<��*p%�J�;X�t���w���Y�m_m�6u������s�(Sq��,�DxY���ė˒��8+�nDym�g~
�Ꞌ������Rc�W�!�� -���h�M+I���1�������0�}v��N5��K8��3�Y�T%��6�4
`o���A�g��,�7�y�z��)�j-#sD3�-:���~a��lkfO�ڲn�.3�����O1�]����P.��]IF��/0Zۃ,N�$t�L&B�U�|8'�Q���Uv���,�a��)J�O��0��ǥ�aX�)��>놁W��z������s�W?o)pl.�)Ȃ�dU�����S�8���&zŗ����Usk��{�I=�v��yq/s˅̏v
d��O�Ϗ�#���3ڲH7�N�8y}e��:.�R�،i�C�E
S4&�i�P���A������_�trW۱c���(ZC�%e���RxtK8$jG;�X­��q�a��[�jq�J����U��s�!���'�q��W�����9m�+��[�qx��q�[���_����L�|��"兺bKx�)�lοO��&�Eq���9��:��^_���\66�$������R�s����3\�����d�Z���/'~�+�	���'c�c�|[cj/|Bh�L�f� ��o�ё�������n��D���CXGo���%�kk�*/��(��t<�5+
=�lmb �H�,�V��jp7`Do��Z׹i�qڊ����޲�O��g�s+dJ����g�B�8Y��-}������i�8_�����j�lm����%ֲ�D�<�0�!���Sۊ�C�0����$���":fD�MH
<�=(W$Z_����|N6�[��|K$����熄�L�~ܢ+�G�pe��~z�Iw�$Um���Yl����ĞQ�0gL���dij��A�A�C����q�;g�����JVSՏz��`�x$�D�8]�!:4	�,tQD��J<��P�Mr��~�5#T�ac'\�{ƜX���ߔE�"�9�śoi����>�Z��,��%�8:���>�F��h��.��N�l]pk��3I�k^�0��#i�5�+p��R�ʅ/��!��!�Bk����g����cϯ�w�MWl�i���.zkbn��J��'k�g���.]�����_�����S��7ľ�У#j�	�>������#����U.��E��vf��Tx/���s:�9�͆F#����8�ݷ����]��w�>(1H7R-F|�Y�>�	�5!c��*|�-EPI�M�f�9����EކJ�lX�iM�?�!�"=kV{-���1�lM��ڊ� HJI��(�0�D����hƐ.�!  -a�]�����h$65����y��#��|��jw5��݃sG�&�Fxa���|Y�OpppSK�z ^4����w���^��C>_.i¸�'Y���a2��M�J�3RƟ
lʢ.���Kw>��E�}@�eK�8a
���=jo�P��β������[N�.W��I<0����-�o�S�nw]?��oN��Qa�$ѵ �z�CM�c=�橝�C�?�l������x��XdBuF��dO� ���ʮ��S����2mB�1��z!{�9�<�U,f�ry�Gmn�����=pv��ҡ&�ZZ�!03r����^�}`�I$��|7�,�������adav@�����,q�b�I�Q�9��!��i0�&����3�T|���֪,�(l(�a�׷���Z6W�c2~�\v��<�uN�P�m3�P��x���.^��-�R��p������(���$�<G31���}�wX�������d�[�w��Ye\]�:;�Ǘ�&|R��R���$��<^|�eVmo\�v
@=}�CkR 7q�� 4��y<� F!���[��ǀ��Mטg�u��A���+��&;~`���B:��������{���D�3,+���/�lY�k���O>2j8���jfM>��"Ʀ���}\|7�~`����o��صJ�T�����v&���P��!�#���[��L�m�;���E�׊h�^/_L�z{�l����JW7�h�П�}A�ɬ�8QABuD�#���wj?$jgrO�88�k��]�E6��zہ�{�v�N�[A��� ,�����.�����a:��8T����[k���/��������,���|�D5t�;������5ʸ�8����O4U�hv���O���O��ws�ӛG����~��r�Tc�U�ˇ�����EM���1�W��1�p0��_]=���bB���ǆE5ޅk!��8���So�8&?Bet��-g}���B�Y�7(���k���G8'�Hz���`1�|��T�N.���"���=l��U�U�ev���튒m�U���D���&ۘN��~�y�P�0f3n��K��O�w��=H=ۡUq��L�5ʞO��|Ap|�;!lqѴ4��d���1�'H�'�f}�Bј1��ΏB���M��
T�%�}z6䞧��Z$Ľ�>D8���1���Eo|Y٥X�(����-3auC�?O&]�F�z������?��OL�A}���%��4��w����uͯ��1�)�hSM�ɧT�詤�!���H]�w���nݐ�����$y=�3b��6.�:ﰛ��	���]���,�"�"���J/[��z~#����Z+><!(e�g'�_�">�\w��fY�s=N�,;��OqkT�ED������*/-�>R�:��������'��||��n�D�%����W��%��{�1�Ӻǋ6e2����u�'�xR�#����F�OM�0)���FɺM2֌�H��2��υ=8@	{��S���,���t�ƗO��/q�c��y�(�꨿9̋��;�Ox�Ƕ[8���z��~-;�A���u��Ȇ�x���_�2���:�W���߶�]�
_�a>g���=&���!¹�a��=j%�
��Xch5�q�;�����}ZZB�A�U��W��4�ǟ��X��s("e�1��Z�g��R�fj	����xܢ�	Y�=n��{�Q<�Ř?w^�����Y�vꌝ���Xԕ"߲��>Z��X����םi^4g_%#��������X����n���t�.l����W���tW4y���8v�ˊk��&|�:6Q��8Fυ[V�|��Z��H]�o���~>�ѩ�>j�������'AWV�h��	o���Y�N�	D�������
[���2{��n�]�	կ�Rg����>`�l�,Ռ-U3���/�V���x�L.l��ڭf��
�8�V�"��M��`r��|�{|��)4�����G�g@V���Rv�d�ͩ" Rr�ѵ�'f��%%ER���tm�����f���Tφ'�Ȱ?�.���yQ��ه�V�(Wc�Ei�dD��+���j>� v*��W��x�R��3��/��zc���`�L�g4�Am�3�;Ǳ�w+#ьx.ɯtMQI��ǎ$���_ĉg�{cǸ�Tn,��_ӎͻܱ?<�������@�ٌ���4
�Bg�c��lytl�봞@�~`A3�2��ZhY�	�=v��X	�Dw.�[��{#�ʫ�����RR��%��|:�J08��8hg�y}E6��[���xU7׋�XX�Fժ�q]G�%N+��UB���lڙ{��[՛؟K���e��K�痹H����9j�zV�M(b�h�f���� ��;��-0`C���`0�p㴃䳗�c"ߩ�زG�_�2�kk[ھ)�n�O*�]��������5�͹&/�&��[��"d٦x����m� ԃ[KUC��W4���ڻ#8NL��"�|��s����`���H�OCθ��Tț�;iiK��Z����ב�ф	�Jae���ڶ��,�J��Dk�w�[�-l;�1��/Z�r�rߑ���c��ۓ#������)�yG���4p���K��U/�`ٯ�	�y��84��w�>|cgV��4f(��������f����iF��<'kN+'�a�U9&���eI�_�(|��N�I�_Ϣ��k,>*��A��)���
�A*HJ��g����9F��R���и�X�9�ܟ��!�d�Ki�V��d�CM�"�ل5��%��z�W�&�n���f��PUv3u����SKh��������}����R6����@�o"��S7��ν��=�DJ��W˜��X��:H�3�<�<���o��$��q�ozR�H���s=�?{=N�S�}�Ѽ�~cGUy]8�A�A���-zD�/P:rz�ί)��%Tи{H�������d�1����Љ�P��ԧ�=?c�����'������7��G����<,D�9����,ܛ)Qu�7��s��/�7�gl�?�dss�!�?�Y����2�)&2jKsF�{L!q�����Ј�6�����3.%�`�D��X��.h���Y_1�β�#ǌR�~��TA�	��������!�C�$�J��y����za_R�#E�b�-�c���ߚ׌�l�fӛ���Z�+?6�a�/g����Y��cETx���9F
'd�|њI��/��M�mK+�[�"����>����{�_K�UT.L��]q���O��Oծ�qa����Y�꫾W��f�}��O뙚��+B$�f<9��4��Z��r�LFO�7��9R��7�G0��ϔ�ޏ��F��_�����>��x�h}"1��$s�|��s��fׄd
=�ޙ��DWr�P��V�`TE�%�ޚS"?l�>�'�K����K���X�M���C�v|�e=��e���ʦN
,�z���#D�>+<]�Z���>"��D=>�hb�P�'�m����%���NI��>��-�ϣ�y�����9�jN#��$~���6��C�y�nT�
1�	:\���2��ޘ�s���k&&&��k c�e���i6f��߅�z��f_�M^*}�H��^�A-�G;/���p�뢓�9�ݑ�i��(W?F���-Y�� �mC���(F�qL(���}��_�I'?h�#��'��^�o�cY=���{VgB�=����v�hQ�r� 8^~�W�3ZM���q!���>r���V�^�z��{�7wk���B���uA���A=h�*������5�C#l���r:�����l�����.�X~�m ,P:$�C344���ixI1�W�&�w�:em�Aƪ<n��1J��B��%��֣�A�r{wS��",ﳓ�x�=Ds}�xn������i�#ioG��U��a�u��"�x&zھ?t~HN�(��gן�:�y�d?�ȇE��ڝB��P�O�U iI}�Wp>��j�Whk�Α�#��C��L��(v�+�������1�F����G��������l�zy�wt�f��Y�d�ɩ�s\؅қ���I�K~d:.І��/���X�NK�˕V�*ʮ*e�7�F�;n_)�6�_�����&U1M�Lx͏Π�������\w��B����p����}���� _29~�.➧�9>s�Ys"�v/b�3,e_Wع?R�o�'�hezB/�� R1i�s�|У;(�FתٌX��̽�^6Y �ޭgk6�x�����ZC�/_&���Z	�k�i-~�~c�N�v�k�R	H$���Z{��+*�G�����蝀x5v�Z�U@5�GL����K�oE�?�������&J倃IK�Y���}(d��%_���^�`&7��b�A�D�L?1�OT�]8'A�n�+nr�tS*�_��T�l���������7�FC|6Q�������U�\��pN�X��Ӂ(T6P}}a$�_x~ �i�Ғ�H��g�1����֗�k䓷�hu��R;�4_'5������:/�עo��I��L0u����r �vr��" Y���8dߪ�/�v�|=�-��*�E1U͌8j�y���~� ��/p����������~,	0�
�PY}N�t�����i��3f2�b���!�"֣4٭v�duP`-�\�?R�r �C¸�ФT3o����gs���� s?�6����X�;>4��Bv8���:��~�1�t�s�ȍ>�cI�᪩_n!��)(NمX{��S�I��JeQ�<#��~Hi�;S[G�eO�.��1L(V%��q6�� С;�4��Чjx��D��(8�GO��}[VJZ�(+�u�>�|�1 �{���,�nQk�Pz.˟�y�JVwMr48;o���5�_g���A�'�W�+���5�^3jz�M�ba��V�q�~d�+l�n��}WЯ�cSb���㪡73n�}}�)�~�����?�_6��m��y�����n"���b)�>��-5U<	��yd���Z��	��x+^���yб3rq��f�>�~�uD�軃�#�����PyFX�>m��|�@���5�E�IO5�%�v�]�.�F\C��j�u������fN�S̤e�Jp�f�Y}��zv��X�rӇ�����`F	a,i4vZ(Ui��G
:�yH��8�Թ��G�h5T�3�㴹����4��n����WWIK�+����>�sǣ��R�<r�FYeNBr��4Fd|��"�)���M�%�>���x.F��0��:BWXu����M��V�CE�>�_�����:1�g'�0]x��pa�N���R^�U<��'�6���{)%S�{�'�K`�V������|��aъUoWr����fO,�X��|aϼ �n021	ܾ�[�wBb����~z��J���"A� Z aR
k���JX���Q�s_^�}>�Dk�
�ݾb�\�`7[wj�%�4ݱ"��h�	MG���'�ݰ`�L[kD`C?�V��Z?�&�y3� {����\��?R=b�Q&�9��cB�Q�Q)#䷯�|1��ߦ��N[ LL�!WE`�"!�f@\8�|���S��;��+]&A�x��8�B;��`��y�|�<��<�&T�s�V���c����/P���| ��<�O�,��uw�#z���eM㫩5�hQ2�Y � ��w����l���sfR7���Zb��x�}�ԭ�_�9�������O���2�'	h4#�n�j�R��!y跜A�V��̸���p��0`C����]̝#Ӝ;V�*��k*љ;s�q�R0�FL�|m�=s�V[��;GK�H��8o�Vɯ� =p��K��*�M0wilm��Ї�^�,_֕�RI�o�Hzub�<΄�L3���6]ɼ7>���(�?X��Tu>_�Lc���n�$_��C����}�u��[�e ߒD��w��fX�Y�@3*'��b�c�ט{���0�Ye�X��*��I���ǊV�V�Fv���~��5ꛬ�y�����W�ZW��0�D�ksAq�!�s��#�VI��������iJ�J~Vyky�6Y� �M�V;l���I���H�}.�p 薠g�+���9��6�C^hO<WQ��y�e�6�}�E��濃�?g������k�a&�G�!�ᣛ��f	��}|�yn��G���л�q�'��*����~���yc�Hg[�(�P�5�
wV���{�ڦD@���W �a������/}���W�sx���h��U���)�����V���j�o��Y�%��{��1���Ί�FV>b�NWDk�˶䜍a�:*y����X��v6vԨN���P��L�ν��'�=�/���i����;b1�&�4U/9����D��_������)]|?��&�BO[7>����33��m$����=����f���-��m��.7 ��� ��Ӎ]`^�Ó��_I�z�&����2�����V�aa��.�K1@�|=�}"�~�k8��Q7U�></��Ī�p�{%G~x��c{��z=�3&�8(fq�:^~���a��ڮ�-i��T+0������M�[g���'�тe,��_������tS�QN��a�1���N�34?$���P~��)�X��K����+5�HK����2�>�_6��Nt�,D�z|�k|��h�
�{�+M)�K����:�.��G��S�?��(�hը��0U�<i�Î����Z	��w�	'(�˞68]o߫,K�$0 g�g��5g$�#�GwA� ��Wd�Ț| �\ϗ�t�ζ��]#W-�?��c���\�{��K~��?md�h��*������ᢠ�c߸8.������|t҅M����0"r�3�{9M���W	�������1�&v�pK�c�E�>1V�׹��>�z˚��t��%�âv���Բ�ğ1����׺��PT�|��!p�//�-v�U|����O2~��v�,n y�FUQ���q�I���%ݡ)@��m���?4���ޮ�V�����\v�*<�C߽x�j����z������V�<<��}F��ǽ��yz�O����4�⑅L4�MLڬ�[N�iG�:"��y[T;	���~�8��gmӼb/��)�;F�St�𔐍6�i�
_��qZ=�����:��'��a��J��*��q�qo���h�P�{T���:6/��~ś<��hX5^i�OԼ��+��.�',��mn� �0��^q)�M�p򇑊��*T�+2y�5 ju�v+پ��������޲�]����F,5�┴�C�}[M�H�-��Y�cV��(�r��\��bu$�C�6�p5`@�y�}G:_�!�x�G`	+�;���eho�d����W�I�i��*����zq��ݨ�֌�}H���=�) �����#�>� �݉^�Q�J��C��a�d(�:+3e8�d!X��o!�ŷ�#ˀ�I�a�ո̥�1�X�[��-;[Ml��hg�^<E�<[���s��r���:�R��C{^�b=8���:�V�˲D�6���S�w67���ܪ����ui�LG��'8����=1"�U$��I��@=��-��4��P9�_����Сa��LZL����o�nm)���z	#�����HXl�/�o}�P�{1E������vF��Y�'� �:��վ�qJ���������q�8O�k*�tx=�o/���~n�+���޿�H쓘B�Lu�nݤkb;$�*�� C�*d��.\i�}�±�[�<��"'{��;A{�'Ҵ���N�� ��kJ
������Yrp�]nٞ�>�DzH�����ć�£��F6ol�pt=�i��+g����Fdoh�j�.���{3`{��L���߲~��a��� m�i�+����Q�W܊C�f���}�����M�?n�я�,���|�1�#~SQ�p̻�����h3W�lN��_G"N���8:����\�6���iy(�.|0&�a�q�$`�{cA�I^��"��b�^�t#C)��(�E�vU��9�YZ����"a�-4���tW �X������)�BĒ	#Ґ A������SHR�Zc'��1�f��'A��n���7ݼ1b�6�v�#í��i��?�$khs�ιV�dg���hL�
`bn���V�-Y�3vN�jȣ�/{�P����c��x��-!R���a �@����ȭ."�� s��z��.��5O�7]+2�)g jRꛢ�۷Q<دt|����\=�������y���u��-:�p' �3�t�"�Ӥ��,���^�O(�I�
T��E��G�|����E��Y.X��c���p�SA]ݢ_�Fs�:y8�5~�*[u$������*9o���-��}��8X`��8:�<�c���M����8�}����M�;p�{���0�Yf�7Q�vc�;�R��>���g��N����OJ]��*���b�ɵLuW�{Ya�ىL�E�<�6e�66�	p���:|���"W��W�s �,������2�T�\�u�jI6��r� (^xt<�UFD��XkU�X��ό;�F�m���oǋ�����`;L�VCZ���Y��������j;���Iӧ�E�[&���0+*���G��u���V�fJ�#.�#�8��������k��'���b^Yq�@�Ԍ����|�G������S	6RYi!Cpu��w	��~�Vd)I��0#Ǌ�T�عz� 8���@T*������񄩎�Ǌo��eL�M�B���e����.�=3v7�aN",�!,`ڕr.���z�9���i�K �����1q�ނ�J��|ͮY������^N�)�9��Ocn[�}�ɤ�������z�=�w�Ί�_AV�K_D����P�U�|2���\~�\]��*�ӳ�I����~�"�'X���~����T�����>�I����Qw��,�v҅���*8�!.8V�P�<�����í�K�h�x&*SΔ~�{��H��9����[��v �t����Dc�������F9p����^zE�`��β���|�O�K��$��x����Kը���Sj��JDZU�>��{�2�	Y?-Tg
��`�W�0h�|v��$)�%12m�,�r%��&C+^/Ky�cJL�]0i�+�מ�O&r�+4�y	�R0���yT����9�?U>fS�i�MUU�����qt�������ONX�_R�N>
6Z� ߠ��)��S��m,���K�*�z�u�8A�-��;���N�sj�����%Q��"�b^p��o]�ԘB�o�� ���3B�]�����%������`�re�2�kG3�����|�D����7�����!u�WH�k�;{�p]���ӫ�~��de��v�s�EC�Q5ν�uC�e�?=~�?��4�V�l'�h�t:�pFA�fU����ܧ߷�6�F�w��À�l�Xk�Vw�lp3ɘ�V���n	����B������g�y�j���/�|�	��\�`�y�I�3��oV,<�I*����?v�t��Ol)��:�����,u�9y���]V� Jr�������7�U�)�����R��ؕg��ќK��Y�����2�[�������V�#��L��<0%'�,�
L�b�M��_�j�|^��X�ߩ%�/��d��yڱ�5q����4_��N&NЋh�1Kdu�.Zl��{t�1���9lL��a\gI��8"m"����qі2�0���u���4E���s�&�%�`#WJ�Vت
�^�{�x�0.��;���+�<$�UG1L��SK8��$S4"���-eD�اp��9��.̂<fAX�  �~����l��3������)D�ڦ��&���y�jsw[xM��9[�� ��"ކ��SG��6�NQ�'�Ң�f��3��w�	�Lz��2"��V��Ms�Z��~�S	K�A ��� ���7l�0#o֮#�����X/j+:�$�w��]�5䞢	��7c����6Z�lϏ?
~V�i�Q��[�0�ֹv����{$&1�⑲~ i��As�^�9zs����h�Y�#�o�{�������f6~6�s�aE��=;*���6�F����'b��I֬���.pD���b� �vOƷO���!�Z���	��=� E�f;�5���
�uȾ�!��R��<��0�w�[�;S�� �б<��w�e��x��K5�����y�S���N&��Ƞq�sG��$���_��5���k}�e���:�@s��ʝ����z��cDG����m �&�D ��L���I�_��^g��  �HA��~+▅����k�}�^ �z@5��u̍���<���{����)o7�:�9�@���?hZ5M����%%]��-Uƃ�7Z��;�g�=�3>x �j9�.���9&O�-��}���j˕3�g�4 ߈Dl�r���ʕ�ճK��6�T�e��R�D!���q��H\��w��J�<᳕�u4�~�o���f�BP�൪X�����)G�'���Ľă��K�.{�#m����,�P�B�X4�о'!��*H�R�j҆��u���o�|���W�7���So�C�~����T��7�E��iYE����__���Z'�l���=�DV��������uq�G��5R��'�sEqp��S����BO�D��o[���8!Y	"�}"�b_jp~SK~�]�EX@����K�m�_C\�6rx-f<�;j�
�'��I=jִk�23�|�OMv{9'��B�]�K)�+ÏQo�'O�e>��E=��ZxVqt���X������e�c��U��~h6j	�~"]��;��9#QML��)��<�*�z�O~�olSUNu��n�_�����i�n��/&}}��k��s���F�|,��\A+����p���{�y���j���h��f��Y�h�{�î�����7xK:�?"���q$_7����l)����]=����g��C�y��xr���Y�d҅�Q��F�ƾ�z�����o
yBkÝ�9ĉ̺���,
�"�-(|��W�����q�' ���+Q
�x	x��䃬�~h܎B}�`,YJR���g$g6Rʽ�
?�9��,x���]�c.���)3���ب2kS�!��4��B�,�2��9�p�{�уi9,�����4�1�12�� �v �@*ّ�Z(������=��a[��}����C눏I��}��T�&���![���4���{
���j�a~�IN���P$�����������͎����ӝUcJ{#C���8(3vY�I�n����Lu��ͯ�g�h��r_���Κ2���ڤ��a�!�([��fg���W`��G\��ٯ��N�jB��򣍟#�ke^u��	�!����i�BG�oe���_�$�1>�@�r��2�q� s����B���� �� �#�KY_;�;{��G�a���0/��lY��[�̸��}��ג|�+��9݊��GC��g[q�1�D�]���>�|=�9����p��.+���I�q(-0c%if��#}��蘾�@3�K�����!d'vu]	���[��(C>?�5GַȪ�9�\z6��
v=�	�?��˙;6Y$/(����U	�ց���G(�}� (�R�����RȤQ׺�Ab�����-�����u�Łq���0ʧ*gj#�'����7�`q�Cq����7H���s#M�� '�X�����}	�7־!��>��m1���8��A��r]��D�����}vù2�9]UU�RT!���/�pk5��:��w%�ʣ�>35 �yz��q����4�ܼ%T�>�qQ?02�5�y��������9K_��2�;�}���]V���<�A�}��~f�!�S��:���Sv�r�6��
�hahI�r�-p��a/?�<��vX�&K�:d��<+Ёx��Cv����f~�������lN@vҏ��<�m<�f���؁�х�������ͷ��DU��q�[T�R�V�S.A�q[��<�n.�s�N/[���,�܀�(�
x�ek���ٲ�+M�R`��v��5�F6ׇ�u��"���Ͱ����W��'���wL�F��Z�qpV��#1���˯��%zX�N��,lG=�㙋z��Մ=
*ψ�_����2N"�[�;�⮳?+����ç5h�@?�����M(!Q��e��XZl`�`�2	 ��|��zH���z!Fk9�'�:����kg�*��3�2���[�����p��^�Uy ��?����s�7��]X�� Yw�m��ſ�z�,��������֔�r��@}�s��@�|�����.T��z}�U{�s+f�a�𬴽�.J�֠ILV�WviR��)��C�Y���R��Fw.ۙE�>[�R����ɪ�_����xƑ����ekP�=ⳋ������rB`,�K�\Ru���'�Ń���ʕS&��8�
�Z���a%ʥT��ܶ�N�Wr�pszH˭����|(O�?	O��a2
�2�p �����˪�~�@D�η��App\��9�^8�FtìD���l����]h������
�WN����L��R��o��L}��|�to ��_�����r�=/�����d����y�
���w'
-؏8Wzf�Ǿ�踫������	�֣<͑X	��n=��Zaj�s�C�`ooF��>ד冼م����n��+�7aPB��aN"�7�!$�	n�b�Pd�T�#����ARI�o���$���8S2l����fM��;��UjG�hL��K8r�v��� swm���I����pZi�4B~p���4�A�/xf�������u����2�N>��j�e������Ԕ�o�M�u"�8Dh��2��XddS��UQ��5J��SӸS�9z�G2�y^�ih���bW�{pgK>���Z&��
Ж�lA��kn��k*��/Jdvrb�mdP|<o3�﯏��(Ѽ���/t��C�}y����W��l���[,��C�����G4��'I�����0	`ekSd�AԌ����	}+�)��ꡆ�r�Νr8O����[r�8�x�rUq��@�D����A���j�aU�̹�w:0��mf�Rh����̲m,�ذ���ܴk�I���!�L>�tL���щ�e\�8g���Vʂ~!L�A�ҹD�=s��%�Ef���(+~��E���~1�p�ݭ�<���b�||.L�'�:oN��A���u�����<��)��N�w���鞓��͒�����͵�d�ƈ8���D�.b��n-:�am'+qo����Vs%A>��ig 	h��)�2��'��F�J7E_ʓ$Ɇ���t��@���M�A�e�T�.����"��!K��$��qx�'d IXO�se�i�j�[0�o�����$���
�w�#f6M^n=�+��|[��b�ƥB�J�Gc��`���\6��O��W��) �E��h���L��J=�5�tǿ���z�&��AeC!D�@�����i��)��_в���ʊ�/�`$�:�5���� ���c���[�g��7^_pj���]���~�<���T�#����@ROq4�QWh�G��H�YF�xh����i�p�����O��*�I~/~�e�ctP��d�m�⦜�=���d�EZJTĨ�5Na�94A���S�����Ӂ~��
#�0���vD�V3hZ0���h���k7��Dz�4Kt&��`h��d�t��ʠIJ�@PY ���60p6���Σe1����'^�󎳿U �8͉S^�m<�gu���j�ɤ(5�������Y��
���%r4U�HԎT/o���(2�6�������A���j�����x�׿纶f�x�� ��\q��D�Jb�_�셭�k
{v�%��0���N�#�y�"�����Lq܍!�R��)>r"+C�S��Џ�j ��G�hͅ{Rx�����&1�ƾ9�
X�3�ޥ�m�URe�r�G#�$���v(�ZY�N�N��==/g��4uל����>t3�.��w=?h���e�p�Y<iZ�c8��,c�=	7�^.�@J������X6|iýDT�R�X���7/����������:.������,�eY]��;�2�ʷ��2.����I�9T�_O��n;{zmJ�����ZD�Y�b�A����G��o�������(54��q7c���Vt)�%m�����������E��V���V����_)m\u.#j{�`��=䴜�55�a�q����?K"_L״�8���ʂ�"@�^8�Iy��ΜpXn��*����L�����^^�{�c�y_:s_u�����Z��B��K�ӫ�Ym��!� �p�=o������^g`����"�Z�k��U�X:@���Red��#���J�aJ:�0n"]�Nbo��c~���-��a�XtC��@��[0�5�ʵ5
�;�$��Sv�C�Iu��R��#*(�A��/De�<\����jP����n��~����xGӢ����F���FF;����Px�=[8Ϣ�z�zHb�U�#·̕_S�X��fQ3o`-��ǁ�ͷґ����7&ݴ��D<d�++�ul�Y�͆-b�c�D�Y#_����\*�!�6�R5�?3J�e��ޘ�Z{s�еꫤi^�zs������ѵ��'�W��C��E"9����������������s�C����b�j\w�U�O��M����;��o)Z�-��{����	��{����%V��K�]��xPЩC�	I�ۜ��{bzv|v��v)G��KG�-^I�[��.������g�ݟ��SuJ���J�׬�.<�ֶ~��/������|=7����t�����,�u��8������`Q�.���d�z��x#����tQ��%}H�a7�fhл�~js E�6�@����⦒>���R���J�7�vT����]xIf�UX�Z�s���B����:�����õ�=�HjN�P�Ú�a�����#�9�{�/A���̙;���9&���ڋΘb��L���1<]�)��W��J�c"�:�+8Ď��{4�#�]��umo�W���V)N}^
t������<Ty��N�8P9H�e�7�)�����hhLu��*Llz����F��ҧ�uVo��uS��Yڪ�嗿W�I��b�w+'����8�U�Un'��#�đ������vHhT
�5
l�Ζ���}T�z��(���t�A�0��:��ϋ/����vJ�6^�m�y� ��ޝ�6z*{2?h�HQ���E���&�������a>GǇ�8Zu�J�%Xu��\ԣ��x��˘u�@|���x4�}�>��qkā!�7h+l��BT��#���`@-�ga�����U_{����3��vw[74a�ӿB�XY��ёK�˱��G���<���=�k���.wWذw�O��wno�Dq�[}�lr~���e�>�/��>5�.}jܿN[.�� >��c�}V��Ìᮯ�eps^�k[ȠT�d���4ml�O����m�-�vL������*���������N�n)�G�j�O��J�+�d���B&�^�.��loy�9=ƇI��i��f���W�"
����#Ńȸ�'��c0_��00��qNsb�L�cW#|�����ʢX2�ޣD�"ާ�qA�$�3,zj���[�n�E,
��Y�>ͭ��|�;����[u�2i���$�֙f���R�R��П]�w�kd�.��ղF�Y=�g����4��-1�'#�D�=sc��'?O!>�$fV=�I8*B9��<��w|���t#oܦ�s�T92�}�/t,��ˇ��;�}O`�F���|~u�[`���]_�ZB-iiބ�����?�L��<B�Cl��e9"V�2�U�\F;�bz�	(?
�e�Q�+Q�=M#�Z�'������O��9�*}�h�ӄ�������F�Π˱�vԚp�s��UŐ�2S�����t�J�]��J��0ťv�c�rM��a�.��uWsb�5���y�؂� ��xt�h��P����x͵Rڠ�oeї46�M�J�_AI�a�̠����R�uFVyP��S��DZ���şhV��}_��l�1`qZ�F��O��".�_&��0����9.3���а�[X��1���a��o���x�<`w�r��z�DC�]���vp���YB����x�����g�m�ȪXm�6B���a|��a��&�Q�8�G2Q�r��L�(- _D���净�ʂ�&<S�l���*4d[�[����fW��:��l��o惊Qa��Sˎ����������J��A�4S�O�G]O+#���� f�ǃDѨw^��D��/)Q��GM�����̗ mD�͟ǆ?�H�d����\Y�+֒2���nB�M��o+��۵������3n������K�S*�t�4�q8�r�g	��迫�_���pM)IRE̪��';e��/Zb~���_���?c�LOM�ㆉqN7cb:�M7��4ӛ:����Sӱ�s�4�tǏ}����_x����~�wRT����9�dl߹�E-$��J�`��P3\6M���
��<HrQV�������!�oݣcϋh
UT�!S�N�7���]&������VpAYB�K���nU����XM3vц����b�_e�35��|4�*���O�V���+y%{�A���UHYv'�Rj��������%����ؖ�����Lx|y1p��0m�25�>ލ�%�����\ �[�+H"y��C��l$�?�p��<��@��sx��"��x1�Z�r����De�b�r�.�.�W��"��t�z첡+��Y7��T�ћ�E f�)6���ėH<_P�W����gI���80�i���0�Yq�!)z�,R�]g�řc9�z���K��~>`��VP�>]#)
9hM^W;�<�i[�I��Y���]u\�z��$�c��i�7]��h��K�7��Z�t�Ji�|��#��y��sN��YJ�Y���$B�S�����}P��Vғ�;�'����ir]���Ga- ��0�}'���H�\t���Ɓ�.��l��O�Tu��".���sL��?�}~�$�$!د$z.p�
��챍_���2K{r�R��&�Z�a��J(WW��>OYQ��5z��|^�6p���Jq��!�R�$����a$R{�W�(/P}:��wv���J���CYx�X��םcIxdf/p��]A�'�6�h���&��b����(�ln^7�*�-��xþl�n �"@�/
��>@�o��=�K�X`��� ~�km�8�JLu�wbT��Cȣ0��fY?�����Qw��?��Dx.�u/�nwj�ҫZ�I҉�!��g��QN�'����}q����׸O���S��J�˹{��K�Ī(�M���zn\��y��y�.����l,�0���%f����vM�t��z�����b��T���r7�ڛe~�*he�{��)=����,vU�4�����OO�Tl�je\�gk(̥@O�Bov��xCOV�o�Ӯ�]qx���<�3��0���i��������
r�t�xM�kc�kᤜ�g�ޛM2����"w�Kb�t+�4U���q���K�Ø���Ģ������&hةC����_��F�°�N��Ӊ�+78����V���O���Hu�(�6���%p:7s&%�z���Ǫ4^��ˣ�6��mk�$.ƃ3���L� q��3��D6L\r
{f������>��
Z��h�|׊�E˱��5k�A���	�<BZ��h�L��;�]��K_y�*.��|Q�I)�p�MVA]���>m�V!��\�'_��>eܟт�I�F��Y}�[Nع�aDFf�^�>�"�dG-����Μ_Ћ���k o��GyY?F:����͓x@���8\�RZ��W&�^��.:��M$��;z�G��;}!��9��`x��V݁� h���#�?�3��~I�h�-��!9~�h� �G��фFy$��,2�V	�>��$dI�!��]�$b�/ ���G��� c7�z���%I�77Pt%m� �=O:.�.S��f)��̒%�5_v;'b���W�)�l�K��髲�I�MK5+6��m�ف��'�I���\�C�b2�A���������>���j&a��s<�3x�֦��Nk옻��je4��i����� �m�w¥uQm����3��êJ}54��L���X�Xy�(`�s���MFNÂw�-�Ol�F�M��[�C��ϛ��͎�ˣ���`����ѐ�GnFj4˛XN?��e�y@��Y8�|���p�O�?I�y�tӄ\�Qb�s<�p���؍�,ި���9�7v�n�P�5u�m%���� (>ܘ�'����S2�&$~_~DAUiA����`�w-Ó(E�y�m�ؖ��4�:純��>iw�;��g��g�Sw�j��fG�Hz��+�ʮ�~ip`�%�U"n3x�]H˷b��k����f���>��6�Wa�_СW�C;��r	P`Т5`X��>���on�&��c���c�ĭ�'�^���0�o�����N�`�\�:�?��:x���7�����o�����[We�������:G��pЯj_�J� �!]oӋ�~d��+�b`����5�K� vV�1�.�G��J鿇()9�~��	�<��	��9�x��~�>ۍ�gS�/@���5��*hҪ��@.*��1E4M���Y��G���m';��Y�\����o�Qr'�"��u���att�O�ë~ۼ{�w�W#����D�-��s�H�)Lx��k^������mc���{gG������Q�Vb�����/�a�e8��u���(��̄�_w�7cyc��e�vL�֥�9���}���tN"�_�pJ��|.ӫ*�/i�Q��H:Q�9	���8�$و����F�L�xFhKS�6t6uN:ł�t�,"{Ya�B$o�ӹ��P6��ܟz�m����B�w���Q��K� �+�Zx�4��jQʤ
.�?�I���t�s�m]Ap\ W9�����j�Mdpy�m�����S/�<�\Xw�ﰷ�͚nl�����sjd	N���_��WV��*��ʩ�@��%���?������G;�|�Q#6�:���Z���Τ�����(�h�؍t�����δ�DA�]��Fw�oğN�+��b�CX� �ڛ��^�N�E��ZB���3~f�r��
G
�/w��5�&�r�*9Sh�>8�J*�glTD��#tE�1I����/�xF����~r��ݒnT�y"�>���}y���$��d�v�M7�_���� 	]�M7��7k=�ZD����� �|����]!t�����m̚�d���ِ;�E�Bұ�eK�B�1G�$�w��6�������mL2�2D��ra->D�cߖ��;�7 �T7B)���+�ޏ�v���!�*�3�{����&�!��*��ܬ?N�Ĳ�pyx+C2�������%1w�^��Q��6H�������2�=&��2��:l A4�u����W���C�#>n�Y�|��9o���l�Y��yi�������
	WV]�r����5$��r�w9�+���|<Z�����N1��my`���i�٩� !�27̤�7l�-�N�����}N=ï�g6�vI�&�_4e�������N.�U��]��=���͂}(|l7h��L�+��T����O��f���0�(�~��ON���h����F�b��ژ,U
��@G`Y�� 8)� ����<��A2j��C:7a��|D�+��Væ����̏\	�R���(R�q��\�q���]��
�Go��#��L����57��OOǣ��d(�Vק��/�[.��9W��.�W�&��)j�<�r�"w~X��M���A��
��x�4[�s>dj�3��Ƽ���׽҅ؼ������n̺<J�
n?���U��S'�����Vn����w/5�Lӈf2*�Ǉɰ�,�`:t����i�0o���^.
 캢Bq��ďn��..����;(��������wh|��H���~wd�f$��7���O�Kk�QB�[<�\|���.g�ꃟM���R�g,� �I��?��M��1�O0V5�>�dof���Z��v]��9���gl���tE[HNn�I��(�כ)�~ۡQ@ϫ��#	�>p�O��5�؃�����淯}��d.��j�V���� �09B�V0;���(_�L��5D=l�����N~9��Df��|�� ��t�9�6,A�N�D'r��.�����o7�S�H�x�G"���=������~\~sԣ���U>��2l����sB�π[x���ZC��GĮ�~ӫ�%zҘ��H4L��i�����X	vgN�y���	0��~Gw��^3v(Ѵ�K$�~2ewJbB��=A����|u�w[wl|	6��~�f�7% �KC>M��x�"de<˭���D�@G7*,&�3��9Kj�!](��ܞ*��_�K��}0�\���⦟	�����r� �E���m��_V۳({+�� 14��>�^N��d���S;��\�v�I����������o�<�u�r��Y��i��Tn�LمsW�CD�eS�R�e����O��*xL��W�jq:|���A�_9X��+W�#�W��bY[(��M��Lb��ܮs�(C��?�֞�JS��/Xz�)�g�����s�U{�%�͜w\��i̐$�� G��r?wԮ���~ʆ��m����8���|{ϣ���+�`�[�=,���M�]i8[�,7�)��BР�|5�Ju :�#������JS�N;~E�|b�wz�K�B���׹��������T[GI/�6�Dv��%fB$5�NJ��!�,2�ğ� 'ZV�Hd�қ�ĩ�S�A��2�eH���ro-��L�_3.(�ߊ ����UBBw��?���`�W�Y�գ!k��G�����F�v��MS�|��8䘾���o�`u����ˮXI�8�ޕ5an��E����E�'l�$�7��Z�3�'�����b���HO'��~R�����I�ք�H���Q5e���a��]�HV�O=\_߿�I~A8;�g�W��A2'�'3�L?�-�[�J��W�"��&���-�l��xث��IA�IL}��c��R�E|̟.=��H�J�CH�����Bw����Β�c�"�Ѱ�޴D��1�ݕ�K����;뱇^���Eu�UW�/6�⬝��.�J���Zbcc��/�2$a��b�+'�ώ���S5�L�6�z�tAk��v1�O"��g�f�}����v��bF�]ͷ��8^��@K�^�~�����#k=MfD�wY�	�au��8�z	~���yY��z,.�?��۔�l�ܕ��8~_w�ȉ!,�ig�z���1�JCJv,��v1���E�}SO�_�*�
�lV�L�x��4wq��&�JZ	�I]���q/�*<lTB����M�m�q �H��I��/se�|�>�����Ӑl��A�Ⱦ���s�x��:���+�mpE�����2U� \���h���p�_���F�ϔ��3��]�=��d�Z��0�
��8��ڧf��6��x$A"vk_ۿ1g�/��^6耀�󏹒�p�p��̫���lq���V-ffW�d���y���O�%���D�>_O  �9s���졞
gȹIෑ����N�x`O�K���C�;��� -�tt�Ӧ�'J����U�t�6� |t ���&_�T���R}���}%{B��&N�dWR�<���{'zi���T�F?n�St!li��@7�+W��=�La!��H�q�~r�&�tve���F����^e@A�r`�Tv}8ofccC��hu_�arӌ�T:��]���<����F�j��7�^vb��>0򫺤��u����[Uӧ��?<�8�5�(���e�aȲV(O�eD�$��l��pH��Ȍ� �ݦf)����]��ͳ�Y׍	W�4r��������-�38������֮�[G\�8�Q��ܜU�s��)J��"ck^��7-�Y�����Q\��v]zvr~�����J��]����������)��.+�v��BZ�?J����e)(�켠ϲE�f�[�A��o
�	Њ���v�/s_5�������j�w�s`ƞz�F����FLg�.tR������s���0���cGkx��>@Y�IH�MO��j�O1txg�y.H�
^ ��%��D�v�;<�_��f�E�9�7�����;b�9i��,���#vӁϣv�=r����
�H޼�%���n0�3U�&����_R���&My�C<[���"�>�^9/	2u�ۛd�.hZ�f��P����:B0+��O~!�P����[q0�N���Ϝ�+/3:�4�f�)�=��5{��S�w�^��q����_s�Y��H��hl��~��^H�ea3�&|��_58-<n� 6�b�>��j[z�v -G�/؝������p��Ty��?i�?�Vt~�#�pE}.ʚw#���׿��ͷ2��]X���c�_�!��ݝ�e�ؓ��-&Qe{%I	��}H��&ׅ��������جDc��?@�?C����f�KB��������zj�&������Y�������՜TF�,�7R߻� �8�D�H�#G�Tr>�M-yQ��p�۫��'��,��}����d�����T���t�|��*�4�1�h��s��m�/�Ea�!L�&���)b̜ eٓk%�".=��]'�>j��m���7��	Q:�����G!U�Ƶ���_8�=H���l��m5�#1����2��\������G#�{M��i��O-`��A,��M}𒼽��]9�����5#�Z겳
�������[@"�Wc��+/fP �a>���'���KY��A�}��T�EA8�h�d%Y�-�$q:U��a�]|&<j�R� '���LR���:��L�J7��b�Z����5V�V�����P���y���n���o�VN(YV�$
`nz��}j���ף�F����1����V6�,o6�媋guK��~7�VG�bc�Or�*�=Q������{v�+Oݪt؍�w6��y��Z/74��h��B���:�/m�d@��e� �C/Y��.���bS�]S~��?ܻ�$Fh�H*��F��`�SX�F�	��N���
��,{�`5/_$1�v�,7�P����}=�}ѕ�-br�M�c�9d|��1��s#��3�4�o�Q�z�5��SRd�}�&�Ë���J���OW$'����h�5�]'�ך6�Ol��L*�/ة�Ȉ\'3� i! ���ú�5o�3��h���r�Tm�}xx�`�+��5���S���⃊�{׃ۿ����>sT�7��D��$^��CO���?eY�x�e�����+�^�viO%�Q�J�1���-a�\�2�H���k@iPCq-�mt��K?�'��;������ r���_SY$�Y'5sl�R��2�-����TU-�*�Xp<`Z��oHI��u5w'F�h\��;P��һ3��f0�-��=R޵C�A��XR>	�gʖ�L�Q�����w\�W�U�L�C��dL_K��]�C���oDQ2��
�`]o?��o%Q*Q�7$j����[T����07{�r_��mc�V#�Pt���p�������+��j�3@�L�����1;t��!�j�wK���h������
f�{�g�\b�;=��VZ0�'��x��J8[�����+ˡlN:�q�n�Σ�J4]ι��)U�w�3�q������� jP���(}�~3�V;����Aـ2v�16������Oؓ�_z��;�V��j�J�9~��6��P~6��2��c6������.p���A+İ�ʭ�Ū�W�L��z6�O+x_T��bE|��2�X�#�0|� P�����)�CrKv����0*�~߫���B��� �ΘV�yyȕ�ƴG7���nD�w���H���iZำl�I6��3���@]��v�5���,�^�<���v�h�������hZ����n馊�=�݈?��"����2�~���aCfP7�O�9S(~�g[��_N�a��ݏ�������Z�]��0���GphK-�]��P1�O-O�����L��N������i8�cx��V���zAg�ϝ�s�=��f=o���Գ�خ�A��꦳"V?K���ߦ��s���g�շ�w٨�*ַ�;��a�M4a��cT*\���2�$�&��z�\& 7�f�v,S����ܟ���5�0� �sV����i�� �����n�f��i��d�4�V�V�ܞ"
�F���� �)�Dfݨ��A,�5����E�;
%I��Ш���I�~��N�"-����t�aF�f�$��P?�I���3��~��Aq�IW�m0Y_B���[R�3;�1��z[��=Z�΢U��n��>��\���m���f���^�_�z��5,W;�C&1�dΡh#��uJ�z�둥na������m2M�̭Ϟ6�z��tRIE5����D9Z�u�(NU�6
��%��|������@E����0��;�����!`b�|K��y�3���ɦ����m�Q��鯇_Ed;jS1h�oFqSHX. ����l��p��"�zu*�)Fmh�V�7��w��;Py�I~���c���z:�p<��_X����W�B<oYd���Ȁ�Y$�˩�Gͨ�r�}~Q�G�-͛��T 1�L؁���Ζ��w��;�cYu�]'Kz��!��xu���!�Qb'*vrgN^۵�Ñ��~O
,C�(�֗�S�Θ����f�Fɍ
z�8f�/Y�(V��(����md�V�I�㛋����ab�"w��^��IHKkW���T�wE�6:��_��Z��$˃�T����3���1/�3/�5Z|Q�=�߃�����,>RV9�6�� $.VA)o�F,ˮ|n�+<`�V������WSB��Qng,S=��+1~^m�2c�I؋e靤�v�O93�'��_բ!ȟ��=���^����,��Fx��t�6,h���[7�#��e��%_)3����+o*�8�2� ;1\�����U�D�*��QD)N�c�t�rx���8^�.�>�`���a�@o#�x�\]��Y��p�Yt��[C�s��~M�[̽����ƍ���>�t�Vt���b��^1����%�O:��a��r�#���	+�uv�{��! R�c75�o�,?st��a)�N~��B2-�r��Ȱ�l��w���-�ȗsY��PD
}�mp���ل[KܯD���a���w�������e�H��
	�[l�>��ڹ����g��������UCL�W�pv�)���2�Te6��)�N[���4
���vԆ
�u׵�L��7%$~��Y!-e����4�f�4�UuLEJ���?�ʟu�qZ�Տa�iA�����;H�o~5���c�Ы,ce?���d������]�y����]����aR#��J�W�b�'(��tI���2���g�@Xk��a<?N�Ea��Z��{D)m����Ga�5/]�T��Q�����ۦ��w�{�vի��pE��5�dPY��s�r���/a
� 1�3뗰R�˧t����Ժ�w��Ux�c R�t%��XB�k��wƔp�(՗lFﶜt9�vQ�T9�Y����IXO���N|nbˢ��I+U��3��ڎ;H���	]�r=�:!ߏ�zc�ܶ�&YJ��Ʌ�/��|/\t�z�ͥ+���?���1./O	/��߫�7�[ޏ�r����Nv�w���<�?bCz� 0�{oAKC3�p��3���0���G�t������5C�- �����q�yv@u�������e�[j�)�Z,�#jJ�����46	V�wGྸ�';ϫk%��1��pb�}���mji�}��TY�����#��S���M`(N�8�'Z�"�5	���<۠�b�}<&��1��̨Է;�����t����j�#��ËY��H��k|���;�~Z��z�����c~-|������/�4����Q,%����G
J��!>=[EݞDv�D�DKF/2�٧��"�CQ�������~��wo���"�V��F��|N�Ոd����HH���i��������Š��������w��mߊ��HR?Xs�l����}\*m8TƜ��,��fݝ1|=�(�TO��P�j��&3���wR��~���)	2��z��I��b㫫o�h*y����3�ΗL!_�xn?�ay%����4�������`�Nq/�H>V�-�hĎr�#׹:~�8�@�!R?��8Q�]'����O[\Ij�z�\ϛػ=J2�򬝐�M��IW��j��㸲��"�|�ȉ�r�W���z>y'�HU ��,</s��+f�ˡ7����3� ����ޑ�a�g�mW�ID�au�rbەrgp��5t�& �n���ҿ��	J!a���O%���W��པ#���slKig�eP�ү�����i,}�Q�3'�x���@h�}9�^1*B�(GC<�A�^2����ue�t���� �$L�]u7؍-�����yZY\�p�d�Z�zLĀ���H���E�q�V�X�z\k%0�����wt*���$l�Hǎm����j��#�t�E
m�5t*�rm�i�4���ʃԬ	�&���v���Y
^ЧW7N�[�	+{p{���/�^�\�[^��w���~��Q��p� ��}PO�hÂ/���x響�y5�S�hh���)�02+���c���s�\���ơWx�}��Z*�.�*��\��M
ߝ��MS�4��r���.U2kE�-0�a̪ZB�o�ܮA���:�$�vP���O��=u�|��r��4�dM�I��zN�hO�g����Gǩ�S��m�j��b=�����c�[��º=bS�{�(�����4��uW����'�G_��g��÷�ZY$�'�*W��U����·������6:�/￟�lA�w���?��u�ϕ�}Wyii2rA:~�ϝ��Lc�#��%2uh����έ�?b�c�R�g/u(�����I��¡�xF��������G��#�wi�H��7�iU���`,9j���V��r@�_�$�{�{���2o�tVDJ��Ͽ�SJJ�� �`h$T��g%WMl3��湦�(,/n������V5'�;�9���WJO`k+,� �Nx3_��6VvG�9���N�n*�B��ׅ+���5E	�]"{��k_���"�>;U���;�ܪr�����tDMM�{r�z�L得G?P�>긽
%��vCo_?9�{'���yZ���u�	_H�������ɩb����X������-�dˆSB|Y_Ԓ<����g��S�,!�x�M	�*��+�>��K�3V���c�f|���gy ��2B�m*���U\I�L��(��o��#��Z�a�6�3���>b��g�|�+�J{�*t�S�֨�.���S��Ԟ��@(E mMs��hnϿ�>U:þ��K����wUp��:ɭbG1U���Ak�D��ۣ`���:6Z����K�^���䒹7���0nkѠ����\�׈����?��������w[��#U��z�1����h�p{?�=<�rs|�0��.�ŀ=3���a����1f`���o\v6��O8h�R����E� �G|8x�}�ΗYHJv��~�.9��w!�;���?Ҟ6v�f�d�����L3�o�����#���0��B�{�w�ʲ3�U����؜��/Ͽ�"G�zLJ�΅�ʶ}�e&cg�ָa��'�l����E�>����9���Ս����B��!u�?]�|��P$����U��b�Nm�+_۵,�n=���<c�B��<RW4�k�
�v�Dsy4H��g_���ߞ�ڀ�G���򴍼���{Q���3���;�-�H������KWYi��?��h����|��Q�^J�&�em���,���^v�r)���:��:C�b
�3��,p�nJ����/r�n�gO�zqɐ2�Z��S�)�Bcv���J�J����!��t��K����昖�+�\E��2�_�wr�J^ś5��fN!�LIb�fF�;�ٲ��M~nX�>�Gr:��K�B���Kg&'��#F�;���2�7�=D*�&?G��2�מ�x���$��).��WlyZ���p�N5��M�7ay�����Z������^��kr�|LD�������J�q�����/�Iu����H�L��E�-����{��X��(Rq�Y�şM�L�w�8�n�ܨqU�R*1�.M��ȩ6%��X�s�Ѣ9��O�����8�I[�3>5ᬎQwh`\ݟ��)1�$�g
�.�S��X�T*ޟ��C��:���3���w/%1����Cy�vhB�ٯ���j����N�ke�k��˺������̹�?Ƴ�뱶7���r��m����W��Qzm;?��;H+\>�t�[��α���CZ9Ky�F����
��<�}:�f"#���?��K����b�{�ҿ���R�U]ޫ������k.�F��P��I.*��::0�Nf�����2����d��b�f���F���	˖9�{����R���?cDhR١���,�Q�w�߯x-����2=�.�P�}�/��<�'E��� {1~`�R��ei'�fq�M�k�k�#+�� {�o��e���I$$�lw�7�`�<��]&t�i㩺�) ă��ɜT�|�>��,q��v����껿�ک�V�fx��[��:bb�!~�N���I���H� �����N�����=/�Vl���*|j���YK�S��~����`R��'ȹJ���K�sC�n�mos�;���������������{�g���m���_�/��_���[ٲK������!����?җM��ʓg�S�ZVx�Z��Zls�t����	��[�Q�P�
�%Q�D�9���<��I��9�v�Ms^���P�9j��~�ߺ����k̅�+�R�g����&�5�9G>\I�n�ZuS7���-|w8���js�I޹ۯM�>3#���{���2��*������KУ�ck���[/Y����Oٝ��ҽ5_�ܷ�*�y���H<ho�a�$�b�̿֠g�����ۚ_`z���r�G�wn����vy���n��dFrr�����Ea�AK��_�������	����� 7�s:Lٝ��_�K�!3���e�i/��d���7i\�o,R�	�~R�1�Fr"�=��͠�_�Дz���:"���sI �&�*ek^�b�Kn\�$M]=�:��4��M��Z�0��o�,l "!�c�}8�HRs��[�Ȟ�+����З��B��
ڈ��ō+O��۫s�m!�~/�7��P?�j��5��[�����������E����o`�6Qyzq��B��g*�ܖ���-l	-����1���F�·���2��d˅E�o���Ԁ��T7'TA���r��d�WI�i	�--���q{
A�ܳM�)>��8�I�.�����=�x��ӝ�h@$o.�|=\��O[ړ��ߛ^ܔ_sE8���'C�K�ll7�~�$�^ר,�E[ד�*)?s@����ZX��t���9�+��[i^�J{t^�|(s�����#
�W8˘�׆b��)�Q4��z8z�؉����`�������'i�Ϫ�_n����u��:�=+� ������5q�lYx$&[��ĉ��[7;�w�6�����E����������2��'L�x�#��b��kQ���nS���N��cs/N��~��2�Vsp��=
�BC]з��O>�gx$��Y}F�G��K\}r�1+�t�VI�t�/1#�һE��D��gi�6��~�4�� U������w/+g��O��ދc�'>�b��jX�9���v��D|������D�+�^~���)[$�V#��*���p��ŦI����� �Ԟ���&;.��@��ߋ�_x�Q��[V���W���z����x3�����R�W�;�u�q�7�f��[MEs����@#o��n���0~ �e�V��f��DGm�^©�Va,s{c�-{�x7�Ӆ������6��W݅�%`�Y�9?*\���7Y}��\��;�9���S[`!�V_�0/T�Q�"ɘ�p;3b��z�q�c�H�Z��p2����ˠ<�Z�Q�D�^D`J�4��ąL�~4J۝{��g��Ň�?��[x ?�
�f�L썍$6��߱`�!�/VD��	���Ь��b�1y�*�d�D�x��w3�Ϙx��X�����G�3�N�G8��Y����� ��,:��d�8R}n�c;�6E�>��.Y�$a�r���y�I¹5�f}Mm7{r�+rN���I/D�g*��3=K��>�Zu.-��h�q�Aη����S�.����� �STܡm���I��4ƜT�7���!��n�=���~��m��� QT���IɈ����}��zX�[��~0��GN64mBb��%]���˼�������Fa�0#���A�P�VW͊���{�-繦��Ƨ�y��$B���"�ɇ�ؓ(�?���=���TϤ��,���utH-�y/���Wa�h��-����Y7w\��Yozض��am��:d�]7��iP�=n}*"Qm�s�ǳ)���Gi��U"���E��b�S[+�%����;�d�`�]+bǔ�3gz�����s<����Q���w~���g�nd�Ϟ4���H�Z��.N෣��B�s-����^zD=.;
�^�}���SS/��x����n��kie�gCvDe�Дƺc��-�LτG��H���BI�ߛo�-����y�A=�|�����fC�?,���O����hʼ;�n@T�4a�Qd��_938v;�yx�.���,�<��2 �*��g���(Fxj60[�*��9�[��ilʓ�*�p�ͼ�RMo�=�Պg����N ��(�Q��)V�R�!��c���Dm޹��a����?UW�x2�S/Wwu1��2Յ���-*$ �G�n�-܄����Ġ��j�^>{R�d��I�\ڻ��K$n�瑡p���c�OA³B��Z,E�D���.�Ԭ^@F~�R-�ǵ���.]�v��&c��(����D`��d��z�9L	O�6��s1ҵ�s*)Au�)�F�f0�$߅�Y"Xf� ����t���R�N��Rh��T�8�]>)6D��p��p5�<X��\q�L���o�5�a�0e9�5�-���V�oV��
����[�qG��[�)S]V��QD5������i7��Z-��z�	������v#�S��b����MH�G)��u�U݄����4G;Ԋ���{C���u������⎦9�y��t?1j��9D5�]�93q�(����o�1T&^&oY�����>%�067�������� �e/k�F*�jT�&�q�{ϰ>E�AGTf� Vr��N�A����Y���JG��z(B�	�IX\F����20ũFw��wz:���w�*�yҿn�7V�I�!��=����d��Ī��"��k�ݯ�N����>�ʖ̨�_l�y�,Dy-�a���%#�^�*?�i�c���-
��^]�kMF��
1P�����������?��9�TM�ňp�׭����S���'������������`֞j�����p�jV[ĝ��.��y�5`�������'�i� �H &r>���R��K��S�-�(,������ ��-��uGȆ޽g�Lu�Ͳ�Q��WP�[?�s*/��R�}������3׉�y��-3c�e۩n������z��7L�)�O�Z��6��/.����_��&w;&����E��?�{N���Հsr��_�Q���}v!��[@>L��🈩�����y�c���&�0���3_��O)}��I�_kͥ��+uX�ۢ�O���Q'�V#c3��o�
~��:Q{�Y�`7G�X�s��й���b����4���� 6VY��S���W6�,�/��.�^�~.,>8�>$��*K{��+
��1m�M�?2��=�-�B�Eq�z�pY��6�W���wBƓG=��n�����5 tq
[��Lh1����	6��L��?�"����Y/��0�q�C'�R�|2��#^d1x"qu�-�S[5�ݱ����k�,e`uq����"��7>.*X��n��zD�~�	�ъ����狱�(F�]�*9�{/-^��c���"m6�m��6]��R��z���
�����<H�W�Z9���ǵ��e���V4.?i���8��Q��y��c���t�\�rʝ)�*L3"��9�:Ed�e˝�7�B6��%��iH��bGO�UA�7^cuƶs��py�z=֥M浵T�����'���(�(|�u
k�'�Ҹw�Щ]-��UX.Dt�.�7�Y��/l�$j���j7��6�fx'>1�����������{ӓo��.���-hƺ��g�EvP-~Y���|��(<�e݉��n�?��u��?�M�Ŝ8����ܘ=����t����'8?��QXC�z���HF�邘�>�q�~��.N�8G�e׿r��y"�/{IH�}��C&�X.z�kK�֣�`��Ja�"�|'�/�H5����+g�Ώ✆9��ȭ��ޤ�#io�n�%h�����6��)ZS�-��)�ђ�O{���wIF��]�C\�G[��wӎ�sD����bh�G*����y�d�������Z�Q���U"l7����]Ե�gag�a��փh���3_��]���-Z�d�(�G:{̚o{
��и�M%�@m�v�ӟ�=�63R>D�98�[�\
of٣�F�5�+���8@��*@'D�v���G�����zEZ�-�N_f���T�ZP��*�#����5;;�&��޼6�݀�[&��`��;�bD{؞:\F����X�~;,�*���~�����q'J�$ҳ�f����F�>` ޗ�[����?��ß����$n!d�"��.)3#�쬬�M��VC*#3deӵ��h�{��{��{�܋k��}����y��:���}>¯�7�Q[�3����j���f�U��.�i��p�����5.@y�S�݅f��V6n��c.���qd�h2X/&�hZ�\�lu\��W���?���y0u��_���ͻ�^�x]�~}�J�Z�7�g!�s�ܵ)fJ��R���uP��\vI����L>Y��|��B�ι�:���	��p�K���T�;��R��\1&��O�U)c&�/�o#�#[ �l��>�����F<�ؒ�P�/7o㶎��*�O����C~\��o�a��
�|ٙYFܫ�9����Ceբ��8�1ԯ�����[�ܬ��-^�2|�1#��'!�ۅyQ���J�Y_�����{ێ�%wb;��)~%uF$�����,� O<��H?�N��v?NP���>�~([�����2��?��S��:����+}-ÑZ�����\�ˁ��c�1k��:��\��3���<v���HDa1�d�%j��b��JED �{��,P?��!%(#���qN�ؐ~�?�2zov����Nˈ�t�9�C.H�M
H4j���0Ж��7"�f��*>p�IQ�ش�rgR��y������jO�4*t��G��	*g<ا��,��)�M�#�+���m���U�r�ն^A�V�Q���-x�}~�]������j�4J��K3rrìF.��Q�rNC�&tu��E6��$mI�ξ5Ŕ�tf�$z��K��%�8-�t��uvH;�ؘ��j������˂r��ޓ���*)�K%W���:���ztH��r��K ��ߵ���h������ٖ�K��F,�d��7�Z�?u,|t/=[2a���Q�GD˃�=O.��?#�3U�E,7W;�����{ľ5Z�AI3�h]��<�$����T����rG{Ky���,�&aB]zy�U(�子�JA5����Rs�1�9�@U��:��ވ�6��x�N�X֩6^$�bXi�|!�%�=�i�����Wy܂b-�%�3��g+WT��!��z��oU�(�>�Y�\�����;�T�����\1���4n	9y��(��l�����js�CH~R	���/6���Ӳ���\[��Mi��ZW����C�~y|z��|�m�y1�z�w�\�&6b�1�&y`d^���%���/����5��6�~�W�3��@��`����h�%VY᣾d��=?�YI.:�wl{> W3�D�y�rN$eD���~��M�
�޾���z�p����f��`��� ����&�xk�kD@�_A8[�b����"J�����͹��>���*:��ʓ'jd�������$���ݕ ��;fS��y|K\���s�)y�6h/1�� ��Ï��*�N�5fd�g`�h�>I�x�[e�K]�S(*c�)���w��:Z����[�h,�o����=����׮d���p��8�Vj h4|��L�� =ZXL_Is/r��~.	�^�b�-J���B���^�b(��.j^�FC7���������@������)#r�w)oM�5*l~���ʍo2�FTw�
�f�iv�TS�J��	1��T^��
2'3M몀�o��+��h�(�l��Ƴ��j�ڷ$L�r��__�]k�n�K<0)�n|�Y~�	к�a��Rz�[&�$吒�V��2G�{�w3;�7�����3a��a�1���;z
�'�C^UH�^���EAQ-G��r�X{�}����MZ繄ɾG����[N�N�'Z���/z��?H�5��}��\��
�K�t�������ޠ��?5�T�=�q��fQT�����x��6����a�Y�Z�cǸ��a��B�TLL��n8-#��=	�N�����)���K���2�ۗ��f��)��+�=��'����h�'.dPo|��)��-�׀ �x��$�D�$��Aޅ�G3��ǿԺ!4�c��I=��d� �8�H���<;�?�"Ec�&3*�ձ�^Lf�1f�k�-�<͸�=��x�:�W/T>�_��X-}�|z�-t�?�?�(��`�{崱l�]����քu((Z�����y���:3�� �K����2f��;�HT�ݢ�k~�`Khl����έ�d�5����,K�525��Z��.K�]1Xo<=�&�t?��[�?�Rh(��ϝ��&��wJ��`��]�Y�V>Q�G��RJ���ٖd�P\�<y�O�'����M��-������\��@}�q�	�3()�����+��ئB�	��F��g�۪l�#Ǒ��Bl�09_S�UvJn??4�^��H��m��@�} �0~�N��ͻ��]�/"�<bW�Xe����Q.��ok-'���H��ѻ�9qfg�9h�9骜:�urx��h��5<o ᦹ|3����{��	_K���)c��כ7�U�7�[Ѣ?��3�&��~���\����X&i��T����9ݸ��T��p'�)�gx[�-�T���*��`g�-�������d|� ���҇�7q;U/C~���>@ģ������qG��9��V��U]���ncs�=)�Q�WZ�2�X�$��i��Z�A���>�Kw����%�1���'�|�R.P	����>�]�7�Tw�]��ݞ���n������r��T����<���S:!�4�~����rB,��� *<Pԩ�ϲ�S����G{��#����[�\5���)K��Z�y�q7�_����\�w��9�����V���Ԃ�y�a9AYy e}C�Xv�]�7�$�~�E���k�g�,񼶿�ܶ���¿XL��.N�qG��1�+5��+%�q�C�/��M��O^��_|P�ݢ]K�e,˭7���U4l]��I���5�߉Zf4���=d7
�v�bpw�0o�n4-Ő�7�
��Xl�_	��h�x�S��y��N)��^��R�5A�� ��M>W�)�:��%�+��"�����A��	X��e2x/|E������h�n,7��������_l��Ӹ�{Z��ٝ�y.M���$_�k�^6������~^Z�lOGk9�,(���^�V8��g-^��R?�K������vw�l���DTr��|�͘��k�M���߾�Rؼ޴�T ���K�M�M�>�b��W��ڷs~?��	,>�{FL��N[�ď���B���|��u5�: ���j�IWs��F�T����$|oY�?vM�7�l&�������6���kB�3A��D:��E�\bj��JD���M]B�Pϸ>�7U�5dv�q2�}/?r�,��87j>33j�hᖷ�Y��q����]��@�)0�. C����<����t;t���޽����uu�#3-�)��Lc����%�NX65���y��O��*���;�rB�)1^��k�h<E�dh2���K�IB��+5e��.O+]��Q����� ��nD|{A���?Ϫ�J"�'��G�������|R��T��|�
���$�{���$e�1
���X�SYl�~N���l��K��$�ŋ�*��[ș�W99
�<9�����9c��S�L�yL\V ���SՑ������hi`�oGҧŐWܑY|Y�[Z=�D�c�̷=��������9��u^�/�Zi3}���k��&	�ux���*�S��/�4�c�}�X�ɝ��|��f4�9~�'�\;����$�8>*IQ��H�&�z��|q�{�pC���ܴf�g��3	�o�Z&�!#���~|�O_W(u�yxk&H,�{c��ļ�k�M�/����љ_���[���^%?�t�)���|j)B�f=�l�qM鄠��sO��*A��������ѦS��MX�;G�k`$H�Pf��Y�;~��b��>�jl~�.��:���}��~�,5�mLy8"x�(��A���!��{*4�U��";��{��>�K��]y�k�a�oʀ�d�]���"�*:��#��F$^�C��+�jI��f ��u�_)d9�'��7dm<NY��f�z4�����kp˶pG�&$����˳���w-m�9WH�ϐY���yR6��(�rϊ�e��
��"^!qY�j�'iO�+=>B�/?f��-����̻���!����?5���N5v�>��0�tKV�W��fl��Z(��n��6K� ڮg��ml�yJ�paK ���KS/IC���{hz'��-[	��S|�R�f���9�z���ȅ�>:�,z	>+IjG=�Y���YH���>���߄8��������qJ�6������g�]oD����0�p�^mQ�<�zH�l�/�?l�x���P�Î��5���W�9��(#�*�D������)R�ԑ��H�V��Gy�!?ڷ��m2fu{���koh]�.ɗYI�Gu~sTc�]�n�������ܳ�	�;��k)����@/�F�;�JБ)�%��pj�k�s[�qn �d3-�i�n�G�J��7213y���Q���#Z@+jN2��bj�B:��IX&FZ(6����|�M�埭�����v�����A��}!���%l�޿�|N�_C�A��qy���#��5�WhV�qr�����"�C/����m��Ŀ8�|�Nm�ſ�������$�ș继$�C�ď�����v�3����P��#ߝ/ԇ�X��0Z*�ɕ-4߄��~��5���SK���.{jh9��c?�W�Q��>�A�*���_r�;�:�z�#��o<������S�C8�8�Q���]N+�m�?X�r^"pyH�E&�(䬎�/,���k�:VA�r���_a�2��i���N]�����6g�"���*�}�m�����*��$����Z~�����,��N �׸-۰������<~?��'"�٪�����7F�Tg�ߺ��h�d��r5�����r�-���S�+-��,��zB����l/�r	�[�#�vħ�&��]8����#�͊b��}y_��'lx��I�yG��?|��D�����>����&�����zs_8�����V�.͝�򽒴89���Y�-�f��E��MhFڻ�U��|�MO>)����s��H�Ƚ:\�M}�r��Xm3j����a�<"��%�%::�J䓠u���=��n!�f-m����ו[��Od@ׯ.��~��LmuV'��%��z� zH����DpѪ����B�(��
4�z]D�cߛOQs��<��#�Nn�q�P�����~��0)�֬����`�05��6�0]f�c��D�,��D岴�����u�u�?�5qo�H5f�w�SgV�&3e;Q�ٌ?���̔o���<���fz�g�搈���Q����>��%*��ѕqCQA�����N�m�r�ExD�=���<ex�M��r֘ͼ�^nO��2��`�o��������@��<U��&���v����0�7
k����1^��Ch���f���g]ؚΖ��9?����+��;��3�k>ʌZl���ȹ~\��HQ�߁��)������_�P��>��K9���R?��Yȝ���w�>�N�&b�"LC߻�^,�~2��=��h�ǟ��+��26Gl�n:��M�k�&H�
��>L�:�5~(vq��{iE�ûz$��	I�|~�4�{33R���[��[E���gf��>�f�^���k�ʹYM.����G?%o��<�`a��+�����oP�P���>�伢*p�-a=MH�5ٽ�z���@�IA�G�N�w��du?(8�����:	j1QŮ��g�
[�9�!%�'K�~��<���m��ȿ�����j������*�D�j&��Pߏ�"Ѣ[fK���\TU��17U%9�%�ػ�l���|m��n��F�C+p���yDw�,����s)���Mw^$�a�/#��7���O��� W{�M��7bq8�����o�����t��Y��k{��i��g!b��"(?7��k�m��1!�+�1�[tr��z
�n.��q3�o�=J�j��uǋ��0�Q�{Y��ᨪd�6qr]�;���/����{ϕw�>�	���Z�e�X}v�n�0h��	���M�	��`z	�9��]�ꕟ~^GrvEl��[{{V�o�L���J?��#>�8<{�0Ԅ�wo9N3J��йH�ћw� .���xE#hzdHH�ݪ�������jꊦ�f���=픤�A�]U�]�螰iȒ�����ެ�m�k�I�NZ�ʤ'x4<ڧ��x_�w���)W+-�$���I�˅��B|�����Q� Ғ +3��E��r8&tӶ3�����Rڡ�)?��s%�۹�,u��ׂ��ئ*#�����4<��L����gMfV����+{��R����%��R��Ǹ�Ko������g���CL$q���]Q�G-�'g�M��a��+��F��Ê�{թ�}��ܿ꠯	L�w�5����u��D���^a��5�敗[�%a�����$&����)�@w=�	��SpAȝ���P-����_I�3��w�Ei/5& ԅ�_��x5�B�\�E
�iߖ(��u��}�^������d�a�F` �q��I�~N��gf7h�%�����ȼ��=����J�~yڬd틏����S�.2����zorDN��N�d����v$껒~b��� l��9�M���I�gʋa���R��䰮-�3�^�O����{iqKӶ�3�!���{śZ�J#6�?4Q38�oE��7��O�0�#�"�6���$n��.}��(u�r�v�4�#�}]S_A�����������e~X�2�X�ǺK��=���^���G8�%�Et��ÏۘD��	�����~e��4�|�m2e�ծ�Z?d'�}�p���hz{��2�\��F�HӚ�%?V?mO���s�:�y(��~y����x:��3��gN4̖[⚽�蟱ۮ�ÿ�Y�8����9��+33:�yE�{\�� :JN��o���ãh�?�<�c`(�+�ߙ���X���]/���i?~��N��A�������[F��.��G���n4�>EG)&oS�T��{��xVh{���Jb��h;2���T�1.�@&ح$;z&�ؙn���M]�c�Wl���Y|��Rk��Y'��	ݾ����=Uw�^ׂ���*�A�J����2����Y���~���Y�O�~m��9{2�,�8���t������?	;>ޝv�=	s(�����]ے���#z�ȧuF%���]q��M�lj�hv�-��ݧKp�?�,��/��J������l �F���߽�����pЩ�a0�!ټ,."��A;��Skr$�<c�Z+��:�7���
��/NT͂Fga9�T\H\��ͯh��9о�M�Ѕ�Q��]��)|p����|ra����#�]9!��!�dQ�J$e/�����V~bGN?�6w���=�\:��Ug7!Z�����]!�7_�(�|�h���/�J?�PT!��ҏ�Н�^�	�w���=ꡪ�P���UE[��1�nތ��r�>����N�s���^�����%�R�&�]�Ba�-���Y���_M��|t�g-��I�̏�'�f� v0���l��Br��к��΃���]ov�hʐ�ùkR�v��>[���f�"Ύ�N�����L��+�	Y���s21o ��nX���o	{�~L����6h��I�1(<Ҡ� e�SCRS�ۑx��x`moʿ�+7un��&+�.��xCȬ3���f����+�k6����"5��7p�-�8�}H���1%�գDnZ�)5Q�	(��*�"��~V���S�u{���1�IeDZL&@���Al�F�ie�E1�����cݣ�n`R�/�g������;����L�!�mg��Z�8����$W*�@>��M�)���t�ʊ�DH-XeF�v�7��_�E�UTKXI��_�>�#�����
��@�f}9z��6�]�k�Q�|��	»u�;��K�m��p�I9v��m�zR𑫞qG3]}�nbv�d��qY��괯�Xh�����ࣻ���3���v�����t!w�ɝ{�5:��ˍ����ן�H?�m)r�d�_'��#�6�� ש�S��>***���1JRYIֵY:�1�	�Ν�]r��d�z#�:���N�$�Ɇ*ǡR�q<�N�͹ȍk	���Q�����/���{/7�9�N�!�{>,1���|�G�̃�����E%��]��zpXq�� �#>p3�݌�i�#���/=�ߩZ�9S����,��{�����|^�SH���3����3������T��6n�ߌ�м��� �*̓Ǩ��Ap)�����%/�g�h������i'c���_v)J��(%��L^]{AJ�ݮ�N����Y%ӿ�>�V��x7(��:���K=��4R�!�+�ͷ0F�q���$.�ܜ��c_�^b)�Q�F�Q��k�=��[���#'�;�#�H`U�/�<2N�9�ͳ��������g�����{�(����x_��Ŝv��B��浶FPr'�'���%�t�3�T������,�)�]�P�,��䅷�?5%yX��m巊�Qb��xb�]6cbX%ZɃ�&ݣ�ʚ�>���^�Hjː2w��^h�7 Q��oE9 x���3ڹ���u2�5:���A|,��!L��¦���7d˂���2D��qJ�s��7�fX����I-�؈��E9{^C��	�6+�ԪLW@=6yu�s	�:��.�Лrl�q��w��E�L]���vѾxQE������n�����r��腞Glo��Q�K���$�źe��MF����̏��hK����I���>��muZ�g	j���	���4�{[�w��޸0oJ���`0[y��)��h�^ȕe����M�{gS!�_E�Q����mO}yNL���8Б�C��92Ds���/��ʑp�4��O�I*r,��ڙ�Rc�U��傓K���%^�ȏSl��A�u������f��^��)�[�׼˔���{�ŧ}b}n�E|A�Q���G{�`��`m�E��K���R?O��ys��(��1D���{غ<���o^EX-�版�>�xkf�B� ���h1�8:�gq8e�M��ݦ��3-x×�X?7�0���^�@̗�G(�\)m1Z�M��"���D�����@��m���ƥ[>��y];�u⁩��l�
9�aD��g��8h������lc�ݶ>�ZmMR?+����7��^=J�=?%�������v�u;���V��xxw��D��N��T��gg������`@�r}{|�3z��6�t�kB����r씀!�Pձ�o�:�m)Pv�`����Ak�����_���$v\�[���ee�:�K����b���uZ�'��іQ����o;2�bi+ē��,9>��	�m���q���ס^	Pݕ��R%R�HK�y���45Kn훼jA~77�:3V�Hk�?��*hζ^c�7�G\�W�H�_��"��א#M$�;���`�?��Plȟ�o� h[R8�&��Zl��X�E�����&޲�-L��[�pؼ���_憢��F�����:M$���q~��E�������������%&+_�?�=ݸ��j������@`T�x�B ���K������+}GXv�-w%����܁L-�����G�����!��ε[1W>o�^3�--#f2@4��tp�����2�f7qy��oQ�h�m��叝b
�� dN��F�Q
�Ϋ����,[�y�ہhF�Y�tt�y4����׊���5��oodi�_����wU�����O�o��M�o�����V�#�6\E��<�=���5!��,��.'�_�ۙ�W/&M�0��ד���U�qo|��xr|(
��쾃���]��9N�l��K�n>SU�1Z<1ߐ��K�J��U #7v�|��""���捾����d:Å�QJ��[�#m��j�Oe���.k{.��dΟ/�ڄ]O&�>��!B��n�GD�s*�gz���Jw�AM='N�?H˛P\�s�u�<���
���~T*���&�#�o���������_�#��S[�:o�U�A㓨<7l�AJ���/%��?�lrz���\ߎ�os��#��.�cz�:��!�ɷ�H�Th�V?L[:pF蕍 ���4Q���д���l���؟X�D�2^U�NF�����St�7��~z?y7q�����N��u�E�6u�t;��(�������g�&����XDws�A߀W����,�K+r�S�*z���(d�w�����<8��VUc꺄�ל��C�䀖�l7/��j
�xְfA�d3c	�>�)>�y��^��/Dz����MȭR�����a�'�BG���=_J�!�S�grZ	���<�0��x#;�IPV��H&[���nO4k=�	 �m�W����N {�g�N��(p���M�\�C-����t� Q����%N_J0N�S)l#�U�f�d�2�R���ҁ��;oH�z��7����ʃD��B�ฌr)��]�+t�X]X�Aw�������>��'��������^3��0��G���		�����X�9A�rԵ��یi�}�l\��jU��Y�^^����ne�$�0��y󆜾�ǆn7�,l���=�����4lty����S����*=m�"C�,�� ^�0l�h��U��G��$�OQ��6���	ؙܼaJn�z�$�A�����2��eɤ���L\�0�˺A�v���BV���<�C/0kiÒZ�H8D�K�5�p������������|�/#Ò�}{�'�3��i�C2V݇���q�L-����qN�j\g�r����H=ч|<f��1C�$k�'Il���0nW9�n�rx�./,^V��7Қ�֯���d8������O����{W�x/�*�Ȥ���a:-Q�Ƀ{OS����<�tݣ��/�i%���,+y��������⧴d�g7�{FTɗ���ޚ*�&�L�af�;�J��QJ�:�;��賉��3zX��-��e��>h����LQ��7(�S����J~���Se�H������ �>���?~���eԲuf�-���Y��!}� 5*��D���88�+��ܵ�Gkϗ�E���tI�5K���JKun�'%�����杢C{JMZ��Ս��jr����W�6wqf�n��r�5#�gT�r��.:�/�J*�ߩ����?�j�;�����V��զ��i�}�M�4��ȭ5f��͟��ICY,��2�S�g�^l��oؗ?ٍ)��ltSc���wV6��D���_��u���Z�|��|�t?�i���i�Ǌ�#�+���\���"��ݡ諯����-F+�-L������"��;��%�7�@C/�2�Qc��c�h����{���V�D2ٮADe��Ϙ��Q���;� uC��+�$���;�sw��4Z��VYwo�Ú�b~4d?��ǘ��޶#zM�W�|2�3��{�`��ߧ�tY�\��+���+؃��a�|3����YJu_��@�GG��6�����@�撍:�Xj1�_��.������E����A�
�ao{�`�M�\��G��Ӟ_�pn����k�WY�هV��ڑz��\�Y�y�~|��Y�Uˮ��E��a�}��a��J���_|��1A�Ξ�ށ-�8¡��ݑk�>�ׄ7��@��5Q�wY�����6�,'��!����>����״�z�v�[�&��JR꾏�*���Z�8k4�TUXh�b^|�HI�ෝ�����F��ɳ#�\�=uγ���x��(�%�5O�B��(�Ѝi����3���F=
��0��,K�Y���]�����A�����I�&�j�G@�b�(��5�p������6��K���b���� �͘�x��_f�Ӻ`�}�.q�'WO֮�D uk������s�.��*�)����nS"��lj��Y�L֝��q��u�N�Cv7>v��yAk���~�leV������Du�n�YPY<,��q"���-�^���m�=���<ɇ��
����d���៱*%��&��(�&]� :؛�M�??,_c�P��kG@�ق����x �7}a�!<F��Sezp�o��0�uW��Na1f�8ŭ�l�E���"J.�2�;0� ���	�M��N}k�Y���ɦ8J�Ȧ�F,4,��F���([-.K!�ße�.�`la�G��hW��'�)�&��&«PSp7$�����gc�M<p�U^|,�&+	Sa}��i��P4�~C�4��
���u�5���=w(���yT�j�wg�-��]_�Vi`��䳏���
"~�9K�E�#�������߶�7��q�f^A���Qv.�Sj�Go.�ng�V%܆��Q`+��$�誌v�B��:'Զ���d�I�.��T�;\�q��T�{$�e�5}�r)U�����0|��#8��:Kg�/c�e���V�.IF�i��7)G�r�����Ƶ�����D�"ŭ�^K����>e��5�'��W�)����>k�5m�Z��_��p�1{21�gpx��=O�{��WN�t����փ�h��>�F;�ŷ���˺໿��ؠe��=zޠ�}h]��w�
�� ���@�o�_�00�2�0z�К��x�>I߃V�̗�1��@��u|Y���h�xi��G�4�c���c7�yū��c���n��K�n�E4/�~�|ȕ������kT�Q�{H�)S����/ �.��6�p�G[��R�
�C��4#��I��v�C�iu��_����͚]�{��UY�!�?����'#0����?u��r���ic���LͰ���n�y�2�o����v�e��n4���u�]pM�Fҷ���������p�*pf6ҥޝ�iw<�_�%|��+"�����1�'_+��t¥'�bol��K�UI�p�7�C7��Q���}{�?���:/��j,��lP[��.͌�m��:F�_�CluS����/��ZSZ���~\^�Ɣ��b;
e��*�P��
;`6'բ��?-�s#���KBf>`��u��?�����&��1�-/ߑ���&]�<k�8�7�S�z�$6���y�,}��~\�ɡȄ��%�G�� �'d��?i��}�C�^�q���H��)���9u�k�����B8\��pX������j^R����a���1�Ƿ!I4`�iY��U�������"^	u���<��w�6M{^jT7��tC��L�����k?O���1p)���"%À�D��8C��o`kv��*�t��H�
󙃶*o��Od�B{b�^H�k�M�c :>��zЦ^��hv��$0��s_��u�rX�L��+@2QXa�[}��
�u:=�n*�l�-��6�P���w����]��V֒��e�Y���M8����C.��[zR��"�_���[����� �����|d���.����H�bZ���}*���bI�Z�����Um��.1=y>}J<v�=��a6��V&_��d�s2
C3ݕ��#���y�SG"o�2l>͎w�՞_����������MU˼&����4C$)�ڢ����v�M�i]eP�������"*~��ܤ��8�����:IH�x�O�6�)���U�k��)���U}��I��'�#캪��m���+�o���ľ�LGl��-l����[ay�z�;�&��ʽ��ؠ�S�^���-4.��\�`�Xҍ����	��Jy�"�SZ�IԱ�xK�H��������K���W!Z��6:LQ�6)ST�(�طXne��֋���i* �	����T�;��ʪM����0
�π$ZG ��;7�kb��E����F��ژ�MN��K�K�p9�U)�Ŷ���bjAX?��8N>��X�]�~]��V)�`�O,1�H��ʷ��~�o:f֦wK4&��f\��Kj?�R4�E����!��U;+~�W�l����vy� ����FmϞ����;�;7�АRV V�2'�xtc�Z�Q6itGU��$�s�#��X��u��1�oe�}��
�X��������{�c;�tދ�<1<�؀U����<�ˀ3�q��Jצ��ےaY>�q�Ȅ��7�x,Z��T�=0���2�[��� rvYw;�8t�ܧv;�٣�k�����}J�z�,콋��a���("8�I�,�B�`����w>���5���n�o�֜^���@[�,�uZ������ܭ�	t�<=���7�Mj"�y��������������2�'�'�"��2���ʆ㴓���{y��Q��2b�aL؀��Y�w�	'ܖ��Җ��$���Ůͥ�����j؏�{�i#w��A�^?�{ܠ����C(�O��b������:��q>�T[,���`Һ����Rʵ�S.+M�;��KwQ�����ݱ�oG��a��y�.)�����H����m��\r7�c����D�H����N�����UnTK�5,�xE��;���2ҟ ������G���Rg�U�<+o5;�k/6q��:ݴ��#��r���b�$���JP0���.�T��e�a�▐Nr(��D�_H %Y,�aIMw��'�v�8�r�z���/0蔰7,}m\75U���2��TЂ/��9���P�5ڌ�����l�����=����jy��'h���;]ؔ�� �z$�j�����د��t�<ڢ����V�׽ܹi+�������y�%��
�`L�G��9<��@�zݠ -|~�JPms�|�^kR2#����]$������S[��t?=u������k�M�+o��^
�^}r��9��$|:��@۷���q�_A���2W��sik��0��l=(��&n| �_29>; ��O�/C�/5;m=�62Us� �y����7sDv5?`�9[op-[jn�S7������w̸-/H3R6����j�d{�p�(��6�G� R}f!F���q��������Ֆ����]ǳ��?����6�bMFMT+��Jy8��;�L���������D��jRE�q�	+c%0+�DBa)e�f�o��*��3����j}Rb;e�'�l�~���Ȁ��|W�
ya����S"�cR��I�"��ݲdW����<��� ���Uc�&�d����Z��)f
���8�dٛ��@�2=ʍ;S�����#��,��R||��.�=�����a9�å� �����yJ��~]Yx�Φ]�����k&�Z��&7H,�{���욎��70� f]��EL��/�DZvM��E�K�k�T�;lD�S}�p����!�cvJ��ݮ�H4� ���3�L�J{$\R~��5����_g�>$��`������`��Mٸ������	j"� o��۝��mf�e��L �.�C�g�ȗ<��2�F�ⴂ�y��d�ǲ'��\Bí:�V�,� �8	�Z;���q��t�z��L4�ʈ۸����\e:ܨ�W��++�Z�0!zC���|X���	��`o޹w��v�K�X}m��Y�q�V�;�ذ���f����[�G��[��N!��9x��ES@��)��T��]�� ��˙+g?˔�8�rx�9�G��2�}3k/�%�L������Gh��5�l����������I�e�$C�B�v��穒�FU��?l=������;�/?�o�:�b��@��"�� ���!�%S�-m��x�΅�k�kf��Y�]��r��*���T�Phc��7�5~��Q��w�;��������Q?�Ll���u#Rv��}u_<��w�"�}�Z�)r^&�y�xlЎ�<k��MA�^��w�S?Ψ<z3q_�{�-�ʟ��19��קK�T7������/����$��9l�~�'2M��m�A��������fW�r2�j��T���A�F�L�%$D%&w��X/ٰ�.6&"ʖ�ꢽa�l�#/F{�?<�v�H���a�m�kC�e�����'Rk�THu��|���
un�U����畓�(�
�O@�i�c�._$�d�Z�;bxzz,����"iQ�A$Z���0ȺOY�nÝn1)	oȐ�g2j%:�
�<�̈́����z��V���2b��;���7��^X��#�gJ2p�nɅ'+��tn������#��� �>�cf#M$���-J'7t��9fAO���ߴ��,4
��z�)t��`	���S#*l�&�+9;H{N���N�>b@��.;�q,��F�r�)�o��߯���.��2&��^�C%���k<�s����k�n�!�̲�>��H�e ���N�B�VAt�{���s�/d���I��d3&�ƀbC+��~]��Զ ��T*��~���*���²7��Q~7��0���*"2�<�4��L�/�z'`�x���^;>�53Gsd��65Ǽo�_R�^��p=�J�栺w����E�9\A	M'*����"��6�o�q|���1�"h
j��� 	%M��-ux|�SļS�Ǆ�o�RFJMd7����h�������*� !"!�Q*�#D�;F��"!H�tw�)��`c4��F��?���꾹o�s��s��ܧ�8NH�u�+^�U8Ї���ޞ�x>� ��u��}��@6��S��]A|ו�Ƭu��e�\Q����%�M�Խ�5w��b����/znY��&�
�����÷����d�C*&!6�� ����Y�GL��\&E���s� I�g��Aܾ���=�_�=�F�z����J"��ȗn���0\3s���ٔ����T[[�bt)���%�\��z�P���'�Z�����~�.ͱUu�8]q?Q�j�-9J�A�.C������s�	h�w����7���o�	Yّ�+�eOu���p,%q\܄8������Ǝ	Mh�o���l��0�q����i�|�&O��].KUv�A�f�r.��l�j�����wR��/n���1��0dn����)4M��\a���g��q�M��j�/��,N�oB���Ux_�@۶Ok��ټ�֋�Y�+*2:0�2�T�K�/2�O�B�dT�ֿ���
H�LP�7�rs#�-�{b��#�(�e���YVÚ��#��"�y�fw�ƾe�P�Js�@k�e�NO����~�{��g��3�l�l��p��Lѓ8�v�e$��)��!�N���K�˹a��E��
��|R���u�T�?�.�6bȄ�O��mS夂S
����dr<4��TC���������2�v��'��-������o�g�N	�fԿvl�wJ%0�]����cG��Yw���M��r=�v�ou��qo���9�����{}۬���ݛ��ʤМ���C����vڂ�KN5��Ȇ%�+���/�}�3���װj�"72ec]��r�織�~�ԉD�ȓ�~�P2*;qc�� �5���(ě�++a�!���8~5K����-�&m�AB9��T�Y���Ag���D���?�p�����T%�����jl7��v<��z�ݱt���|XC冚./S�t�Rdn�
��]Qj��	�]z���*���k�Kɤ��Ȟ���Q淦f򨽮LB�{_C�$���讽}�uGA�����絮���O�|��-��9�x��Ũ&������b[�Ƅ�cO %I�W���|��r��C��<f?�b�����T��tq^�h��N�m�} ����%K8D�E�agl��be9aK�K��#�2;sՄ��X1����-f�BŒ9��u��������-�V��4�Z07y$d7��r��57`{� !�r�Q`�L:�n?S�����#�㗇=����MɦI���Ղ�iz�_��!Ogf��[������rO\������L��um/�om���2�^,̷��U�>�~yP�Z��Kd�[�WB�Ǭ�)��q�K��|��aZ�9*�r�������_�+�1�	�{ꔡ�D�I�"��K����Y5��B�!KR<Gz���l$["	�f^�?�+�e{��q�ԒH��h���շ���C�/r�VA�=�c�*�;E�"K!�U:T�R,]��l���$�d��7G���n\��8s(�о��4`t��'�;�%[�ې����-�hhE���A	=``��U���u;�h�Ϊ�VYt�x�z�]#o�5�e�	��*�͸<R˃��'�U[~��憼��ZRB憖��6��΀�F��BD_��I����r��
��G��%�e�\Fl[믇��I�Y�7��j�uTj��v��?I�6DN�	��O�,� ��$��_�@L����';x���n�6(���r�;B�@�s��mƻ�YI�O��s{M�..��讻)"UP��s��Q�A�ee(����Q�d7��QLa˥��j�&	�:N˦��Ч]���-~���!��g\"��\��lZ���G0�ӟ)��>��e?�=	��oo�90�)t�Cַa��W� miK�R�U�5s�w.*Mi�E�Aؼ����J�P�1�	��YH3��v�F$Y�<��#;|٣Q��u�]�Pȗc���-`jx��D�f��Y��isibg\c�ڙ��T���7��m>>�XC��,Ż�z�`Ɲ?`��"?Ǻⰿ��_w�<4=%m�`t-=�?�}�׹���g��r�5D�^���7?l]���������J�-�I�8Q���N��ɷ(yO&��O$m�U&t~H���[��>�Oξ����-1I��E�g�L*�<�q���=S1�hY�ίv�*pe=�-$�����7����U�	w6s�������p�j�+<3�(�]���ڗ<(�3�|�o]���r�YA�%���I;�>=~J0=�C�u��q���_��O�I�)��TM�
+Զ�3o��x�P����hΓA�G7�BFD��
¶�@|����/����T����wc�c���֋7Ĩ��Xqq#�[��o�I܄�_k�l�&��~�+)��+e��Y���߶��k��n$�=Ǟ�y�q��)��lM���	��Ϟ��2<?D������O��NzY�H,�`�xڃ�/�]C�z즎� >��>|�GM��AǷ�\5"̋�L�a�r�GzfR]�a���"T��gk�pƙ:�m�={"{�_��6wk�^?�/,� �jL����]��%�+�n%�<�pf]ᐍkE"��O��*r|-k�Jڰd1�x	�l���]�y�H0F�'8��9�z�oh�oR���j�ƺ��B8:Էt�g+hj�5��"5<��Zd�81�;j.��!���V���d�E��\���DG-7�Y�2㻦�2�
8G�b�ٽ�߳�ctS{��Rk���R���j�z�u��gi��^�A9s� �<��t������z�ԡ>�ͷ�/}p�
mx<b��3�8 ���p���B��d\n�4J8C��B��&a��N/�39v&h>�g��=����V�cl�����5+�m��s��׷g$�Q��K~D$	�n �r�{<�	Pf^k-(ݻ�T:�*�r�����\6o�4W5��E�Hl����~`���)ʹS��t)aK�was�#ۯ���w���8�E����;�j�wA'�e�&��$|�V� C�Ki��e̒f,_;����z֦��@��)�@�����8�1(�ݾ�npʍ�S>|�?���}�o�����M�:�ؘ��ҡ��r���y���2�Z��\v�=�^Q�
������8?]��O��)�����H�Iz��ա8*6���'C[�;e_;ds<���1<��IO�t��y�0J[0Z�}��~Lc�S�{���\��9�b���E�[�^�η5K�q��]�D�b��;g�\����sbbj-{�8�ӳ�'��� �uK�}��F��*�%��c8�k�/P�1v"�I;����E`��!R��%�Ƕ�ّ� �5��b�Ik\$;��Ġ�S�����Ҷ�� ��E��;�_Z��w���?���[�����-�»���<�nr�z[ћ��2�}޿b��m��n��Z���qn���8/9
��y��z�W��RQ{��S����o��R��7��A�5n�Z�l7��rB��R��x��\h�c,���y8&U���B,�|��j�#�\a�u���9�����6�>3����_R�Ef���%u�&��1�.L�'n,�l���P���5�Kkݒ3�#_KC�u}"��=p/k5c�!�?�*Mv����Vܿ<�猕c�: J�KP�WvSKY̡��9-�ҟ��_�����7o�Z
�a��\;u=�a���|U^jH0�ኊ�f��9(|a��/c�k�<�n��3�R�,�.���w{Wv0c����P�k������ת��Q�.���`{�W6I����, �	����t�/tg�	����Ðz�vA2}h�K�Ԥ�(�@6�R��*�^:���{z���	�R����6juX�?[�P1��"����~�^I4w��!��rd�����j�a�F�Fu�a�Z��|��
���L�R�.�]Oux�_���������I��^�]+�?�����|��lb%V[@��i��5-���l���9�.��$�0���~ܣ����I�h���t�y���{_z�@H�b7��P.w�p+���zI�ܤd�;�S~v�ǵ}�[�g�.�t�ׇR2{C��v�·!��m�����l�vf�?��"z�m͙�'��/|�fE�Hx�vC3���p~�`!���5$�-�֫���Hl��y��A��%���eg��T��)�O�.��`lS?Uũ,DMT8�*�ٔ�6�����і"��
.)�?��1�����H�!���s���Ӣfz������r����X�1	i���ՆS�SCU�~��q:������T�+�Mư��d�y���(�Z��!߾�T4�����N-�v�1�t���OdRq �R/�������ˑ,�_é�@�cְ��q�o��ڪ���r�/��V��%���8S���g�������D��h�1�uP�����{�﫯[Bf��.�[�jj_5{&]ߎx�=T����*[�Pe����L�؍eH);5+��0ϲdr���B@�����*ҁ�HO���<(�`WP�o�����&��JS-:ν����*��G�1*�o����o��Y_j�n$�(T�h
�Δ�}8�Rj��
Z�mHD��5; �2�k�0�%��nD����j±�H��jw5�;c��R�2� �B7�`c@��X
�5���Q��V�$�LI-�zOi�y$Ԭ�����'����1�^}W����˴<���T�O�����܍�ۊO�� S+\n�3H�i�釞�qRv��é������{/���=]����m����,��ޭ��7�[��3���!~3Nl��`�j��
:��A�H�?�ژ��̰�9�j����xq>�W��|�p��]�<�Z���g�Gl*:��3�U�?�`�q����$y�]a����yB#$:5�3D)Qg����rLט}���5�=)�����r�� ��Z�',����a��d��d�F��y�k��3V� �:\��������w���adl�/�}��� 8�:���JbY1<"v,��~��xp0-�{�y\'�JA� "5,��F!�迺�1=i�۳Az���@#D!1��]�#�b;�����g����#+1ݯ3�q�(WCbu���+��o_.k�[���ʂ��Yg~���U9j]'�魙]H\�o�J��~	�yd�����8.^��/̳y�y`B���2�ơpu�g�_��s{�����ȹ*Ğ�N�GcImg*i6��		�)a��H9����󀡖���b��20l7�Z���&��p#:�.�Z���3k�&��T�{O���.�N�2`񚯆���%ݘ����י{y���.�!1]R2�����]*Ҏ��]�y����u�G�O|8�S�a������I���,vֶ>w梏ۓS�����s=d�:ku���ۑ���x�(��-9�%���o�/q��0ȯC���$���
��U�r/�N#��*Op���	"4���95b�<��w��&i��d�ɨ�Im��<ҽ�Q\>(�t�.����A8�%š���Ecm;"|}}lb���>��^���:���}EQJ�ԗ!�`H�a㑻�B֕ʱ�%����<}�M���<q`I�g�yl�rxߖ�#}0�s��$�I1��E�������a�T��0�ttB�|*U_�Va��������Ql4��n@�G����ՈNk\���� �� G�xr󰳂�� ���~qj����>�i�j5��k���Hq�sG�#��+����케�[�5��'�}����ǯx.۶D^�Ll*�֬��؇	�н��ʎe����F��w㹛~4�^�Was��$��)h�4<W���Or�%�n�N����*�]�41�� �GZP��/�8�"�5��8�{��["��O��ȡ@�]a�{�F��(���w1'�8���=i����������'.�pķ�"� փ��B j��+�@e�ү���(9;�����t&}g���?�~���o�{@d����x�w�Qqӕ�W��5�p��?��;y���T�"�"~���^����q�����{b�%�b��!-�3�Uxx��Bϖ�1-�<��6<T*�J����
�J:U޴&=�ҷ��|�����e'X���z)aPy�5w���i�2�Y	��X�"Hzɐ���C���u�sB�	X����s|��B�$o����od�$oK���RF�O�ei�	'�F�|"����-C[�������q�؜;��}��i�!=K�W�M�#������к�Piy�-��8�t��N	M�}$�k}����!Ԓ���C�S5nU����_+֚�{�=��7�|y]�zݼ�l��م\�,�\D��-��0)z���_лo��T���A]���z�};��l��ܝ��ő
jl6Jݢs��( nF��ط��R��o�${!m�n�v�S&���5��(��/�U� ���v�Y��YE���ks\�c�7ǻ���:�)G ���� �����ާ��8�Y�;\�T�3�B���t��̏��ȱWt��Đ�Y�4���ݎ��L��� *_���N�:b����dܗb���G\�9��� �v6u���'4�Wd�Ē��.�)��čzݎ,��Y<e���(�����PP_�is2�%�J��5g��]���~�� ��;Ĕ#F����U���f��^�����w%2�����ۿ�&��2��
����0<�����!|w����)�{�}(�|�����B�q�3h�=.���l��b���4�p����R�0��?�f�8͵V�$)X���q�_�es�)L'��>�&b��Ɵ�n��o�o-*PRi�5u+�y���>���q���JsοBe����v�u�#��R�7�d�y%o>��^o������`���L뵺�c�T)�%��aR$?Er� �G!W9�`n�"�+.y޵S��)�XW�ӌ�z>hR�������b"A�G+E�$�agxK�bIf��ΐ+d�*%rW��ON�דx�x�	��%��
oW�O��}�T��&��DfxK|���G�~O7�bE8�k�Z��g�i�����Y#��k�}����Ǆ���+sl�F7�����}�ũ�hНD�E(ut飹�<�:�5;�&Sx���=�U�(MԁGE~L��h=p\��+j �kZ����/��8_��f�%�����j�}�H�c���re=o4��&}b��,���bJ��JX�0���~�g2y�*Rc��<9�e*�T���Nñ���w�Ȩ�l�M}hE�!=��c�Z�5����Ժ���Ƙ�,�77C�����	ۀ�ˬ�w��eu�Z�r�5/m��E}��ݠ���n �����p���I(u��'����w[���
�d�ڌʞ�kl�P�3�pZ���N�<:8��!4�zy9r�����;򼆠��PM4���3�|��z��֜�\0��۝j�,�֧���N�Z�=~����
���(�E0��;�[ɳΨ%�)����[���z�8���A͎`P��Z5���R��0 Ҋ�o�G5�G2?v4,�(��i�?���BLm�|/:U�pA��X�㟐ʰ�Y������R��!b�%iS����m?��Yi �-�v)�`���[�ez���QY;֪��n�@W���P�Ox=�|(�jF�"Z��`��^ ���FwKq��/`�W�Y��*��ʵ�|TVgt�4���$+S�@�w¹�Vٱ�+t�i�H�>��yģR��N����0��3K�!�yrբ!u�r�<�~R��x�E�-^��U��3���W��*a������m
���
��p/b"ƞ��K*��Ec�P?�iΝz��U�+�ZA~qd%�'����ң��S�n�Ƥ֥�q��(�?�T���Ѻ�7�E�ѹ��6���F��F��|���V6��!	&r]��zsKa��T�v)T����v�yĐL~��\�z/�l*ۭ�. 	"�����_�Q��sޏ��&y��1w���)U�����{́G��y&���	{T�k!�rKHB��UO���}h/�Π�~�[	R�(���pX;�X���o�]��QJ��s�($@���,mR-׊�c�CKv0�<����ا���n~۠�c\>�j_�KE�s��Q������bO��7\,e�(��)�
H��]��U�7;[3��?#l���I��&R#U�P�6�}d�~��C�dξ�횥��2v���rBY㉍���/ޚ����a{T������X��Z-�F�F���D�������ZT��u�@�Q�������u�K�a8$֚ݟ?\q����T;�G�옄(k);�8�L�H�v)c˞<`��i<�%��|�sЎ����mV[_�Rс�T�A�6�4��$��wKZ���Vu�4'yK���ɦ��i�5�����on�U�{ͩ��u�[���K�
U'�J�I�@S��|,�8��	��E�����E������j6w6�T�� Og\ߵ�_��ߎ�G�|������e�-����	ѿ���N��!5�P�9<���F�F�Z�Wic���H��-A�%�t(��uI%��H���n#�t���U����.�|�8��4-�����:~3�K2��Λ�����߁V�����c*"~�r��&F�y`B��'�x�7ek�	�e�:���̘��@���˱�)�i�HK���[>����ڏ�X�V �p����z(h-�IA���H����`��V�bG�/�^L��ٷ�h����H�.���E?E�F�.����B�
p��	$���¼��0�gd�y��Y���/��W���+O�z�	��ΡR#l9VcDq1'��^(�6��D���~w�)r�m\۲3�j)��H�}�s��헝H]0����oL�:/��B�J���3�1���q{��YGv�f�p>��n���+'MD6��"� 1��r�0���Ϗ��95!�~��6	Ӑ _ô~�rļ|���I�/k_wH�L�5Nqz޷�6Н�k�p���:9�\�_�Yx�_IlΔ�[2 qӈ�A�,
~��iNÏ���*M<���nb�}�`�?�_�8
/0q���M|6s����ٓ9ʫM*:w�^Qm��)_LW�nL������iTt��L��F$_�j_��.uK-��g���}I�,��I��t���f�� ;|�W}�cƜ;�U�u�͖|�t���w��CD���G��z���L�"���	��B�XݷS������ε��F5�H�A�փ�9r8Ϗ����;���2>峃���hǦoЮ��g�"�1us�$�>�M��Z���od⮖��B�k�d��˵V��%�n�|��[�&F׸&Ȳ���h�1D4hM�By��E$\+M8nЯ��ް$#���'n))܎s*C�u ��raΦ�	�C1C��fF5�ʒ��:���=�[����G�:���u�(��qz��S��r��bs�D���V5�Q�.dvB����������R#�1dj��hr��������ɱPZ~�GN==o�,�R��^����y�T�(� �z:���~}sx\'�Y�	�l��!�yI�&!��/������3iM�&W{BOG���1]�dԗ�Y�y٬a%?����/���*�{�7�$vn���o~&�쉉A�`��o��8D����R=�������Tߺ����O���&K?����bݿ7�:W��`|������|����"ǳ��}��i�z�t���a����,j��z�h�R�M[$��_�/\�Ot���\��u1�H:��}�6�ZNؘ���g����W� �s���tb�xNd9;�=�������:���ѱ`7�5v�p���q�6H�ܨ���,ahɇ���1hə�H�"i>��O�Ha�F��IB�������1~(9����[�t9u�Z�ׂ��.AX���4M�Խ}�E�p��	B�%?^�� L�����Eu��;���쀋=ֿ8wp鈨�e�^��O�0��ϝr\��F���A��"�{��/�,�n���ˀ)��RU�7}�Ug��.Ó�����>���~���O�:�݀`��.7^k��p��@}��`�/Y�Y��2�>�������ɢ7���$���c	�Z�	��V���<M�>@E�*du-KM`k���I-[�c��*�3s���)�ܴ���y.��,S5��cf�9^f%@��DnB���O��/)(9΁B��8�[nag�ԧ��?F�$��V�K�9F�sO3R*�����X�%��<��ء�U~�`rdʒ 9��B��E��bf�}:Ż`�P\�+�����Z>h�.e�j�r�f�_�!���x>yW/b�2��S��KW��4`D�^�!*$Й�-�SI�#��`=��������k}KJq����	��O�x�P35�~�kR��)�+��|{��3V�l;<�^E� fH$r[Z$*+�w��=�+�ʀ��r��js�%KYU}
f�Yo���p;�F��&~ZmK �Ҁ����@����6�jP���0B�Oc�R0e�r��v��;5ydL���.�o������=��Z��A5�+G�Rd�V�NQ�$8P9W레I����c];�i��j����C�~��
Xo"�SP� )�
:l\��� ��D�5�Cj�V�6C�s�q�z��4N"q��z[	��v|̬�Sv�wi����
��>$U,%�jݱ!"d�$�5���#D$�2w?;dw����Y��_����|�#�a=_�x�
ɖ��IO�RZ�8~���Η6um�W ��R�y����˯N����a.�W�{��wrOV>ʬ����$H���9�}�)Gaq�"���"��C�e�m�8{�s���7�ʽ[��G���e���8�v��S|�Yl����a�z��*g�Wʜ���H�m�a�7y��ښ��ɘ�F=iy>�/s{��t�0<�r�>W��#�:��ss���A��%`q|�'�{���ml^�&ь8~52�ُ�ϣ����p�x�Ez(ϼ���ۉM�Wz�*�L��? �ٝ�=��j?_ّ�����]q��ݽ�I����/l�;io��V#�N��I�)}�a��T<�'�d��b�&Cj��|ᔜv��)��D�Z���P)d2��yZx������g������|�^����A�G��{���ƽt��W9���_P�t����iȜ;�`GB�'Ks��Yèo�vk�(餞z�s�k��/'��{������4nIv�l�BW�)~<�fN9<�XVk[��7�C�����1Z�ߟ?�7������&� E�����x2�wb3vP�@�lxʨt���T���?�4��k����⪙�^l�nLi�a�%���
'1�jhѺS�x�����p� ���xlx߀FO�����U�-�6	�W������GDйwV�y�Lz�c��`��P�U���洁�bBYdP�7�X>�v�ᱳ!>�Jn�S��;	���
5?q���0�w`wg�2� �3	��z<u�6^��x%��iYܘlIp/.%$V��Ф]�i�ُހ8��n=��V��n���ń�r�
�~m#�A*�nA��\Ʊ}<|?���@c�h�
:�ʹ(���w���K>��:�̊��X�=I� n�u����	Ah��[U����M�;�vJ�N��[~��FV��N.&���G5�[6T3�wxd��N`7%��"��z�0�9U�#�߰Cu�i�w�>nS�Tz�C���"�`���3�h�jR�{�$�D͵���>��f�lM}�Q�p���1��Pc��F��|�-r�*�Hw��3����dϏ��<��vJ=4(v�dw��OBf���x��fE�Xߺx�1wB0�9 LZ�$;��Z���C6��q��~�dy��X@OTJ���������]�D���㧻�5H�0#Ο���1}`�Խ7J�E�0h#"ud��<ƚU�l�5�]뎦&B���m�7	�l�La�&�����e1NJV�S�!=m]~�Ώ�m��?�]���~�)�Rs����i��jr87k1$����Bf3�eYp���P���������vfJb��N�C����g�:ؕX7$�u�����J�� @�?�·#�M=:#{DҸ��M��|O�r���Ҕ&2���?�Uk߈����'p�Ka5TV9ސ&5w��\o�-��)�i�����߆���;e?̖�I�Ԅ��@��_�=j+��l�O��dC�*f�k��ȟ[�{�2�r�P. �b^������d�Z�0�Nm>��Kd�'uZ�i<�B"ҢU:��7�"SV���}�=vY�����vE��ZŚ�P2Z ��	6F*\�N9�ӗ� Y���lOs�{9/ien��2����6�������q:U�0�������T<؟i)h��Vz����yT��g��D)��A�i��ךr�m(C͸';uC1���d�2z�v0v�8�䒯]J(A�)��L�@�7Ц���#=Ӆ�h)�+a§�O�T&���z�vFCJZ$Q��Һ��ح��	"�����u�'��[̿��S���r8����^��B�4�M��*���R��"S�G\�d�0WH:}��x�-�;�x�m�}����܏�\1deo������%�X�uݺ��	v�_I�B����-��.pk�81-�ߕ�rL-#5dqՒ�I����GS�x��l�x�������Fj�el���O��Fr�!{�QَV�rӾ���AVv���p	`]��@�Y5�I�Lk����c�
;Hz�ô�n�K�MB2`}�h��s�lC�@zq�08vE��5��F�d��}E�4`ϷϽ�}f�N,��w�>��7}?�*R����Ua�(�\
l�pj�Q<�����瘲��$��Mr���3ޢ���A�;��"�����|n�-e��R��]#}M�h�	x/���/�U�Ǹ<<�E	}j��TЫ��@F��'m� u	[�yF�H�k��"�/g?��4�U������'��U̱�N�:s�"���e �r��w��=�A:��PY�F�f4�C�H���?��C�N��oĳ��c<�>�ɶ�Ea��<�]~l�m�l��Bl|B����7��~���ҕ&����Yz����H��j�����hd����(~$�a�(H��}�8���H^�����wD�?��5��>����ҭ�v���ܐG����9�;>�i5%�9�gځı�QJ4��)J
Ri	�ir���S��3y��q|�$ث�ذ������w�9J���[��T�a��y�W$Z[;#�Ux[,@�PC��?�W�!�g,��9쉙S���%S8Y�M
&�pv��,����A6W�A1�V{}�1�C���s�YhQ�(c�#�R9
�pD?'���w1A�G��ai
��3�v����s�zj� �O�Ų���Q��j�Đ���H,��T�s����꘾�SV��n���:��SK�[-�_�R����2���σ�rs+����������d=Vq0a_@;���̙��#Y�i�ɯ�>5�hT��[ދJ�E��9�>P\��S��aꭱf��^�wG�@D	�� pl��AζY�����--�Q���iS��8�@�s"��G^�3�Q���H�ani��
���3�4��N6M�ћ,6�5j���v�緂��{7�W��4�~�2ع��8z���I� [��I)�4�!H�L�.Cax8��arW�՞�ǵ���R�L�l������^k�xտ(X�~�����9*�{��'�L8�urS�J5���#�$,#j�C��M�Ss{9ƨ1�6��D�0 s��YHߧeͧ�^�bih��.����]��B\d�K�,����|ͻsS�t�le�����<x����V���Ɔ0t�X,:=����=K�Tm{��2��Ɇ!�%�p��/�����Y���5n9��f6b�����:�^�$�w���ߚo
���L�T���
�0���x5C��j��3ë��ʍ�K�6!�����,�Ⅽ�j	�]��!��3����DЄ�a�Pxo�`2�{T~�ش�����qD�d}���g`09(FaD�b�씜ˈt{G.���xǪ�� B�(	����a�8�ک_��6|M8�� !�sg#���=�n�7��Y�q���dϴ3Z%�nص���;��orBh�;��f'G{��R�}]9�6��,�=("�{M( �F�:�5��%nB��ߕ2���;Z����T�:i�n��7t�Re�Я+"�{��L��I�%V������Sg�h���X"Q����FD?�ʤ����3�(��"�?�-��mCja]1)���\�z��s��9��P����C��y��Yw��"��wg�e�^�o<2�����}xd�:�9��)�-(/E���m������D��,3ؤ6��S�)�C���4tx�&[��7�cr���M��M(��ӷ����G�ZR�U)�m�{vp>��4g���'����{�?�/A�I�`�-@}j�J};h��	�E�TT����vJ��zjpҀ �az��&[����Yo�0??Yx"O����x�}Λ�j?A��t��b����Y���@b�nYl�q�]�b!�h@�$���r���w����m.��"[��@&����h�g�/�S���È�@�����a� L������I��ӗ%�=�/v!�-���jpr�v>&T�7��x��j�I�Vx��I����.b��d��aXH�oc&�uu˥���1 .�NrSS�`�Q�xEjM)����A1��:q���HUL<�o+\���+���O����+���Z Wp�I�8���l��j�/�Ȏ�V�0ƛ8�~��SA��>�gH]>�Ǿ��P��u��t�Y��Dd�MW�C�t�4����0�`W���|V�9��8�=�<T#n��K�Al��47.���Y"��C}� �^z��Q����K?ɞ�2":�\b����7t��T����c��E�қ�r�����r�&��j�@���ˣw��t����z��p}���S��Rš��yeP̃����M5ip!9=ļ��V�IѢ������"�&C�nL�V����e���Jy��sl<[S�:��Y�P<K�۵2������w�PRǴ�Q���66ԓ�=D���o#L#�Ƒl��̇��4W�^��d�x�&E�H��z��G-#�6ze��<+��������K+���
�|�c����~X#]Ђ�AiE����A�����B�~� ��%�}�� ^>��`f����/�Лp��.{�F g�E:o�����n�u�e�jo(h"ev�!s���ˎ�� sBm:s?���:��|�d�E��Ϲ������D�1��K/��s��!z~_��E��+�ڔ�$�"��%��"t3H�<z��fZѯ3~�7�����!�:����3�u�M�R6ày�hΜ��:��x��q�˕u|��fD��P�� 2A�/�҄�Ġj���k_����� z�ةNg�Jvk!{}Z=���7j��1�q骖MTŒN^��z�'ǆ�gV�h�0(�?a��MK�L�KB4 C7�7�� ��������?�U(���<8�?���9�޻���s`Ö�=��{��A����	�[t����{����������I�S���ڤ��hgY����^~��䱁�w��{��?���G�peȦ"�vt|7,�
����oGbFB�S�Y��?�$4��g�*[◴UȆ�3�T��`|�D���?r����~���+A�[���6��%T��C�>�"+P���P�:�����Lѵv>?�h�;��3D���7�/�nd�W�
���Rm���٥ [mͰ��L�=YNV62u�x�%�%�!*��T��{Q;0�W(��wu"]2s=��:�g8����O��D`���A&�r
���+ϛ?���w�U@P�{�0Ղ��<MZ��=
YmV�
_|S�7�}�2�@�y�Z�$0�,�j����?BD!f����p���'��[;�ω�EMl~+F�����뎿G
=E��ZL��E�|g2!�KL8�u�u��!����Ks��q�5�]:�:|o��Q��w^�"�W蝳�:	'Ӏ%c!@#l��>Pn�2W��|�;ԒY�M���=I;
b�Fq�κW��{�l|�2�B�B44�~�}diFb�R.��ۨ\����r��d�W�����yFM:.c��$��v�ٚk�P��P�݀k
����c�A���
[^�.i߂=�nB�j ���K�r��H1��V�J�'jF���M�O:��b���j��'wL��ɞ��8��n�O�	�Yݽ.N�&K�ʼ�c�o����櫪v^�lBD���ؤ�2(P��7�ۤ���)��)O( ��,*�W
���_�n"��8D���+g�R��yK�ycg��#�Ѥm���<(���t���7Q�W���ߤy�r!"�SJ�,�Yƌ����(�'��%ڼ�KjRW��{�)�Sܽ�``��g}5"oH��9"o=o�-t�4�Ey�B+E��7�%^8=���d?@AҐ=/�<��G�rH�X��sY��+�r��2Nj��|��y���B�<'���#@I���̧s��ސ���1���P���6�'�,C%!�la�w�d�^�LQ�u�{){($[d�w�A�){v3�΄c���5����������{��<��>���b����ݗr��,�6�o�V�_��x�W� �Wo�B��|� �,���,���E��>{��)�������U�د<���A����g��o@jV��������L��勹��4�����+�bO�5)A7|��{����Z�l���SB)~~fȞ"��uq_"N�Ӿ��Y�z��۩[g]�)e�����\��;�����n��'[G�E����L��q�j�*���+�0�N��i���R�[|�15�bs.#�:sH3D+du���=�[ý�,`�#�kNs�s���!mkk�|�|�����Y�����ݡW�u�yk� yQ�� �K�����g�j���T�龏Ӓ��	���A^�Q<_9�������j0�~�S�=���PpzF���[�(�َ���g�ޱ����9K��	�ui��q��:��1]��*�n�P����5y�D�꫙�:���ө�	%��_h�.QQ�BY~�@4�f'��sG�L*����g?|=��;BgR}����R���9��7��PR�QhRK�9_O��l�ݝ�ʵ����S��M]d�*��K��]5!ho?�P�?]�x�f�B���=�K:�Q�.�]*�ۇiŗD;E��
us���&[��.rt!x�Tw��X~��� ���3�\-����g�ZWf]��*�x��.Y�L��׻���X}K(��d;�x�4��J�J7jϗ)Xߪ�[t ������з��'%��[�_��0�_����a���Օ)A��7����k�Vۋ������?�S�:I�'p�Ǡiς(Z���4W�v��l�Չ�%�5���n�:��kX��W��޵x9;Z�� �N9=�����Y5ߛ_�
�H=�@�8�ṵ��E]�V;�C��+�=(3`2��QU2\�U��ZR�P��1q�J;�c츅D����θc��iXP�W�s���5�nݽof�'yo�q�e��9Z��k�]'����5%6�#�_3����N��>TyL=L/���tp?r�_�U��1t�$��#���O܊QN3���漙\��qO{a�w��|������dv�}hRI���G@���`LJ�=�+��G��t��FP��^c�f�����w�W�/&/�(��o;�4�\��:�Y�4@~C!�.�¶X\Z�x>��*�ez�&]��mkk��N���D��ݹ$�4a�zL��S�}���0"���X�x휗�]p�����j�n�ؽ����+F�ka���ΙΥ�j�k޶�����)le��;O�3�39?5��b^�T�ܝ����:S1�.حH<�y\X�f��N��| �>[��N��5X�\0�Z��c�˟��M,��[I�ʕ| ���?�X�ң9i۵UEԓ��R�_l����FdR���7���q�N�Gk�u(���[��t��̙��
ʪOF%Ǿ@햄��1��zQ�ϠP}�����S>�%�������}�������JJ������������h��W�G�4?�ԋ�bKfY_$6���D΋[�����Ӎ��%P��x7R�3�ߙI�q2��~Rj~Ys@;OM��a>�p`#*�W�ʨ�"�"dxy�oS�3�o���������HbQ�Q���7׺��㶇�^N�j�Nѳ�ŊY-"�
��Ѵ��uLԒ�2r�A�|ڂo64�U��*UϾ�/���C`+�g�)��V�,C(��S������ԇ{�O�HyG[a�z7�K*h8���X\X)]�4]%9i�KK@rY$�n�S"��$�y�������ɇ�r��c|w��w\<J�b����9��D�y\�!�p�>D�/�ߏ[F�zg�Bi��-T�[�Ϗ����0v95ȏז����߉��22��!��Ɵ[w ���$���ei���;�D�+k�Uhk�{���aD���]5Ǌ�T�)Ej�0�|��7}����a�B��G	\ǽo��?{тf=��e��k�B4���/%:�����]/�:����^/{n��n��;d�}�ޘ�zx���m�����s�S�j���D|�!�7:��o�K�\Xe�j��Qi<"�OMEk���O�)r�7h:LQ3�A6.�C�����w=�p�G��&�:�15�n��2����A^��ִ��U�3�vڭ�Bbd#i}u�(�p+ަK�+L���^����؎�ʣPL�H��}��&�p>�s�-��0�#K��&��A�}�r	�\wp����EGBfuuk^5��aOp��F�v��
�j������� �i,YWϝ��&+�	X�L�3;Xf�� P��V� ~W:g�q��"\?9�.�b�Bdi�g�mZM�&���q��,4�J7�C/�v�ߑ�U</m|�`W:@p��Z�=~��A4�q�>��489��������9y ���m����o�EL`s�]�J8���E���v�<��iY~�$�2G�ה�4gŊ�O�"�uӇwÛ���FtKo�t�@ ]�:{V/sI��j!`f�x��	}Yr�tI����GL�J�5�1��b�A�3��2�q�LA�fj�V�����$�y�Va�)b)g�9��s�/��Y�vV�#O����G����p��-/ ���g��=�����!��+p;���_n&B�L��� Px ����^Qd��D3%:o����ʿB)p�]���>����W������Y�=7�����8q�R�(}���/^S�9XT���w���^G��eS[MJ�YhN�Y��/�&�j�GY���L�l�_r.���q��aE*NQ|DݛZT�����kq�bS x��L�x��G4d3�hBX��5�W#�mG{hd�^����݃��U��q��g�ҏ�Z(X/~jN��KwXsZ����1�^������.GE��t(����/b$����t�S^{�!�ğ	q��ή�o����8��)�=Ŵ�K#nJ@�+��#ݫ�Ҷ�p�#�F��Q|f��Ӣ��߸ܴ�r�Q����JSx��k�;6�@+�h����bs2^�^���@�N|����'L���USG���)��%�߆[�E�s�3�UW��+;�x���>lk<�EǛ�_Z�~�ܢ%dSK$4o??��[�lN��&�sW�ab�2[װ@Ap�*��3�<���d`/;׬l��[�{<��~��l��t}W��6Ԏ�8&�->�H�x.��k����~�m��26U�hN��}��`{�x0�O����E�,�xᶃW�%&OA
5���3h��0��=��B��"�o�ϓ{I���Wɘ^��/����7�W��cf ���a� NP�/V
�+��WT��co%������6�����6� �ͤ3����=����ྖB�Uy�
U�3*���VR:~L�;0~�,�� ����Ks2t8p���:f�7yD��N���R��\���P���0��Ei��CJ�n�F�z:�X'&���/nE�P�䏌���[*u�/W�*d�a	.�(1u>��RVMqL6������<?<����A�7���K&����%s�V�cI�;�h���~r楪�1V���R�q�?�EG�o��+��C��X.�\R���.R�1�"�إ���Z�����<��釚_)/l��L)���|���V���˭�h!֜�,��ܫrx��n�"��dw���J�����<������8��Gw�"��c�)ѐ{w��1W��|X��,�U�Ӆ8�lA�� ��<D0v?�o�m��1T?^�� �%�Q�ư�B�H��PIC=�Q}9�n�X�\'g�d:>���:{X��:��7��I.8�c����k��Z���ά�h�D�8��E�j�;i/h� u}w�[$�o���;n�H�V�̕��w�X��J����CܛE��9 ظ�j#0���C���B��b�����ze��Ũ�LXn�:LC�Ǳ��4˘��鹯�羨��(��}�X���,�D"b ������5��)����r�s8��{��OOѿP���<�Ji*�_�?��kq#oů�C�o��O5r�j��Db�XI�7�$H^9�@��C�5?��	Jl��R�\I��J�[���}w�'WN�@�11`+/�w�:�lGm7t ��ەm��/7�+#=[��z�P��t~���h�N�{�1<r�p[6� ��R�[���	yM
�r�E��r��#���|�Dc�vo h';Ҙ���8%osȪx��|ɋ��4�o�Qq~��
��bpp�L�'�$F]�6���c�V �g�P8D_���?�����܌�G�11�y�$W;ܵLC��f����a.��z-�z�u�
���2H�h`N�C 6og���̈́�>�A~-n�T,y�t��ua����4��zu�2'< �G��}��-�Zj�4��ӾN��_�~
�\*����a���_hך�@��{�.T����'jOj-�ݏ�L�Q�qôn���[������4�Mj=x���MoE%5fA�CS�W3���Ve�Z#��E��P*��[�Yo��+�������;e@G��"{�ݗ��\��u�횩����MTj^��+��w����yU3�W���U���W���8לF�í�2�u��!n�o��
fM�"�N�z���ު�F����%��=���4��ۖ���l���O�b���}��I6����̕��]|�WJ��}��46+_FS�����:YLq���)W�����G>���e@�������jh��7�f�%ڻ��s3��^qƃ�0[U�e����ǪL��^��-���n>hH���~��=]���n�C�R1 �'�@��r�_&�vwO<�-ޑ�|��')���75|̱��v���p�'�z���$�b��'�X�x�	���"���sL�?9 :�m~��\K,��V�l�8�
�;��[�N���7�H�ўk���w�����2+#KU��k���Ƒ�*{�<�!׍����P��b����3���d�q���N��d�k1:{a�|�@��6�V1:�$���d�Bc���;�$��C�'v�
��>\b�r�mf�&�㦜<�Os��f�������֭W����t��>_�1���8�j�`��C�Y}O�.��߬�P��/ �^鎼w�����,ؤ���k!a���D� t�� �f�:?X�E9u�Q	���i-�9�"��|^�����V��i�d5��!zY�b[鶽�G���C�CB�0�}͙�g!: a�����H��@"�����lF\(�NM|�,��k�WŻo�g��b�}�Tq��](�lų��'�m�����榑��X�~gK)��Z_���q]��U����7�J���J�+�ଣ��6{(�ڍ�1�<�6}�������@�v̢d47�B�*a5��w�}*џ
���w|v�g�#�J̲��b�A�m}�(��w~R}��B�v��U3��	
��"s�og� ;}��pX�����I�i%	�͏�y�T�J8�#�FF���uhۖ"
��o������8���W��-6^>�/[���k;�Z��F��R����=�j�bï�գ����8����5"�������L�߮MǇ�%&�Ϫ�ȿحa��R�d�����Z  �	�]0���id)xu�����H�k��
�Y�)�-t�6j[=~MS� "�X~�fY���I�`J��#���i)q�+���J���5j3(���SW�o����P�{@3Zgb}�����i��/����E�ŋ��J����Y,�P��f�Ќg�!�$�q���m��\A�8���t�9�a�7A�	�Zf��-0�o��k&|+ii��vpr�O�� �J]� ҹW���mwN렦�u��n��´c���s� kzh	T��(2���;�&I~Y�]�G�_�א:����B]�� k���"H�r���X�x�d|�<� ��a�|�grUn�Oo��/a�@;l�0V�A��k�7_������Ҡsȩ6��D�]�l]5G�j��e��ۏ�&��!�\�9�%�b���������ǥ�F���=Ei���f��H8�gx�z�s�3s}��/�w����d{X�q7�L(�V���}�u�bL�T��R?�Y��U��'G�IJyZ��Y�?6�up�Q����7ҽǡO���h�M�0�%�KVXN����}��{	:B�s��R��T�nvxf����/�L|��؄����׉eT�%�����N������/�Kn����Q��o��:7F��-�MO�.H4�s�]�r�|�Y��>�[�x�2Xĝ�u��
}�g��,�a�� X��+:!����dMB3�����Gn%s�j��t���0�� ����m	{�tM�6߀�UmQ�-}-s^���\m)_��7� �x��-�Z�j� ���F���]�yf���(�8oA�i�9��f.�������3ac{�܈�t����8k�ݯ�u��4��=�~����}�39 ��{��7\��E��	t�9�W��._@��hjM�A�4�D8�m��Ղ7���w�	�߉xu�����Hk�Wդ��]��Z\���%v~e��{>_���~6�`��T�Ԗ<���£��j,]T؞(�`��Ql�8I�z���ʘ��a7�/�wE����B$�'q��^0�G���P�cq-k�|_�ҽ�����몿5~���YC��*S&�%�h�U���7ԊT�V<����t�����x��-�|�Q-�e|�`^���4�]�D=�۹q�٬��;�4�Ӧm�d�EC����<k���� ���VX�Q��w��a�k���	�z��@ܩm��נb��68��Q̲ʃ�#��㭣q��[~��_��%�����G�~ �Ӓ�ZFof#$Ҿ�b��?���1��^���;���=����+���1���Ѱ���9��>8\����`�,�E\���sfu��P��%��z:����,�I�Y-���
�.bS�U�(П��o�Wc�WS<�[i��-���fcX0��ee�&\*�(��r���@�NS���%hCr~L+VJ|�}�v�{&X7Vۆ4yA��Y�L���E1)�]\w� ���M16-i�Y\@m��9�	NsH��7�|�q�����`���1�/�v4�[Â�o�h����AO�4'I�_�$'����}�6�Åu��!�i���>�E@g'l�W�i��S��@Kդt��K���R��W�������ԝ�G6 �٘s���Ř��@�^p��22�.�O6�M��|H���}��<��#@s��˞�ʑ+uY.ʋ��U�k.7���f��}Y��vS��V�s�&�{#w{�S��m�*�c8Ӈb��I�_�nV�|'5WRϽ���X��K#� ��"�_���ZA�^o��w�K	��z�[���G�O|��Ui�P�Pf��K�����˖F����^�v}��~�2�}��k@�Һ��o�ơ�$�1��A�$Gm�g�P��n�U�F�q]]��4����d�'�*��n���Dp>�f�Ow�Z�(�Ǒ��O�Jϥ�'V�::-Iq�����^�.|�~+ڌ%�U��j+QuzF�����Ֆ(X��m���h��+�8K�+�Ͻ������,N�U9w��-"JiY�h<)b�>�0�.,$�VI�&�e�%���Zۻ����".�6�;	�$�f����ӭe���y7n�������U��,L�em��9e���w��V��+���/�<^Ѧ��i�L����g��y�X%(~�S�%r�^᷈��Q[Gq��1C5>�E�{�;Y.X��xÅs9gU��뚊6��?z���'���R��;J8} �]D�Ė@p_h!B�J�^e`�ؗ8C�<-�Bi>�+����T��N2�z>�/�pbJ�������*�\5�S_��,u���Q;=�V�ӽ6i��:MqA�}�Ʌ=\B�5X[�[1`��Q�/匥�Z���P��2�R��S��aUaj���W/�Ǵu�rЬgT�񡳌ίa�?m�f��MoHOҚ�Ws�Y}'��-@���/;*A����Cz��u~���=��uXUxmTk(����y�t~W�6,�/����J�~��M��w���s�}}3;�?��"w�҄w�-t���Ϫ8�%��{8�uN��TD�`�ëW߆�����������\ɚƾl�,��|ʜ� �XK!vZv��-�1&_y�����b���02:U%���"K�t��������h�P���2H��+���nDۄ�۱�ܙ�t,nJ,]�Z�� ���R����5�c+�S�M��`�*��b�3"��=�����{��;��`g�>��1�r��%�u�/���$tO�#/�Z��%��ML�)J�S��B��-ĳjk�0?��uP�w�ۋ�)p�UЁwǳ`�sD������^��^��Aw$ϴ-N��'\��C�O9Ƚ�7�����U����>�uk��&��I-�k6A�B�m4-R���.�+�<�oM7��fMeH��X�X�ũ	O-� 1���XE�Yt�
��ﴒKO)VJY,|�<�П:3��r�0�:�k�*��G-�|7�Z$�"%�wF�r�E�W�"-N�T�~�;/(�?d�\���\�P+�k���� ��=��6��{��3���
�l�C���?�M����.P8��ٓ����9���?	�/�c���Ջo\
�	Z���."����(�ڋ�\�v+�V�lo�N��Y;�/�y
�F4Q�6�o�� i+Y�������ѧ5v�χ��i������������XvL�Eg����h��So��5�_�tR�!$�Y.���b2;�$-<���u�×�\_|-��s�E헊�/��?���+Ր��1��G�q�_�1Y�V.ۋ5�qw����m�q2������f����p�N�=LL�h�v�C'�?�pRqC�ِ��!5@:����.dHʏ��?P��̄Y�b_P^Mf�ѹ;�Kpϒ��^��3α2"��6�ךv�u&��,џ���/;�g��;zk�:F-�L*#�^�һ���5��6�����N��Qc�۷�2̻m|���J�짒��%V>nBe�p��s;�'�~h)^�8�"�+���`�U'�+(�`�X��Y�,���h�M��_��Qu��g�t��b�����i�K��0̕a%=���a���<��apZ�3�Q�p���֨��A}�qk�}�@\NSD��B�+	����׾�@S�k�ȣai�bӓYT����U"/;����\���پ��ˌǆV��"�tf�N�$���D��ƿ��2�R��rx��t�a.)��/@Ϧ�R���,4+ϑ[<�-�X�Y�\e{���gY��+�b�Ҡ��/���vV%*����&������E��}~i�Z�~�Uي)b���Q�sTJ�~�ZZN�W�~	�wp/SG�wx|�*�؞�ūVa���Y�l
���J�WI�Cn��-����.���dש�ݹ#��v�4x���>���Z�������>�/(���ǩ�%����t�X�╣}[�}:)@iܶ�՛��qw���u�c�
�w��k�4D� �F�j�^�@�Sp��|n�b�Η�i�	'�n�.>њFE�Q��� �~�l�1��G��q�wI,�5�Jҁ:�	R��A&^C�]7N>�f���n���*��l��8�+4���K ��=���R��\ ���4l]�7j�FUN>�I8��w�@4XinLj�v9��K
��u�E
���/��)���ؐ6����?�?`*>(R��e~)d��4J����1�֞Z��y�{��q{d���s�
D@�cBVvq���+`g(>)�OƋ�a���/d����FT��R����ORUٺ[��aߊi���˫��%�d��nEΩmNG�n�>9���k��[)Cq�B�ñ����A��n��[�d9�Aĥ�}~5��V��+<蚽4�φ��̠ȇ�"tutC�=�Q�=�5A^��f����)��F�m�v�R#C�����~�Z�'�����C�~��>��8o�b�b���x�p�n2�W�F���"J��X��z�7ǐf
i��[R�h5k� Q�b��^�Z8���vjH���~�כ\I��.Q��wC��=����^�	uٝTv�'9~U�Uнd~�!,x�x���%FG�p��������'n�aħPh�=�@퀟H����u}tb{��;)��b������Ƨ�?`�#:��eI*v�U��8b���$ݰ�Ϸݟ^�^���4q�ƭ�#��7��"NC����x�-�KU׈��7��O9�	Ol�+���;�[�O��������"	��ۥ)_��L"yy9{-�wj&����"d �Qr��gM���gSx��U���fZ��f}�8�e��Ϭɏ������,H��ѿ�Qy)�!FDZwDiP�w��}$�����KS����)V�CF5������4�����@VmnM0"Ѹ��f(Z���8����0㺑�)�����	r�?j	%+_>�P�	�T��4𴰹�Y8��y�Z�(�����W1?���v���vr�=+�FU��Քͥi0=r�mr厬���X�-�rq�t6p���d٘��g���/w���h��_qB�}*��/2V��;^T�A+���C�
?z��(In����HϬ�!�F��5���? d�|=�/=0)��Qm �L.^�-a��6�Z?wy�e�Ο�_�$]e�mX��a"C��[���������{� �sS	��īA4Ȳ�+�4#/��M�b�������ɣR�Ok���ʳ���STP��_E��Б���8WZg����)!dg�|��(Wȝ����S�l��T��F)�㬾¸#=Âtv��żfD[G����<��j5�^H�OIm�w�*����](�dsB�`A�{�q�W,E*�'���9M��J��ƾW����1�?SgtM(=>���� k
/$��W�����b�c[w��{�퓈�}�c~sLx�)��?�ʯ�la��9��Bsyg޷�sB��5�J���O�;z�c���F�H1����+�ͫ�&$+����5V��>co9�n[:�ݻ�ư��?!�w���y���?��?S��8��ɶ�b.��ZR��UUF�
���ʪ{�2xŅ��I[:ht�=��c�|�g>R
y|%]���.�U��Z�O�-�7?%���tt��sJZ^d��0�pn���_�����泋y�%'�2)N�q�����/Zx?��j�pc�+�������5ӳ�ӫ��
����Ƀ斅Jb�U��Z��ǡٰ;g�N[�֣N{���\)X�ޭ�&��e����4D��T����'�ai��M�8���$ ��p�F���SW�ܼUa����s_�?i�RPqD
!����N�FTzIh��jZ��J5������VD�/ُS�T���jlYz�H<��]>����§�ǁ~���=�R�tׂ��R�������5 )�C�[��ƹI��0���''1���̪85Qk �s�P	 v��� `�9TI'<��t�.g�g0_�Lٽ>'��ktW1�7%Z�*pg7���$�R.���i�פ��D��&C2V|����{dXd�:�YK� �r�G�L��b�$�S⻃(���Y�UDSm\��Y�t��Ts˛�n��@���,_���2L��\��v_�\(��Z$5��J�%�;���d�{@3���2�{~"8���n���x�ůlN1Ν�Nan7�ԿZ�Dۿ���ia7�z�Z�sk>t$G� ��;Ň�JM��2u��0�y�[�����rg)�I�G0q߲�q���"�pCW'�^hLl����-U3���в�u���`!�q��#�Р�1�q%u�\a/̬+�`���}g�W��~��vM�
Ӝo~�bH'������}��'}�tZ�ZJ���G�����������߹ �\��ǌ��J�zy��pj��dU�;t6�e�XR��aP��(C��^v}�#z�J�B4�]$U��ER��U��\  /�x!8oI��$�8o�e�ߍ.He|Kǌۓm�8!�܊��9���kl�@+o���ZsU�U�9����:�<7�Y+����s��v���w�����0�\����SN��8�S#�ߦ��~�n�v�F�w����0y�f��%F�����ž�d?N
RA���NF2�q��(6S�l:Kf���;P3���B�E������Jj�8$��A�m��:�-F�U�yw̸/�.��$W�C(�-I�L�\�:I �*X7Ø:���GJ�������;<�9�2�`c=wD݂����#�(	N�\�;�즺�?ϸ�'�ߋ���l\%�(F�[��m۟���I�<E����M�YXP�RK[���)���h�[T%���E��S�D�4����G��MҾ����yn��Җ�)-������a�8�<��w��0MzA��i��N�R]D�1�����?(�^J��p��\�"�7J%�N������	Ks�c��
�j ��[p^�_:����m����c-�D���N�oXx�Dm�i�0{���S�;ǂ����~^�'�B�Y����k�PO�;I?���ƪ���rŮ�C����q*0}�(��K�&B�)ah�dݼnBu����BY��(�bH�f���E.am�nƘ�ֽ�e֪���Y+Ivh�^ ���7���T�9�cD���o�F��tp˳l�����L'��z���4�'��#0�����̵�d�-;_֥j`�l]���J#�i�t�n;C�E��[�~T���X��$n�J]i�z'�|��$a��<ױB�t{p78�����������hT�G0�GUO�n::?t�Z�e��9Z���skP���]��X���Q� U��F_v�g�̕}0���pMFw�|�7��dc�k��b�pO5����놣�Zw�8_�$��a7=�lf��_��ӌ��hʛ괶����&�ٍ�)kB��)��3��P�M*C�f ]7����no l �� Qp���kt����/�+xЛa�a��5+�}6�7G���j������vG��݂��ujF�wRs���E�}�$�&HѶ���:�����+�o�F�I��.��C���Ͳ�m�R��M/��!�_�%P���8/;��� L���t ��F����0��/L�s��.[��b7��5--L���9�U�gQ9�u��G�v&�%�v��l�av�@��ܲ�tJ�t5x|R�h;B3���H�(�x���q=2n�L��[џ���ͫb�<�(}R򐻐28�����[|5��?�&<z�$F��uGh32�����U�d@"`�H�T�����W�F{WRM����ӯG��*30�Nv.��/Z����B	�'v��'�5K_,��|��O�wcӟ�y��r�g��%������t�ٳ���E����F�F`������G` �Ϥ���Mf��x�ڬ��QE��U��S��e�$�/�g׊/�^�!�L��<���9+����M�ܔ�v����݈Ɓ��ע�?�8��0�S��������}4���}�q��Gx��rZN���#�h5�h��!��N�^�mW��|�����B<pp�)�\�`��������I���
E��,��,Ue�l� ��ౌ�H�5�7]klS
�C�.��N�����2o��Tc�~A�2����d�dE�CÏ�Z=Qԇ��M\��	5N��p�����E��xr���׳����m��<�AM���_@E�/t%�G73���
�+��y����j��o�����LMѣ���T#�F_B�����p��4~��%���$�8�T�D�{e�%�zS�<,�{k�f�7,��j����^xa:P�i�0 4�3$x��;�9�~�]b���5�~��s�S�/�!�}M��%7�ɨWo�� ��UzK�t�n��Q�F�L�_�iNo����z�P����e;��7e�B��3[Yp�X[��/��R͊���v���\�rC"21�Zr�n�<Kd���������#cT�"�7��@���t�xϭ~�A��[��i������ǁ^M
ZF��Y��$�f�/�A��cj��$���/_���+3�����|�3|�����mʏ$6�<���	:h&=�xT!xG?34���� �{?��:�ngc�.��VCW7*����y~���TH0t�D=����̊�����Z��X�>�g�У���"UF{w��?9�8)����VY8�{��kO(Ⱦ{�n�R
��]��������?��bWu����8����� ����~��lxGo�͟��HgP$/�5#X���L6n�gO�Wh�R���2&�Ѷ`�&wV��#xI懼{����t��ݘ.�8��𘙮{�~=)�z��-�$���e�^B�-h�xqU�W�"�2��`jn=�e5*~��T%���p����g�ڢ>��!�-�:DmR�.�Ա}˙ɵ��#l��|�1�/.����ɀ�j�q�״re����"өDt���Cbk���>Ѭ�V����TNe�
��������@V��ѧk|(*/���D��
-irYF����>�s[,�V�C��7+g�*�o���m�W>�?�M'����P��G�Ru�N�G3%�Z�j�k�Ó����U?L�p�pl����0Ӌ}|����,��ro�����P?*�'�^������T�g�I�.앙�eP(�=4�e��B2�[�ݮŖ�`>kL].�o���3����=bp���r6�-vDr�5y�������11\o�g���:�������gEփ]���G�(�Q��5*';^�6L���+��ǧzJ��doc����P�&��j^��A�`ݟ7LL���̗�Z�#=��co��2yi{����$�	�p2|7��=�O��M���+e@��>�=o��3nd$���SO����n-E�穖��|z.+mwK�0;k�כ��A��q[�S��G�QMY�5"� ��oL*l���}�� ���U���L=� T�.��T��%�FM��b!{�N�G/�o�tf�6�`wLO��m�#&̬?�_l�����}O�*XͲ�ۑ/>%�����A�iS����+�^��}�����M����Ax�Φ̡֗�+��0Og,�@6�Lק�Yb��>Ϳc�?��:�dW�L�~��RA��n��i�����Ϋ|
�Y��!i�I���Z~@�����	*2���x�����Qo�f��M�i�h����f�*A����CkZ�����I�!D�,�v�u�ϯQl�k�������ݦ\f��Ӭ��.xRd�k��n��Q�{��oEQ0Z�Ұ�Y���w;�3鳩�t�%m���98 ������ �� ���R~�i S�3bBA��Ag�3�0k)�b�D;{� g��/z��"6�c�����t�f�ͬj\���N���Qc�Z�������e��-t�aj48�\5$��s�m�×�H�[�ǤR����)r�g���_^G������13H�}X��=A�?\�~�9:xp̰�e�Km_�Rz��Z4O�~@�:��7�P.j�/BI���&
����3R���`��LS�����'��Zg���9J�u���2�ד��vPۆS�a��h�1*:�������З���g��S�ߞk?R����z��|,��O�3�Y����x�j@d��t�Ϣ�;�v�i={n�H�VVZe�9�C$4��7�����F15�w��=w#3�<4l{��s?S��nUh��N9=������6�[|��R/��׊fY�U��؅r��bc �B[�H�8��v�9͇��,fJ{�^�K+��WQ��˜�d�]��.AG�śfm��V�{��䪚 n��iErI���6t/��؊ڌ�s�/
*,b��@���Z��g�Z��9� �aJ�4f��h0/����'������#p�i���;r�j��A���-�T�Y.`�,�J�i^��8n	p��&�Lo,tq�I�"��D9�)���o����k�/J��H� ��!av2L��>�>��a�m���na�!c[��ԍ[�����⧱�q�-��n4t���}����X���e_�,a�6 J'ˉj�Q��L1���u.���?��lY���r-:4�߷A�����W�	u���IC�4y�e���	�\Ĺ���v���/�U
�Z~���-���S^`E\U���z����B֮ь��gddd`�T�;�DG�F���BU�{��DrD��c�I�U���\�%�>�1�/�E�������n��#�QuH�=�����;��nfA�;o&|���9�wY�Q�qqJ���8m{�;zL��@Xv��5��_\3��Z�d��&¿z��a����s%����#ӿ뢡U���i{���2�I@_��m�+݂';t��w`�_L- �z�d�w�P{�Q��r_��d�/�:�E��yR+y�",eC�f�|� B��z;��t,n6|��]S���4�|{Jнm~_i���ݍ��������H$��iO����u9:�!۴�A�N��w�W���ۨ�P��}�o�}�h���
_�X���q�]�n�
kjEsHT��V�����s����o�O�%������x�WG�}�r5d�n
3����ǥ��1�����@q��wǁ��p�˲N�!I6�}w���;�i���������ֽ�L���>�ӊS
[x�my�i��kpd��T����b�h��A���5�v�W�N��Y�2V2 ѐX\{�l�����s# � Lͻ7*��K����4�ݻ���,����/qgk�����AU)JI�=�Vq�<w�-��YZZ�j����X_U3U������T%bLT��� 	b�{��߽������t?O���w�������Z��ۉ����F�_!����F��ڋ D�5�<�K큄y������A�k�X�:� ��}�o��L�X� 	^��=���ܝ~���v��y�����?�m��a!.�s���D��(
s����!�����B��ﳣ���^m���ҁ���.�cT��Xt�W�d�uo1h��{'	�b�=Z��ք.�zz�p�����=^��6e�dɗ����x����n��:�R;xe�7,���\�^Z<���R��iٕ�%���:ۄܐE=\W'4��A؜�9kO8���ia�:�p��+���X�)�-Ġ�>V;5���:�2�Ǟ��������g�5�����(oa[�2�e������iUdOXpZ����c��?Χ��F���������,�??+:ڀ�$}� (��Pva��2����d� ����=�1w>ӱ^��Q��T_k��qfư��Q�@�h(S����󹎽�p_��bnB��d��qk��#�]��s�^*;F9��`�e���]�b����Rƚ�̌�r�����{�Sb�X��ر�4�)d����7v3W�n4����W��C-wiIII}�+�7�\8��m����>�OG��0x3�������������6����e�|u�T�q���H�9�̓��<���~�lHV#��n��(!��p��{	E���D�L߸ޒR�,2zYY�"�������-��b[�4��)�,�$x_��  |����S�+���+�M��c2��g��d:^��lG:��Sښͥ���q�tSPЦ�YGB��z�O��ɣ���w�F:w��;\ͅ7rWF���_ygX�AB���9l��h�[��6ԣ����\����2�f���y��~�!GW��;>*e�F�=��P͌O,��y��O���
�����2��|�^ ll���q��+�������,�p� KN/1����O-�s}�.�>�幫��긄y�d{Me���A�@�#�1I%���AGW3e$w�82&�,�k��~T��?J"v(���;�����>�����5,�?;*_w�WE{�����US����d9U`�F��7��P�� �sj�G���S��X|�>.ף�����o"�9{����J�8	"@'Uh�j�d�Hu���
&b��k�Y,2?b:�vu���qM8�
�4bG�>[���v)�[/��Z�C��=N}-�ɔ��˭��n��˼�_#��!��&� >ɭ?[o;��|6�`pں��v�ؔ\����<z��(�thx�YH��06�&�hg˩���E��2a�?t~&�*o,��Si}�n��o�F��~�����%-����Y講5Np�qH 6샗��G��X�[�ŕ���|�R���塯��		O	�e�|]}��`g�Y�"�^=�l׌λ*Y)96c20���8g�L&����x�.����3ؾ0���n��k �p�:���t�i��y0W�=�=�z`�'�[^�sSxxԃ�4�����I��KR��O�D��C��^X�����(;v����G7�*���;s6[j���%�zi�b$�l뭴�����lӥ1�4���˱�\O����7�/�jv��ߗn~�N�H�x���Ɂ/���P�󏣱�j(��ҙڢ*�K{������4o<��hkˡR\����|r��M�.'����P�.��/�/6P���dJ=��lJ?�~�~����''vI����E���m���ɩ3�=������]1�r�p��;�U?���p�lH&����ʓ�7n}�w$��'FrAK��L��2�/M"y���)���[����-���w����ݨPi8zSck}{*�d��c0�iq����>i����o��&���Cg&n��|8�W ��rՎ]eiBXq�8��q\˟���"֗���)y�]z����S��*��]�a�!�Z �� N������;�#w�_|c�a�(^A���E�'��,���]�?��ϋ,J���� +���h�#ꨨ��8�| ��;sՊ�ɝ�t���jAה����P->8#V��Sڵ�8�X.v�g^��*�[��T����j�V���S�Z���[Xq~=�Zx�ұƖ��7c# )Kuԉ����M�]��;�U� qҺrXm��O��l���w�|��1��cx�GBZ[|8��Ҳ��������'º���0N���E_.���k�s��� ���Q�{��*�"�t)�X�>�8z���Uaڭ+w��3-<�s"����J�v9g�ɜ"[�F���y+|Nq���d�����"��Â������z�
��WB�� R����Y���^�#��{r����Z��X�����	w����T��?�s"�����^B�BZO�8k�� ���^�c�-�
�=��~N�t��@���˲����S��#X�eo�8��9��O�i{�v���������i��:B��
�e�#����6UW5� h1��_��G����?w�}�|�u���\������{�Oqw��A"���R�p9�/�C��A��2B�|?��z!z���H��O��%l��qe��	ݚw���	w��9�r�i���'j�q�5�|ŨKK��!��	��e}��G#Wv��syj�u�����W'�݁�'?�Y��d>fIa�ё>��X	v�8�fL�oon��
WsW�9g��h'h�Nhzt|�&CN|c`�p�)�l�0t�
ߞb�0]t]��M7����z!w!��d!v�ۺs���j���
<�r{)-�vx���vx���h3�^6���Jis�뷉. �`Ｖd���VZ1���31��^�_���M�;V�4��L#IWӦ���Q�C��}�2��"�؏`�is���_�S��[��by�7��-ܛ�	c�;�G�ƌ�:%Q��L�^^sC,����s�, �V����:���oy12~��A�7�B7V#��J�l��5n�o�.����r�狱5��:��Ư������jG*��8�uٹ�%y<X���Y9ኸ8Ԑ:]�}�ϛ�^�ѽ@Io8�S�4��A.ղ�؜��&�Į�vpK�F�s�7�F�nXTx�?q�%�װ;OOr�{S��ⲉ��ð<>�*�9
\����B��	J[L���m���L�&��*"f�sV'�T���6�/�
_}Db�}��VUN�yNZ_�%�+�R�x��֬b���-h�b������`%�^�c�ܫhO�׵���)���d��j=<�v�����K�h=��7����TV���E�+))9,�:R���y{��������~������2l�>��Z�9�Y~k������t ;���!��#�%�h5p4D�T���8�gl�ٙ����N�8!��s�c(l�"�,휺�kw�鋋�������3�Y������f��\�@�fu_{��g�A��C�1Ym���������B���c��|�����&���F���+��;�&f�\��?<^e�i�ⓚ��۬-�`&E�Z{�o�~T ���L�S������S����'?g�_�Z�S�ۦ���!�����e�y��}n�E���BKwX��\����P�A��Om�>�[�;���[u���$I�����ŋ��,�	.����lLE�v���쵍�����	��\ :�\sssۘi�S�y�pIke�D!�<����[�񹹹��G=S�Tg��X�
^�A��u����I#��,�`�j���(���d�Oie���lz�=�j��9vi���K�%�~o�⟃�&_ow�+ª�d�$�p�4�\�$e]\���g���R2Z����tw�@l�on�E��+i�/��iF��� ƭ������X�Z��\�-��1⑞~��-�Zkķh����~j�F��'S�-B�H�+g����3����%�w4���7���	+ȧ��S}\-�1D���Ç�i�+��2��SF얞���vY�g���ۚ��^֕Dj^B��P�!����r�_��B"��?H�U|�Iݸ1�b��Tܜ4ӓ��/���0#=�h�q�;͓�	�?6b���o�:U�������X��� �ֆ�
��/b<h��3ҍ?�\��;eͰ�(�����jr��̱2��{35f��Փ���p���r�������D]��-�Ӽ*�(g�ջU#)7���0|x{�h��6Q����u��ߘcm�[W:����F�����`lVIcݡӏ^�ӳ��_�wz=�ɰ*�*&$�����{H�A׼\K�h]����!�>����:�!��`�uQ����X�G�{u=�'�݄�:}\^'yM
'6zM�G�������S�q�d*��%]l��{](�%n��Y{"%19����/ɨe�Ú����e�Y�-�]Z�'wS�Ug[����Ud��Z�("���t�i���Bs�aU�{ǫ;���Cpȹ��8���)&U?��%Zٻ`'���voXU^C��Y�{m��k*���ۜt:��~�#=�E-��[�#ݎ�E��9l�a{W(�6��m�Q`B�n�CzUA��?փ��kuV%�v�!�W�V���u�{r.e�y�-��Ku���#�x��T�涗i���1Xo@�Ź��;�Εu�5Ӥ��?$U��3������켎�X�Q��g5��UN��d�/�J�I��e3��w1---ٴ!��0�L�*�R�`�~bZ�Ͼ}��D 6� `���������?O���h�ߥ	_	�OtJ���2��g�k�K9~��ϟ>���BשKP�N�� CS=/��}�.k�>?�u�&�ㄺ���]^s��-{�^�$7D�|�o�����${�������1o]5���$����,N���V��Lkxñ3��㠙&�>�#�]F[m�.su��X%�2Aǖ!6ױڈ����k�>./��v�&����'��yudx����3/Յ�ad��;������5uكx�`�| X
��+J����C���~�BJOs.�_�ܭ$�H.[Lȋ�l�?��q���1���<g3�^~�?2T���i�>��ųg_��O�|��z��!��.`� �j�+;\�7O�V����6���@��Ψ��d��+ŷ�O�����2����M��13<��)��aR�CEƀ��t*�<_��m�W�zW|�v�D���BvN\<������z~^eY�z�ZW
1L��u�Vj��@����������V��Mci]�AAR�H������:==]0�+������mb�M+ۢQ�8��a�(�O��6@ݣ1���:,�8��)��-�����t1k�7ܥ�WK�����n�65�}�E:������h�ϫv^�����{d�F���,����ÏW�����H˜�;����c��U]�	���O�e Q7@�� QDR�<�S�MV��,k�wB��d=�����Y�=�E%����FSKS�k_-/�%��6�ɤ5��S�H�MuN|����|�����!0��{��ZU�u2���I�!�3b2Y<žy�}	�����cAnkC��&��cH���ߖ�W�9��.�?m\�ڳu���r9P�i�fk�Z�-����~1��d1��j{����]���p���p���6:��S^�D+��ݒ�б����{��O��h&],�=`��e�������QK�$�����0��-�/^���G-s�q"(���n�e�*v9��[%�`ɕ% <�&q�9�-|����d�e�!�R`oo�� ��Fz�} �C���9�ړ���,��M�&��K̿}<��1��@(�s5g ڨͼ.��Y�ң1���.�d[��A�D'���U����b��N�b�2j��V�S�:n��fs !��J�ΎA�ؔ�"f�Ɖ�^� �j*1� x�P'�L����dwN\^ĪjQq�Dz�2�?����b���QĢ��C�U8�̟n`�E�GU�$_)`��1�>@�>z�|�dJ�8����ß�orϩW�v�/_��\	�����ڗ��a,��p�8"p�8� �y��ɷ7�^�>F���h�%���������yaRQPp���([?茲c�#Z�Ҕ���5�U���H���-�ø���iZ�Q�ZLa�"�*�����^�[��?lGz^���2��fͶRK�����A��ړ����/o��6�!�y�2d�q? �Y�*!H1b��ʡ���Q��6Xn̈����f/��������٘>��d���bhDL�\�+V(~�c�A����l�)�Ox1��҇�}�Պ)2C����L�C_��B;���d��
����w�5��!�yK�+gs�L9ٲ:�j^��%��<qd���o�e�ڠ�O�k�W隞�����4����lW�3{Z�W8��0sb	�(aaa!��MJ:矧ҵm�z�Ё��X�~�V��_�5���*,j�v�a�I�l=�dw^\��%|j1�(;ᩐHk	f��H�򎸌 ���� ���OGF �z�SL�V�s2�F��%�^�'�)wdr��؉�hc��թ̩Z�RѼ�:�� 4�S���>����́zZNWSS3��g�(L�d�=	��ʟdbN� cW�2��w�"��[�ҶZ�D>X��ʁ�aH�[N��9���
M�P�AFp�I��L�#����'�������%�F|]�c]d�u�D8�ɋ}�������Bƞ�K(�.�2����4,�v2��׹��#�t�;:�U��\;��50ssbT���\��5��-�ˎ���M���6�,�-�r�)�/9��C����L��f��<mQ-cZ4�9�]UU0uݡ!@��2:Pl������B��#�9��Kہ���Q�LajGwǷ��aS���ӫ��sW=y�� %h������u&�ɺa�ư�;7�j�cH�p®%[�;��7C�z�C��j�CÑ�!�hރ���%A�.��+ @BY4Ͽ��$�%�s4m!G�ű&ش6c S�pQf��^�tI4�H��UK'!��݁U�*NZG|R�~0�Ҡck����5��ʜ�9y�%[���xN}�xUy��z��R,(Mɲ H Yؐ��t�7�f����~c 羅�Tq���2>��aRUp��[6t��h�J�r���q�e��� @LD�DP�����,�p!���ڠ���J�9��)?��/?�]�g��z��rc�H�W`8���s?�T����;���	��}P���4�x�ܸ��
�_�w0�-��Ѱ��-����:4R�����,�ф,2��A��;8bb<����<T��OcBU��[��E�sǀbbR�*�Ei�
Tb,;yxh�J�	\u�i�l��=�����{qE*��21�4�l����R��
�p�̡�SN���W�er�f�Nej.����[�Q�� =e'm(�(��/�8fP�M�^rSU��~'_��Wo�� o�B[2�V�F�Ou�n��j�^�{[W���s���HREEE�G�e/s�ֹډU�g,����#�!���]�+���yAf��^LƬ2�����d}'È쀏4`�{)݇�1vS�		re[���+K��)�8�lr�G��gwi�|�1�D���M#&�SeW�b�������ܜ6z��ǳ<�z*���Y��(w��h%0����zF��3�^�CZ�}����<�:���Q��˦�K���FxW�AwRG^�R�����.{�c��� l�%�[�C��hӣ��cPǠ@��2�͹�Y��I�;J�"���V7���[\-�0�]�Q�2ѩ)ȉ�a������^�(��jUoT]�M��z���p��j)�1��~�1t�p��U��ͱ�6~��<ǳێ�UKT�O+%�8��^�1V�;���9��%�u�g��R����z4+�cr���(gU qx���)����〉~�|�i���Dm�rv���m�%"�h����yz�#:>#X�D���2X^=���@#l�f_7	�a���ڢ��$[������:��l��?M���~�����k2���6�x��{�s��a��|N������-E���2G&����Xk��Al��b<���Q��*pB�ޙ�6��5`d�uku��DjT]Jt���pě��h]�,������Q]�<�VNi���v$<{#.,��v��sV��/��C��S\>��{ܮ'4�|�xb3}��c�>��o0W��m�d�뤲��l\����uS��Gt��uei�u7�@"�@;-ݼ�Z�� P��ZWmF�}G�0��-_R������ɓe�ā>��W�3��Q~]��؊q}��pf��pEJɀݖ�N8e��Y�)w��2P���Sd�� �B~X�k�ܧ����V�h(.�gƥ��#P.^>�|��Sc	B�*�K~0''ǔ��Km<4ӓ̓��lo�Bi|a�����|3��CJ�k��D�(�����L�qF	{aBZ&��\nKC��m��]k�r����P�kj~N���Ox��%F�op�ޓG4]]]OW&� ��j��3v��Ī�� o�2�t'��t��T@�`=?�l䔘���H@���|�YW��Y�[q;�X��R�w���I�|�J�&y�᧐�#��$z�f���
�Zvء�>\<t����0L�iߚ���21��Ғ*������6�ACgg9�R�L��p���
�V���J��ὐ���#���'B��I�4x	Th�ql: �v�hC��:�OkO>�X\̟���*�M�00�>昬|W�M�^
�`��I
�OK����}w(�]�z�������a��ё�����:���<u~��Cs�R�#NB�nB��lbF�K[��� �|���ccc�����i3��uuex�T��me���*-��ɣ���_=bp��0&Ӏ��bat7�n�6�4�z��+��,0��c9J	!Em�����x�z�7�%��L_վ"����/��䗛�~\E늖1����lud�o~�N%Q�HT/�Y�e���=*y[C]]�z���$�f ؟ZC��m�-��3DI���>�k�\�˵�?�Ȱ�Q�LV��M� �P����3-���n�����{~�+�;�l�>�OR*�A3�;5K�	ҏ�3�NX㽰*-��ޗ��u�ss@�ad�hK �ttGMLxpodi�}r�boAo_�%9�� ���ݎ��������%<���ee�&)0t��e�H���'��=��e�Դ40X��>�(Gh��m1hW�C��e�{C'w�wK�,��z,����su1�v��f�`Tf� ö��-w�NeJZV�ҩҒ�2A�uŅ� �m2�av��`���v�]��ݮGh�f���1�J�8�4���6�ks<z�C��ʀIw�#�R���_�u��3-������`H3*�� �s"��kġ�[����P��!���:�aX;�����l�ܘ�4�
�NR>�����61�ꕢh1I��{-bc�w! ��\�><���ĕ� ��9�SWٱQ�@�>~�:O�v�B�q�]�}�f�X�yN�y?�ȤSh��0�b��)v�0�v�й/ý���]���\�K}�n�w�hF��z��y�+����ҸL{��]_�&��>�l�
헍�)��{Er"2�_؀k��G���QLSn-�Nrv��X�>	�ܖ(�X�8X�'eVL�v�:��Ԭ�cd�qy���b�O*\�I��w��՟Z ¨��X��_E��nd&U���H�S�#�lύKG�I��Re�|[�
L>��
��RCǁБ��X�4���|Q�|h�8%A[(e�=9=;=&KˏH갞X�vc�:vd���T�\�����P�B`3/���D���-LUh�|0Q�z�cu�1E�cX=�z����um�<_�c�HM�&Za]��-���n6���r]T���(@��C�lNN��r� z�.x;O�wԆ��� ݗԧ
����8I�ˊ1��qj�8$"g��-\11QfQĄDd�e����AK���{ºv-�r��=�(�Ġ�'�cjr��
}s�b�e$�v̺��[�S�S5��b�/Fv�v��ckchY
a�;�t�OMH�7϶<�x�n���У�I��x#H$�n�8�j�{S��׮�G����0��Ε��d�zQ<_�֓��p�ߛ�^G����6s'��m������A����������l4��n��;��ݤ^��+�M]��=Ol���lv�ݬ)B(Ö�Z	�H+NPH�X1�;�ףU��
Zg�o�����ٸʈ�X���k�&P�LS��:����hg�K&K�2�R������������]�4��I�m���4{�v��p����;je�+��H���S���_�|�Z�3*��sqqIV	2y��L�r��Ў�! |%�/�����Ȩ���M��,�t %�<�a��h٧O��JL�@��|���r&��,6�%��$�y���l�[�cϠ�o�p��t��'w<O.��d�$�d`=�WO���H~�41�{39�6� �^��I�y[]����'N0z��K�o�����; �
`yh�_V�x��Itj�#)�oi�����V��`G�xX��j���}�HF*yh[��zk���F��+��'In	�D-d
ɘ�2p�ō�]�Ӓ*'�o���k��|��;+��g���Olk�Fͯ����k[�G��?>���! 8��e}?oe� �M--�G��:4����_XW*L��f��S<�@�v�v���A_8��W��P�	��e��� ��nx��R�LM�Gt0��&vJ]��$akK4��V�k	�1�>M>W?�oa,N���ȗ[�$�2��u����t���M`�4�� �s �����k@���Z���D<����	/�1���{�!�z�������<�}���:�
�k��Lqc�g�j*�d��6��v���,��V�-�][�C#��7�h<��c���c_N��qpӽ���� �(.�d�(M/PlG77WJZ.\�ǂBoyc�?!�& � ������ �/�x�̑:��^UOO��w,����/���]������cܛ8f��lr��k�?�P�Kϟ3]��;E�u��S��H#aWkɧ�)�C��ex��_�o�9'�D�E��.�mB_������W���P��ë����ǚ�`H�9м������|}�(�ï���'��Q��H�@�n�2G\��U@��R��7�G=>,�2;kL?@��*�@���D�����y��o��X\��s�sV��/�,&�k�MZ=z�I�=ڌ6Z�K&��FEE��,'�L�??��n0�=�!7X�!�Sq�?�%V��C�	�2�e�{SFv|[��֖DSAoz�S���~[� ��Z\O�y�tf٠Z"�j�c��}��'����������*[�� � �kz���	yVp��� ��M6̈́���s=r�7>)�J �E��������rI���4{��a�!J���ʒ#&������v��\�i�1${~.%=7�XjGl�M��j���C2B�Ɨ7��	��pۂ\]��;lK${Z��k00�ͪ�<~�+>���`��>ȱ/�ol<��N*N2	j��s* lT���j��U�\��Tm�i�~!�$��Aܿ--nvP�4���&z�
!X|��>s6�\[A[�DV���p|xU���L�#1�F���C(<gX��-���{[��W=���(O+K;w7//+I��޴�1��*[wOԄs����~!p�jV^p���PT�x�>* 9877����٧ �X��!�)c`�uvw�2��hĄ����*����^�}�9���T������;���ʠ�?��Q�/Ⱥ�kuh��L`KR�T&��
s}�F<g ����kY ������o��F��SΡ#�R�Z%���j` +¢&:��&� �s��H	X����5ݰF�3��M�Z% ���V���F\ u9�rqʓdW�IZ��%~5��9-x{���-gh��%��?HH�O�\�]<*gv-���|���ͪ�X/x~��^�B<�Ͻ�����<���mll���� �r�ؓ_R���E����".[8�\p�~q �q��U��� p_����������쳏Q^d����/@�U��Ǧ�� ��	wm� tc��fb�K��aaΡ����!1w�ƾNs���A�P	���[�}�	�I�ʲ��__��9�0���@`�'^�~߸���t��^�	�����Հ ��dlߓ��2�M�\j%B/�����[qv�;��*6��A�{��=��i= �%-���:.mr2���+:�s�� ��3������Z��u;7�o�!ۀ�B7&gQ|q�XS��o�7�M����S)�,�=?%iW������3�D,w�1#*��#�s^F����>�5�=������w�H�.��Y�G���gҷ�5��
��5���sf���h<��k}����!K\���|��=�T���t��M$�R�<�4]��+ۜ���P>���k�H�'�(nhh蔄�[�B����t���@�������+U����Wk P����0�Z���������mit��֙++.�Wp�x�P�6`�����6�H��&%�MըY9�	p��.֜�پ�<TL�"{�
X7�!% ے�lv����*�z.���.��w�������E��@�`/��-�u�B*d�3�0XF�Z�A�^|��"T�HRj/$m���7���qJ��G��V����{*��Գ�U��Ҳ¤.`���tH�n� ؓ=�{�Fh	@�$ �B}%!!�ri���.r}@r�.���� �܋�%�����vs���5��>C��7����@:�B��!�	�`o��'�Ç��wq=U�=$m_���@ �N]\����j�?gO��lMc�[_691'uTT�sH����E��F���.���[�VUpp�c�'�<���0d
� ��D�(Jg2����6�&?M�������g�)�`KG�5A��A��ٳg/����۷��� X��1 u�H��}����d��m;���'�A/}��R����g��
(F�#Ե�kK�񡢖}�@C�JGE���@A�~
�3���H``��i��#���< ������҃O���$-V	�rZ�Hls�F����]�+*�K�B��o<�r���'��#��8����9ԅ�����yŵ��r���2k��Z�W%�n�:y����vI	�ӗ3�����}��\�	�(a��ONA ���;!��v��[x z��l�ƎXɞ������������z���Q|��<0i��<�� q�=�tZ��n��ٔY�&�t�sQ��2(�q��SO81陙��*�ku��� ��&/WU%���)8�xZ��y�TAA���}�7�Elz�wh����ń[@ �2@� y�08�z{�˄�o��j!	��{�5�@������i(�B$ʇ��#*
H��υU��> (�xa��h��700���I�u���7p=2o�Qy���EN]��8z�� |�iY��P:r��q���Q_���ߌ�pV@����[�[ǋZ�_g��✿��gq�
�]]u ��^8��vf_ޘ�4{%6ށe�p�s�h SYL�B�O�	�R���U�h�B�dl�Ȁ���ȁv���
Ռ�������r#�,���4��n�N��RpjN��Ȉ�8���\2�Zi��� e��� �\+j��#���/ndiy�������|�mu���mqQ(	����Y�w��P���3Nx�a@]QǀHq��>0�s���L3����L�h�
�k�N��\k�j'ra9lХ����RI��~��'����4=KK�SP�D����^S����R�����$
�i	�9lݽ{Ts��������%йccc�cc��Gj7'�;;͚�8g�m~�k�څn҃�ZG��h�Q}��Y� ��Z%�q���� �.�����2�:oXs��_o�5�zK5�"��*�~���h���t���037'fiY��V��K�� )f�Z��FB�ԫ녅}�5�1 ������h��z�]Z>?���"�ݪB�
j��9�v�N������8ۢD\LL�M�� ܋d��ҍ���3'$>��'ơe�����J��MVό˽{����8,8vdn�.,�� �F_��P��؊���yz<���2�*�y�ݙ4��E_[K��۹��(@�f����d$d�ͥg�&��h�h�V�?�o�o��yv�lC+� �&�&��� �`�ⶶ�M����O�0~H,�u�}�w�����2�3���NgR��]Y���bb��:��*�X�G�;��O��OKL��(�d|�4pQ�2��� 	�؜�r�t@jry-Da	(]�nAq�B#�� W����[PV�++�{k>&1��L�U6�cpr`��x�i��ʧ���]] ��T�Д��	��;;�;��[:W��z���q7�����9����~ke�mu�J��=u0�mheNʃ�8�Ϗ�Ӽ��;2")��C�Pf�d������|�T���h��f��b� �B�VQX�{���w���T9�7�-�tuuuvu=���*qi"c.=�Q�ǀ�|]4�g����Q�� ���=䀎�h�)09�bՁ����9klbb\�e@:W�KH����੡��C�es��C�k�Z'�gZ���t���s��B��p���@?ɼ��'�ɽ�����q����𓘀ܑ��s�^h�
e����[مa(F[[A��"J���;4v�1'�w�$����!GG�O2x<���4�C-�<Imz� �ݘ��|�G��*��S1��ś�Y���q�A6���o�x�-N�G ��?�З�k�EP�.��ۖ��o)�^��$���l� �V�{�n�gcc�{S*�4��(#Qv�̲��W�LZ�Db�X��]������|J�����L!u��Hčl7�Z�G蝨{��?�V��з}NXڭ�{��{�s.�~�n��˾a��K4�XZ\b!
��UH��T6���5�-����B-���Xg\+��t��Iw`�C�M�H�Cqw$Rsu�,e���V4�Ҷ~s
�^�h�ÐX�s"��$�`���|x��k{���6����J�����euf
�͙2�pɎ�!a; ���`� 8���&p\=(x�Epx���Gi
�;�z8^��������#����'ʱ�OojhpV����MgsvX� ��4�T�������4���H��-;&�� �)M:�����N��...���B��'+�А�=k�j)<��tD:q-���~��G�1 Zz��%�C����:�-���,�j����2$f_�9��cK{����Db��~���_�
3弤�K&����RR����M�g�fu��m��Ub������`e�`i�ɫ���}d���P3"�wD���ǩ}�Af�h�Ņ��&V�Q�o\Q_EOw (쑽�3,�������&��@q��ɚ��K��R/��~�n�����ď��snd��|t��J����H��iU�W�e�z��Gf�0����ҝ��֚�O
@�IQ�퀔k48#jn�<�!yv��3�c+�P
������$�&�5ɯI~M�k��C�Dn���I�?KM��ȉ�6����k�5����_����k�5����_����q �Cb�^��׶����_���xS/�S�v𮻫�R�/w|�Z*�,/-~=v��כ���|��|�h��w�K������/��r�s
���,Gp��_�9���{���>�o�7��~���:�;���޹��	~M�k�_�����ˣ�9�áwL���	f}�@ ����������(�Kٛ�~6��3��֪c0����� �^�Vh[��ZRw�}]��d�	�K�a�B �2�A���A���5�X��z�R�K�!}\��ϼ���6^_L]�pΩ)�M�a룷6�n�|H�
�Ļ�#{�m�Gi�̌},C���`���c�r}C#���?"w����aWO������$9i77���3��k9��f^NB�������"vUm��Tsr7�]ܐg��`.�G�w�6��}�I��.�n.�r	Ț����=���bp{/m cO�z�ԍ$�+�IO�
R}� �蓠o�q���¶L�L�eU���M��&�Vۆ��9oxZ����?��ق��Y�Z���cle��WD��a�8#d�S'l�����Ѣ�zD�rgXŪ��4*�R�m�WȈ��h#OI�]S�U4|��?�h�6�E��q�#Z<.W��FoϮ��Z/48U6��	BƙwLE �m�V�y�3,fz�Q���1�r�����&��޼u��aͬ.�����尡���~h�F���>�i{�;GmOGA �������k�_�4�����7��"]Y}[�',�]�P^V�u��I�M�?���E���4g;'�u�:�/�뒟��R�C:��x��劋w��PK   ���Xy�kWq �} /   images/d23d5e93-1caf-49a4-82f1-46066b67b28c.png��uS���?�.��݊k�ŋ��@�P�X!�[qwJqM��K��ł�S\nޟ�}��O2�ٙ�=�%{�+RS]�[YI�=b7:���������{EY��q�}Zey���ّ?Z6���k���6/��e��|�*>q�[_+)k��X�V`!�QD]_���L�}�|�^�~����B��թ��"�1�ތȦ����O�5Q�K�S�q��D<�Dz�<(����	q_�gu�^��i�el�iIW �7笨I ���B��m4�����	��&tyaB�A\#��>��***�GFG}���<'l�1&.��8�4.��7P���o�Ƚ֚N�L~��=Ttz��Y?9��i�Y�C�}y� ������{s%�Yt.e��(�~��y �1|�[�}bzx��	PI"
��x1��Y���q�<�=�Eq$��i�����i���Q��y��h{kK����r��o��&��1��Z�۳��L�q���6��<��w�����R�Z�����!�o�O��^�v���������Q�µ�ӭN��ޏT��CH��Ψ�OM'.-��(������� �ظ�_�q�%}����������m��f��˝�ߥ�w�w�?��1�=����c��M�Q{�a��%{=Ҏ-���5��˝��K�g!,��t)��&��+*`O�K�?�v�X�'���m�h�Q:t�~���V�<�8�����
�|�~tuT��lVXhrx!kD��Rٴt�!^�&��u�a*�8�ƕnP��ԕ����-Q__?��pn��G����F{��@5<l��.�9�5L��\Iߡ���Z`p�L��#�]�9X���p���.��B��u��?�XpQa?v�Aj[�k�������	q�ʍ*���.��'�46�����NN�����)�#Z����Oͯ�ו6/���2@��,;���uw{;r�w�)�'��>��9��02�?|
���$�0�5I�@J�����soӭ[a�P!z�����p����_r��$�y�sґv!���j�n*v8�GJ�@�(< �Wc�>�F�7Zj�o�&e?����5UtywZ'�7�Kf�۔���M��IA���g���%�qrﳵ�=��MPPЪ`(E̱�m����[����J���䤅����ɓ���ps�sn���ڤ���f��mܬ�w[��U ���~��r�@���(3��vɶ�	B���;A��mVS,|�:�dRI��ƆD��_?�A�M ^�	>-6�z�7N)4��� K]R���������`�j�����5�3�+m�t^�y�>�Bg	[��)��~~�;m�Y����+�Ǣ��b2(���oP{�(�4�������c�P�����(����©}н��[zyݻv�M乍��V���N,�[S$��{�� ��FK����\��x���������&�<��7�'N3�<Yf۠�!#�B�f���ݣ0C�΀����"[����뛞?� ܋�#�f��a�~ͨ��t�5�r\\c�Rx���s�vu�b|4��(���x�qتe�a��~Y����Dn���8$'#X���?��~�R 1yk�`@��>#P��j%r�W�ڇ������t$�̯3�%XZ��m�sM��&�ch#�^�temɥ3V�m'"�Z������J+�k�y�ێ�]�uy=�>YMl���T�q���AB��h;=�� �z����3l}�5�1�@]g��q��o���.��Ld B�
QV"d�RS7�p���

(B�ˬ��g�V�������T��2F��)���/��C�z�Ok�x�g��q�g��5�]��V��W�Դ���G�y�<��	�<��WL|q~��y���"9�W�,_��[PQ1Aj���;rK���"&�����X'DL���ai����NKp3�%���f��C����4E�^�fa�'��K�����������`P������MJ�_��k���!�=H�PYާ�H� N�޸x�Bå��}W��_�}��2��v�i���u���9�#����v>n�Jx�<��"D��a_�zp\�_��>Z�3��đ8��G�p+�]l?��f+�lm|�ޣ}�s��]�ӛIr~���0{�:=dg,�z�
���r&g\�2���z�(���"liUj�}�˻ܝ����~�>4�$m<"F�o]<[�����u��e'#��}�������3zB���+�����_Y�.!�Ǯ&	���6
k��`��ZH��m@��bNH�;�d`M::��&�I�Ym����C�*�y3�(���F�����^Q|��ߙ�Ԓc41Z�AoA����ô"s�y�>�%��t�R&����J�Mt�����6�5��������,p�� �*����>~?�IU���ą7p�#�=��ʽ7t&�<�B��q���'%�����K��1M�<�e3^�]#���r�qZ=K���7���T9���"��̔k����fG���ܽ�f/�W,���n����o�cޔ�^��;6��L'$�R�D�a��d>U!�ٽ���-�������t�VH��JLJ���FНzI�_Y���(�xh���M����'��s��ל�u5z���@Q0*6A�f+�XME�Q�B��E:��-���ex���!�;^7��������r��!�:�t'�*$sXK[!)N�[�N&����(2Z�4���T�����۶��р��ѕ�cR���`Y~�k����^k^7�\�bs��h�:Ͻ?��m݇�$�>��$��I9��
�~���ۘ��8�P3o��VS��Kn�B�hڞ����d�����|��p]ň��H��
��0���tZ]CC6����s0Ίl��oi�]+�#d��j��{����n2L�q��7��UC.�g7�)���.�[�B�]'��΂���Wd�-�Jz�QY1�Q��t��i�, X����v�8��Y� �y��uc����������L��r*�Մ��D3�W�{��vl�������+~�jV�/�)E�z�3���-�ϒ��Oʰu�g�_i�X�VN�͞JOί����xШ�mɆ��GA����TC��Z�)�G�-?��)����S���������K &N��x�%^�>�8~� ;�A�����/�������/?�*we�ӧ�9h�p�rB���3���s�[hwJa�o��$i1M%�w��3�}Λx�~H4
��3����F��t�f�t�%�׻���'w2�G�"��S�$te�?��!.�l>'1�KX��Hƫ>^\�A14����H���I�o�|��c����3o��#a��z��W�I�w!������j�t�p���tb��J^8��L��;K��X�%��M�v���\7�����ѡ�-o�l(s��@i����"�l3�w��F�ͥF������)�9~�?]�����/U��>�'��7�J�-�`�~;�����n�$"�1�BIK&{M"���;�\�1I���:�6�G)u�����p�4k�<ʎa�{���������EBB,Ө�硹N��d/s��j���:�k�앵5s,>h,	:�mX�I����Y.�i�&@N�ņ���;@�mˊ'E�Erzk;�r��k��H�bf�Z�a�����K'J& ����i�2u�<�!��ۉ���0���v��d�Kɗ�K,�J��ʚ!ex�j��M�D�F:EC����磘͐dˡ_�Sޜ��?��sB8����s�8�M�D�s��!�q�E��]���̭�DM��0�n�v��R�x��
�BR�o�V�b���k���'o�I�����\�U���9��[>�t�Z���䞲ex�$蜓�xٯr�R9�9�D�������^��d�X3����x���jx[ !�V7�R|����h|����k�teխ�٘f�ӂAqC�)N���I�M��u�%'�M�/9�1E��m���P�k�ɠ�{�Ǭ5�R�#���������J���mo(B���b,	x]�~���\��\0�=D5ƖK���P]��1��ؼ�]#�W�]}�q���oWv��RC<���2��4B&�Y��*>!�J��N%����,���`%Q@�z������o�b��Ii~-Yk3���~���F�Md�4xBH@$j�X���ρ�r��?�pщ���
�P���Ѱq�_�g��X����{fJ�Tѕ�oP����K)w�e�G)	����k�u���}��z�I��	�~�N�19i�xD�W���n�Y�o�cP�H@H�n���z;�'�;�j
��=�h��T"2�]��%�^���f�͕/X'��H����[�@�E�8�D�M���syP���<�)�Mm�Q���]p`��9i�bö����s��D�}N��kQSi�_�[��e F�W� �� �+�j_#��hx'EXY����z�H��m3V��4jԛRJ�����y�m��QP.n5�?;Ca���
�!�IMM��30`���@a5� I��XF��y0�t�����p��-�'�uD ��&hQ��):"IX*�pn�Ű�w�X�Z���V����6E���<�����q!pK��Y�x]ű�D�i2����HJy3���X�`�2�{�Ӥ��ҫ���0rֶ�Y�|���?�$����fy˞]�ː�S�	���*��}FaVkR��x�̍�8���M��	!�����o���9�-�^ܸ	%��Td>ui�����-4{ �>�R~[���<�r2�۶- 盙-�WaDư��$�@<-=,�T��}�{�2������qJp4D���</�r@�E�� f�C6�Jy4���ZC�s0GʨD��u�lTO�"uK�o�J&F�!�%b%����!A�1�z�>W�炘oV����@�M��~.K����]l�N֙5�h?��� U�QF�|,���W�_��)>�d-"��Y;b��.i��[�����&���&�Ω��?꧵Z����9;"˂'��H�(�&Ge'�������a9,��{K-������uF�c�!��sRϯ����j	��g��o���S ��4N��i �u�
8�w�nw�����4ҍc���#l|[ʊB��|��xY@��`#rfc<W����D�[{s� v/,��.��}fv��6��eS]����o�_�����EI)�]��O�FY�x�\�΍�U3��q��
�"�3g,h��4��Zm1�Q��=>�	-��ˆ_U�7?%��y��=-A�?K�s�X~�/E�Kd�����MC"�9Gֿ��\>��/.+�}�wpT����%�O
<Ґ�@���J����[5f��F2�E�%�Z�B
� (�r��D�8���,!ͮD�գ� ?�y�3��W�M:SDZ��U��>8&�j����f���M4�����-m��Z�;�GӬA���иyD�J[�}p�Y&�Bݹ�P@"�I�
?qRpA����$�_㹿K�9�,`��)k����sYH�!����L�Zd׬�"���Y�B��c���v�	��a(�yY��ߪm� ��� �RRR����9'�@v��٢�}�, ��!��i�����Tsq�&.#k��.��!/ Ē�5�т�,����ˈ�e�=�R2�8��'���q]"`#F����p'NrJ�C��*��G	tZ��q��%��b�P~��;^�����6�e�-�HD��"��k3������\4qO���a��jU��Ѝ��[j��C���@�h����������%$��[�ݍ�I�p+2TA�2-&��9��HgvVF�o=���a���5[��&@x�L��%go���1�Ć�o�s VB���~45�ۍ�2�ns!��y�>��5�ȫ��b�+UX���Q�"�G���n��T1�Ae)��$u�SfS��94�c�%q�^(��ݞ������X����ѼZ��y;}1%f8r�RE�X�C�'�R��WY`o��p/w
)��1Š�|#�?c�1B6xHk�ӇYexM�&����6�Y�R�m�f�ز�q�@�X��z��4��}��J�#�S��bohh�, �2E��n����r�c���ӻ��qD"�
�DQM��@�5dS5�#�s��Or��R��B���B\	���C�c�
0 ���~h���"���~�����Ӕ����D៱@��D��o5��j��XnN�_.h��,-N�5��IV�tr�h�-�\�W�ϻO��ǫx/��ɔu�m'��>����*�uDp`�����G��K��đ>�	���e��O���-���l��%�r��<qT1�9��yU��I&}���K
c���~~��s��/����E�����Q�}��~/�6�w���5��q4�;A:��W1G��}�Q����5��|��D�W�&J�7������G�q����O��~��+�'��^�?-��?��(W�X�~�p��c��}�a�rS�e�2�̷H��<�m�}����5�x���"�����&T��c�+=\/͟c�;;"��~a�y�2U���b.��V�1UP�{Q�./��LE�@.�d�(8�W�%b:e���W�Ng����	��Z�T�m�����Ua*as2��r���Z~�^�+�47���B�*�J�1����w�kd>]٠Rٞ,�;9�M������k�4�����)k�_k`M�>iI&���a�Z�K=NO�e�⾿$�
z�2�Xv՘��tmRD����g6h�� H�ݡ���n��1��Lh���g&�((Nu��(V|�|��$�
? ��5:��)���>�n��Wy)�d��Ք߯�q�F�ri瀃/����.���������6�"��^ux�a�n�
2�:)��Г�I��(nKv���$fr��N��&C����\�r���2�N�B��� .FS��SWj�!�4�����es�!npo���d3��y�(�n�����>A��T=�Y�
Λ5е{_;�]��1ƌ��6��O<�@�8$Y�Z+L!1�!4�W�R�q��`_ʘl����5�j�B�ӗTA�\N�vC�R��6�,�ϟ?�Q�I�@�(ȍ``>��;J�\��0\f�1#n��u4�"j�Ev�.����_� �c�i*o��Ms���۠!�tD��A�(��9�gxÔh!�bI�}0"�
��E��ǯ!�¶ف�FLh��G���;�v��2����z�\���ӻ����1$���A�HN�$83�7g�+I�©7³�c 2ifc���b��"��˛�V"{G�'	�b�����Q�7�G�/Bq���P��>��cϻ��s�
�ά�~z��Q-!��71�a�Ya*�@a���[p-؀�+�*"����']��b������_9�0`�b��F ih*_z�m������x�U����.u��"��Ҩ���R{����2����gyHHe#;sD5Cme���R��}|�!�FE�Ʒ�	��@�<�L�,����7�ŅV�+G���,�8�uIz��& ��_�ԓ��΄��O��bЛ���vi�~E����	PQQ�w��꧍�����ܳ��? nq�C���ig>e{���9�C��7a\������+����9�,T>��E)z0f�XRu�}'Q�����U$y@9�O�BIh�ui��$���+�?�v�=�Ѱl�>#Q��l��X��n�ۚˋM!q�o(kZ�B���Da�f1�&�Sy����b#�B#��t����M��;�<dџ����Uǹ�~��y��C:�e�i�-Kvpͯ@�3�=<"�A*�dW���b�R&"����F�Ŕ��!e�@�c�7�}B<V��(\u���[��me�)$:Qf��EP� �)�d����fD*��U��g���=��:Z��>��R������?%$8'1zUƅ�f�*۵e��_������M��P�D�N�ΰ��l��[%��pN0`�G0��5$tS��mzE��h~����K�Cx�܄��lKMD�{*���8ҳ�
����z�^U��ta��ج��J7�;�gn<,�v��S^6���Z��s��;Ư�n���ھ>\�z+m�{�(d���a�~6w*�sY���-F`͛��bo9g2$�lֻ� �T��A�!���'��5�s�_/{���K�2���-�u���`��*[�ֽS��H���Bl�n1�K�'����M�8���OB�#]oX����R�a�i̛(���I����Q�{�����Fn��=w�	b���-�8�>�~�6G�"���K��p'�O���ʤ���~{l�lGHb��m��d�K#|���~(Qe�|���6��z\���*�wl����W��[����Zƕ���D5iJl�PsQ�Gฤ# �Րr����2�)j,Ա�\���{W2d�	���UQ��ʌ�.D�۰�(\�Nu.X�����Yٵy<�=����e:�p�2�Л���`'��ּ�t�s�#jp�}"��G�G��+���ae�Ç��onO�Ы�98�������w�$�̢�Q�S&���+e ūk�8�j\kA�Sm^R����+�IZJ����mU�$Iˑ.b�Sf�I�G� vy*��ut6�.�Ju����oa���%���� ՙ�O�>p��X,�:D��$yҺ%���9�};G�e���z�\i9U��.�+���ӧ���E�PI'�����%���L�n*A]hJ�L�Z�Ȧ�5CJ�J�z�D�2���$���Ȋ�)��J�5�u�A,����8�4^"c�ѐ-W��ty�v]�/$�UW�{SwP��$�ȃQ��w����t��P�h�oX~f�IԥL3g52?8�_�@��|k�)&���w'�-}�QM�cWLP���ǌE��}��V韬g�L'��x�~���8E8dQ�^j���� v|nr���n��2h?��X$�* �ณS�Re8J�ǅc��P=N1�Snp��	�Q��i# o�1�,��1�;b3�н̡�F�	��S0�q&��Ǟ0�~K-����r7�63j�M}W�mP)�m8�em���\��(�.� T	�`�U��<�h28:𾖄Z� �8B��C���wZ���Q�`x.+���#1�5�s4�ô�&���â���
��~��g9rh�~~�<�10/O�����9W���a��n4v�m���9zG��m'�C @�<��?c3���J�������	�U��B#"r�!�ۂ6w�e��P�KW��Cm��|Xa`_e��J՛��"�֣�3V��p>�r
��~���7=�����Dڮ�1DTט�]ܦy1�v6�Ck��˘*%��B{-R�@|��Yd6��6Ϟ�D�}��z�%���k�����\x��~Z+�%�B����GR�ϵ&8�	&�<�9p��=�V�N�x���ix�D�^O����*����xӇ׃%�0=Y���,l�+�0@�I�WԢH�8�� \�fL�� �d�@��!)+֠wi�L���[3Tr�L��AzH�A���6��(}�Ȑ��K�0�;����p���+χ���yʯ6�u�3aL����Dt)5<ν�7m)V���T�d5z/�lf�����u�IgE���NgP1��F��I\=�3�Y�wɅ/g��
OƵZAl�A�h��������/x_�������S��BX/&{��/��Y�Vg^z��	���Ǖ$݉��� ����7�s$7٤�ݘ*��N�IaG�vpP{6M|�����lr�F��G���ݷG=����j_������ �����#g$Ȉ��]g�n�_B.!O�n	�&�}��������Q4��8Y5�KD��I����E�������v�-8�)�a�55��<2q�D'N��!$f�]�]����u�|-{4+X��r[�K v�9n�*fxy�ښ(���Hu���	� !�o��)�p�{���p���]Nr~��� ��A�ӝ�]I�ӻZ��4fn��U�?�PjU�?"Bw�Fyb � 1������z燫-E��:Wd�iE�b�_I�����:�a�����������ϻG�a�B���إ��RNYՙ�9)��˘([ײ�`M{��֊؊-Hd�M�ޣ:|z�<�<�w��UG�C��">	"a�"B1u���抮.��&��	�0�5/�F�z���!��	�6����ž�ʻ1�(w�Hx�Ճ�h��fU�s45f�Ɲ2���K7�J}w�#������wq �p�R����1kt*���U�S��*!nh�G:u��+�72�`n�f����X0�YD$nG���5�^��Ҏ `#�҅Q��a;��9�( ��Ԉx�Z��#��>i-�2��ŭ�b�Vk~��LW�D�;j�����W��b,�Ɩl���+@���t>�o���QQ�O&�p(����Ի�V����e��l*���,ٱT~i��R)󶱯uc.��~��\�d����T8�V�(�bh'�w�(HrW�r1�k����᪓r?���B���w� �����BQ���u���$�@����r%�|v� � �N�`����I����[5nB��B��|�������B�\��.�d8�(vL�Ɣx�4�L���0�p���-�I�훋i����HUJ��:���e� ���}�Ex�3�S%-_�2V5��t��?K�EWQ���,|�sS��S�_$\�q��_0�����U\d؎�@d�{'���se�j@��!Pe&��'=nSh�?2D�(�4Kr�YTUJiD.m>N����{��e�f�(/BU�^mW�n=]�A��%�A1��
ױDR!�@��tG��sqr��Y(�z���j)�l9g<�!�v�M��
�0#1�~��B��ߙ�V�H8w?�1����vJ}J7V1Ξ���%�g�����	b�a���oL��N�JÀ��l�
�{�O|��W�20����d�R~DԌ�W}{qT�ZX膱�v](�*뉣S�A���2���:.���v4�:<%[o�P���ْ��M�$��18��ȓE�N)��L�T�����dR�,7�G��鵎�b��70������?�p��`Q�|S"
N���oU���P�"/f�O��������"ɹH��JH�ӗX�d��nzs��1��	��7����'���|l�23�QJ�4h��r�2H �$����8	K�������
2^mLuGL7�$����  ���e9��x�O�炍ib��-��D�7X��@�6�	~׼M(mFT>X3G�եW���ִ���/���#�b��#�����ڳ�wmi���h�8q4��\Pj����o�~�cvG��a��5�����h�?늖�k�=�IJs( ���H}�g�[D^�o�(���x��Ff�bOtH��b�����A�WE�W�+_n�?Q[;�p��{k�\�{���@T$0LD0u��?a��D����h ���'e��l�{uHH{��������A.1T��Բ�4z�4�TG���^t`qZ+W��H�����L��0煹|�rg��z]>Y|���db��@�| ���O.���^�td�N(Y�2��{P"H����8���8�U�=�)�ĿrF����4�z86��Pio��Gth�.W�r��E"E���xp�>����Q�PMr�ݲ�>Z=�$�{��#Z������ӯ/�&�kEK�ꨪ%��]Ȓ;�Xk��yN3�?�$S� ~��1�33�u���6:�S?��c��)��,�����3�y n���q�je�4�{�c��ᨎ%�o�^5\L�QMo�3?����bmԶq�ar�8ZNV�/��p.��(�@@��7G�/u�ذ�-9��0B\i��{�0ƙ"��G�4�\(�jW5���vZ��;�W����=S@We�l��� 1F�i!�}�?�N�abeUW��5�LE�1	|NZ�ɟD�^��c~BP�Qf�no�Sb=���d�q/����D�׮�R��dG�Ӟ�X:?���֠f�b�^T��(�(*�ڢ�|[�ST�oL0[����U��jn��BYq����#�[��$�!�N��0%�xa�J���P/+�q��S�v�>������&'���B�(`�_�Ńs3_��W�#��%�p�`
;c
iޣ�>��g��x��{I��"�ǌ^�7b~���^�͐U^� &����\/J/�y���D�A�<_�5�l�"j/�YA㖲��'i�x>,�����eU(C�>��1����k�0�����tf�Y��w��C3o�'K�&o���aX�к!�?I\��+��ۥ��\�J\
l�ѕ5���_A�ݚ?�ۖq�y�j;MS���nf��7A�,=:&t�  �kͺ����/��E�?��dCwLv�:'�DLCF��N���;��.vE!ri,ea��Y�D�_w��E����"Mt�\_M3N|��Q�*4)y^��M�gX��.6i��ԓzޣ�鏠^���w���+bф�i���HI�ڹ"�Gm��+�6�����U$��<?Zr��A�17$1	Zm�߮�G�vb	�Z1�&Q�d?�T��ea�j��Pk�-U��X�����^U����b��j�����j|R�b���MN�m�7b&"�?g�g���O������T���(��E��R~��WJ^;�i�ں�1�}&woe�Eݱ�>m��S����n�*;�E��)����(1?���މ�uw�����Xpb2�۳=z�8J4���2 |��,�eII #vm�С
겶&XԷГ ��k��Aum@��1�7�����r�Qd��ov������[�=�����y'!|��|"������DD���z\jv���|C�<�X&�#3i��9�B����w�J�J��T�7Ka�.�s�Y���{�Z�6���2`��ܸ�Ӊ~��i�G!������E��AHf����l���ÖVD	_��>�$OĩrE�o�����ᶙ����I�iYJѳ(�͂IL}~�Mg�ݥ\��Ų Ϫ:���y������z�]�I��1���x���:=�[���������j��)k�p 1�󇕀�;�/ LU�<N���Y?�--��D��a$5���U1�?�KY$�`:M8-�!���,��t�!=�� E�zvw#͜oF �1W�/4� �>��`��ɬJ&MC1f\����֗�̹|xr�G�Q�U����\pܴ��N�!�}���+SI`#��$�3�,;��.4}�ik�4j&j0�A�C~�n3C� ��- k�0Fh�!i���:s8^̈́��-�֫�{��,��'ńq�Mhn��Q�k�36�R�#�$�=7�4�+�P���( ��@<	�1R,���_�(չo��X ��kɐ��#\ֿ����a#���)�t��?퉶�D�k�4�AX���_ȷ��4�]�l �Y#T��<���_K�� �dVU�e�D�4c��O�Ǔ=
%҅6G��j�;�ˍ͘H97�	�VI��,��?�ä�he������o-�Dw#l2��%Q��1�ڥB�v����0W�&���[�R
is��	�(/|�o�M3}c��M�*_�O�eQt�����x�%��PV�3l�x>��_����)�?]&�k���⋇�-�]��=��KgRicF����M�	�2hi��|$�'�����?E`<��ΕL&Wi�ǧ�V�=N�^r�w�T��g�Z�,]�-Z�i���f�%��&N�x���=KK��kX�֒
9'�R��VگU�(5ߓ��ÞhS�X�"r���$�s��2՜P�VTX���i���l���h<_PWI��\PtM���;��S�6��|Yu��~ό�g�I��;��X*�Ɇ�*���/{-��<é˕g���,z�p�~�z?$*�wt"p����_��"��y��W ^�!]nx�[X,DS�5&Bm� ��n��������(��w�jIzҕ�����݄b�Ѳn���\L�Õ��9�r�	���HM�Zt׫��z��ȢҞ���u\{o�@k��!&-�O�7�������c�I6���
�C��j����C��W�׈��5M��8�z*~�X�{�S���L"�^����6�����.�Z�W�Z�N��\���8�`���W�>JOO[���UJ��E���vD����VYt���|��?�t��.|:��� e���)�	xބTx!�Έ�����
W�jq�q������o[M�T�t�Xl����V� p��	�X�cHx��%�6cN�o�;�c �$#���%%%���2�dU$�ĭ}�С���i��ջ�"N�ҔzHy.k��/Fl2�n�:Kw���J�W�Sf��j�T�h����A�6�~fA�R�D���
�T:Ry05l+�&;B|G5��Z2��<����9�_�����:����q���T�e|�z6d��陛ס��PFt��Gy�]�c?��9QrЅ�3���o������̥�� 4�#���O�^��I�������B���5o\�,O<=#��ƻ����	�3�T��#hQ6d�qb��!�zH�c%<K �J1�好F�cT�b�O0B�Ϗ��_Y�/�FFF0�v]���BZ� �� �i�V6�eR�����R�)����|즏㤫4�M<]�K��?G�� +��k����*]�f�'+)u�<�~"N�6���&���g���_ �VΆ�Pj�>�He_b�_��X�^{�J�7��IM˔{&��?+�%��x6�s%K����q8+C��b[�R��T��r�=�����߷,����~�вF���|���XY. �/�(|�ZE�@˱�����Bz<��O�'�Yx��&�,�!�I~��Fq�?���]vy��hpƻ"�?��Ƶ�w����%Җ�5Ďթ2��c���!�����s\��K�TKP�N 3i��#f,����SbȼRSSW����������[h��܏�]d�hg= �4�;�XO�#�V%���%qU�>muð&�3�|���r����gl��C���`G!1���}�����x��v��7��>�W��\'b!�{P�`f�}���Td^��tҲ#�3�����K��/$��/��W���,a�*���pƼS�M�������E�~��2�m]nz/�M$y�f�����d�a��G�d�.��[-z�8r�
���ȉO���^�Ѯ��8V�L�,����dFԵV�8Ii�x01�.W�G>ׯ���P�!5u� ���ߣ(Q���W�|:x@����g@��*^!�ο��k �Ţ�\.��Ѽތ���Z>����r|����T�LJ֐�M_0L�9�y���6>)!f�t����l���Oj���)��>�~C+���%]�
�B-zq�㢂���l|`�.7J���tYgP&}���gm]ı7��R��$�!����Y#�e�(��� ˨�����p\1���jBh�@ƋT'<	���}�L�&�l4zYǝ��͒S7�H��wt	��D�Z���]����
�L]%C�Dw�%�~F��	��F�7�C�fmɣQ����9�
z���'�qyoio��Ŋ�[��޿)VN�^ˣ�ڭH�`Evq6(���K7��jL�5Q�Uj#�	�킷�1�U�}L%ǥ�E�6���seA&zR�Z�Yt��sU?��lҕޖ/�p�L�P�J?P�y1���!_J����2�AF)h
�Z���/R��>8U����������m�.��F�8��t	�,���{�q;r�!�YT�'ml�I��|�=z5�z0©��O*���3%��E���$�R@�2���8*��LV�ߥ���0�n˜��ҷ�����欍0�U�cA��h�!-T�+ȃq�q�����A��(N~Lq�>yP9G[�~ݔ&��A����R�E��Hc(�.'��Nf��pe��Ka�mc- |�����R���*���(Ò<�tdL?����jU��=�����Sd�\�eF-]�KM�[������ !e���N�M���҂�
0gb��{z'�z.-!�c�C'4��x�SW�����Szz+�� ĝz��/B|�u����F�=Ǫ��;�i�S�	tQ()j>�J͸��(���C�����0��z̲Ҹ��ڎ�,��O�_P�J�r���˧�Qk9��m,uu����4�7������E�Gm�k�ּ@L����<y����Wâ5D�j��uᘃ٩�mI��H�/�9E0P*8j?^~�{�^'���������']�����dĻ*R��ˡu�l���4�/��-�y]�
q�p&)��:���8SC���gQ*��I��
?-�,�6 :8�$Es��$�-�3jƫ�͍����b���M���u�z������w�W�OS�ʖ��'��5y`�"+[��\?ʓ6{��W41Z��p2�bG����α�Q�P����BsT��0ظ��;`.�`����M��|�;���8�G��Y߂ ����;�g�K��۶mۘ��Ķq��ęض�d2�m��;�~������]�U]u��C���<����ͅ����	�BC�C��.i��'qI��1UZo	�o��R����l���Y����_�0=�faWt��Di�mL�fv��X,#ҫ����J	9a�a��;�{ޙV ��]=�8��x3XFvlO��� ӣ{T���wQ|��&C�/���]wo�(B���,��n'6"J����=��z���jK��L�!`����*���>f�tm�SqƯvc�-�:�@�tB���t�S2�7��Gw�G��=�:�a5[�w����֓oU�?B�O�Fެ�<�{eU���V���Z��ʑx�|(v�y�PZ4x�5agrκ�e5���U+h�B!�G���C6�N�$;��H�B���������M\��9�򐷨e�@�����:q�	Ԁ�>�RQ*�j�C�Nf*8�Q1���B��_$�F�+�B9^�����Mٲj��^n����eG�[7�"D�=�W��3nHq���ɤ�r��z邴��ܸ���Bc�j!�O.��c�h�c`������O g+���t�����Bk��vR�X�����g��L��X;��g��|�ؠ��#%��wS���"bW�����3�ؖ�x6���X���^�fn���`8�}fē�0����YJ���#RU%�/?�al���
xl���t(�&3��G�2�{��Z�`R�=J�.%g��8D�A�X�G�fF�_֓�����[o[�����n ���,f
�4���R�B����3EQ�?~&6�W҆���\U��+����a�}����j��ծ�h���ݲcbY�&�� ?�\ N�/U7o��h@��w���|0�ȹ��ؼED���%�W�d���e<,�-��3)��Z�����1���Dx9~��p{e��T؆��e�f�ǧ�t�t�#UK��?8��_�VU-s��%��(&�p�+ \v���8�M��׫&��.\�(��b��tKڵ"���M!�P��i@R��wET�2<�s�!�r��r�V$���t"����F�.S�˳d�\�+U��o�f+h<-'.>��0�J�Վ����f�z��'S�ю���Q+��/�"����`�	������F����Z9��Á�ĕ�*��Lz�"�!L�"�|O���W����l ���}�����}���s�󠣻�]֍�������\����0��rs���ږ��X�Q+ò)8�E#��2�7[a5��W�a�a��̴�9!�e3HQ�)�*i��Ř��M՞�O������$A@�X�de��K6��I�"ɠ���v
jQ�D������XV�c?���̒Q�7�-L~e�(�8��)�� ����5��F~]s��]�t;NY\�}4 @|RI�?��)#v��8� �$�u���t��%����1;�k�iI=E���m�u�id�3M�H� �9x��͹�ΆB�����`&����`�T��@M+��Ӆ��*4���
����**��;їe�N�E��'3	`�x�$���A����h�xc�_N� ^PY�[��m\�٭�	�_(�Rj"?c�k6������Ѐ�ˆG|�A攒d�al�<e_���\}���S@|��r��eBg��1!Aw��N���{y�SnHBD��M��Ə�N�[�g�������y!Y7��Z��܈z��8�R-���y`�/ޱ]�v�
�J��15���|��GqȠ�=N������,��K��� wo߯����-A�VKY�m9�!Gp*�rݡ��wp�qaꆮ�b#�}
�7گ�"�f䩓�(�x�����}gKI	6��N8df�dA��&����.��-1w�^C��10���5��r�_-�� i�!�۞p�5�7'�ۘ�'���$��u �ժT`t���X�!YD�U����)�/o-Ĭ�#��T�^\ ym�	�5\���'�e����-As��R �������5���]F���f>����!��gb��_a�65+ؖb�5��r���TY��~1�xD|�$d`�C\9ά!�F-r�x�0z&4�_����:⠏Ѥ����s^���D�!�Y<`E�N�����^^Q�gJ�fΟA�iI�D2Xͬ�������Z�듹DEh�~C�bv�.�"y���$H�G�>�T��On�%xBn薿,�F���#I��;�I�س%�ո&��-ڄg�S� <��P�Jj�-#�Z��(F�oUh'5e�&��tѾ�-�^�y%�ެ�m
�us���X�H���o�:���k����Yg�ru2.zM.fA���+��!�`;�X���F>BG���ňA�辄��sa�d��x�gZ��ZW�(�����<�=^w����'2�ޢq�ϭP-]}�ɍ>�|�*�ֆ�c̖��P�sN��:Qb4�ЯQt��s/��d��;z-ꃻ�a|�l�&���z��wʻ^a=n�|$�~�6(ô8+eg���U R�V�f�Ɋ'^�(��� ����__/���(�й�W�S�R[�Z�BYA.��o���vo���lqyw����K&�N"���4��f���b�ظ�.:%�jT<*䌗�������P-7�>v��nw	���7�.�ܲ��� *�c�/��ϡ����������Δ�BH7����H�����Ε��:p���	�����M��N����Fk���%B�[#o��}�"}��"�����,<N�iS¤<��<�ގ�iaQ�4�]�茙m�0>ޅ�uyE��Q�o�id�x���.�&Z�&Fp��a}z P�-� |����R*�LW���+����2rQ�|x�#��V3N��􇁬r�j޾r�{��3�q9{�:��(�#�"H�����`DtX���NX�9�?N�����B�:0����aq���uLZ=1��B)}]�u�+k������^��\P�y�=u�X���@8�CA��FJ��,��z���D�.F��@��qH ̭���}^g�J� j�]>�̦W3�{-���&68�v���`3�!s����,���c-�'O�C�|�]�vㆤ���#Qe�IHiY;��j�G0���ʧ&gD�ı��G�Jb���P���@[�45�(�"�H0{��pr���[w��v�>ϣ��!]��C?ա��,>�t6����6BQb`���HG�m�`��E��P�z�6u�ܠ0�S�G	�D�Lb
���=�IH����ހ��w�8�KR ��L�r8R��xfFJZ�j��zE�oc��6?�V;]h�vvy <�b��|��it��G6���R�xz/��W�|�h?6:�,��'��e�
vJ�#��J5lt�5~t������H{��hG�~��`6���f)��O��>t���Z���f�ֿ�h�]�����	�xf������bj��s:.�7S�-X���� �!���g>�ڝ�v+��_���(��\�OS���iҙ]12L��bu�*�!z��������n�~HL��R�Z�ً�K�\q�ۏZ0� ��x���:ƨaB�q3�d~0@GC[30�5x7>s��L���y&Ѡ��}���8>�21ٷ� m:��JԱ7a��S�ڕ��z?]�w�����R�Ӧ\/�(�-B���!! �t�4y�HQ��wuk�p#�C�'_�$��!�;�2���e⁪���s}�v��n�ɦġ�1	����E`�҄���W�s�ʝW!K; *=e�f�b�8�Ok��q;�v@?�r\�~��r!�v��)��>d��(0�� )�~��k�	>����/1Y��z��\g�1�<�3�v���^`@o��_"���(�dB�Ah�r��kƖD+�f��K���Ъ��[SQ��X��yO6ug�k� ��S�p���:��;�P0�N�HA�g>��'ˮ��s�¯_9�(%�(.Ek��8���DYݺ������`�Ϙ���C���#1�FU�1IhQW�f�ne'[?��1>�5@�_�!�L���5����<7�v\!����16M��H�֜�gX�߸�1�~[H���a22�E\5ð}�m��'q��'����t���y��;ʮ���He�.ӣҤ-�h��e�(�b_F���YU���>Y�o@Hޕt�yl�\=Z��Z0r�,�xl0�<�����G44��M���ͯŸ�@n�2�1:Q��&�/]�����xpb�`�����9#�k���?r|��)� �DB���I���v(�X{}r�7AwS_�g�s��x����k $�
d9f<���!���)�p��0x_�W��v�f�M��.e���"oxq�j��Y}��^>Q]��!���r6^�����:�^�o���<s�Đ�� ���KO.�b
J�!͜��6T�z��GZ��f��j</���(Zmo\�z�X�<��;��*�P�lo�����(�=�8;���ku��xr���b���Ӛr���I.?W|DRXA��ip�ɉ�n�����n�������V�� �&dV�-
&7n���{��Z�\�7����sbÅ��$�R�"����I.��A3�<R���`"�)�*m�Ő�c��2�S�Ź×-�^��G�V �����>��J%�$�5�z�U��a%)�ܿ,�w�&{<� ��	p����)ع����%��KG�S��/��¶��x�y�~޴�j�@ܬ���>�X����$�%��g�Y�R}���:����(##�I`d��e:�a��x��l8z�̳�QߐN���M)��F��`�v�?�M���0�#s�N\n:��~�i0h��CF���f�pZUc��2�K�4��┅Eå�̳M�����D��o�;����lP�y��~�U<M���h�`����2Oo|q���rx��Wv��{�/�"��CV����Z��A2��[��]k���|���rB�u���⸴�_����b�cq&���'��$�dlEZ�rmmM���z^\�)�C�/K$q��9��j�������/���s�%����{#u(A@1Ú���%�8_�'�Cd�>���
Y�I����ˍ�^���.�}PK��5W<���:m[� ���h1���o{���:��S��������_�T	4�7�}�h���a%K������M�m�'�����U4���7�l$�vʟ�m��F;R�'���GK�2[���Ð(#��U��gB"%���#�3������e�z�S	c�*N�[rQ�4���u����B��qZ���v�� �	e{:�Pj�?{USU5x���TC�S��D4b�v��a�1��r�D��V�F�D%c��N7E;ݢ�L�����i��QC��K7��'�����~����>��D���C��B�h�p��,9�b�!�I�ҠF?�F��8D�Q�g���c�%��,B(�������Ȃ��~l�� ��Ca���\�N�7�x<*��k��v����8}�ρ>���|-�����gx}������@�z�+Mտ��#�yC�����Kɿ@Փ�B3���J���P��;��Aw�G�Ro!/�F��a 4�uF�G�e��q��qS�`L�C�!�d{ӑ�ر� ��)y{f���C� �E���П 0k��%�*$G�jlfIH;ɯc�/x�fHF�"yc�9g��Z0��G*nV�Q��gEbZ���76
/c�c�0���d�Lq�hx���Q:#�Bb3�yP�8���#�ۮ����T RpH��?S�]bb�NhM� o�޲!�i�Lf�$0t4@�v�%�TX��'ER�JNBkAӥ��p����;����,}��l9��GK�bZ� <��yq��5�PT�1J.31E��t�z?-~"Xh�~l��~���D�-TRQ ~�r�?h!�̣T����'V˜�^P8����/Nm7ޮ}w��}^�E�lΛ"�k��R"㪑v�\��oS��oA�F�J��/�o��Ͱ:pa�2�]Z�A׼IE�C��aP���jdo�A�7s`��3!s��� {�s�:��A\���jɴ�3K�Ǘ��#��ÏD����,)�`ZwH�q�^+7sw�X5�ku�	^H<T�xC�a�Ld%ʭq�qoE�tv��@b�C��[w^���`��Z�M�BD�X�~�<C1�$=��m����[ )h�~������/w��.]�_�i2s�K�3g�8L�Τ�q�~�r�_��\e\~�^n��L�0T5
��?��s�i#��Kۏ&b/�K� %ւ
Po�G�t��i�,�5?�'x�U����YT
���Q��n�Ғy���fU�hQ���,>�"�;����
�����V��e��ƣ0D9}FZh���1C�|��#hB�Xeϛ4=�	�^8'�C�-9�ހ�F_b�ο �^��Ť��'W��Kʹ$�t��3F4
D�P�8 ���u��E�+�)6�RP"%*���?�NapoP!�/�1/ʬ�r@�.o��*E\�n<��x=�O��Ӆ�+�ϒ/��2��|���J���3V�w�
v|�} *��o$��@��㞞	�Z:MC/��iX��X�gw�J�Y;�-=��@�E��>ry_|ygW�4<��6A|���R��10�	̪�Q�'bЯoA�\�>�_V,XwLz��қ�%lԭx�l.q8��3��LuL�%C\iG�<��QN��'@�'8�k"�h���9���QD�jkr�%@GG'A���NvW��Ü�w9x�8����%9m��U�Y���D�yA��}�������*~$�-��	Z��I�" FB�n�����h�#lܤ�kY(^�c7?}4�����\���,@׸�����@�5ب��`{�J_q���wZ;�6L���MA���
}��W�_��K^c��t�Q�x��ɕ��O��t�y6��t��ņ˶�>��Og���sݩ�疁�Z9����zy��.��PH.��)F�+�S��{���i�ŷ�s�8I���SU��﫴4��
�gџQäs��)���?�)��	�w�:T"�䜈�Khm�\p@�=��D��*I�eT���=��k��罄��Y��u���$��unh�oO�*�W����A�L��Ѵ ��[6z>�k���T���j].S�y��<%�	~	��R�ak?jȖy�C�P�������.Ĳ���M���Y�&0���X�Z��� ���w�����O�e�|��x�K~��S�ۣN���&��2��S٪����������MnK��_7#�Y>���Ƨ,��-��H#-�ᖝͭ�U����=3,���V�٣��������2L܂�&)Xc��-���_.�8NdX�ĸLI�=&��4#��:sR��0\U�Zf�O����RysP�S�y5��RX�v��D��cYB=E�BdjG!�_e����Z�)>�7������,�_�U�:T��B��1���	@
l�%I�Ww�`Uà�����Ul�9�)upp-+CeUvѥK*�Ք����m2�f���Ijl��t�� Rӱ����KTQYYLz$@z���sY���#U/E��3�l䃎Ö��[�%̙5h�����s��z����V�D�H�*ï��z�x���Y��Q�ٯ��5}m������Y��pO�%KKpK�T3iEp�)����ӝ,NpW���E7A�4���a�QiM�@h��y���i ���2��%B�&�g*��*�g{Xd�t%�Dt�qſ	ZT��YU3�OKmJB��n�z,Q ���y]���:�Xc�%Fn��s
�2i�|4� <s�VL9����n�t6��.KiЖ�	��'i�x�8g)R��4+�Vܱ�p�˥��EY���ef>,���Xn,BR���Q�<f/Gq��[T�=��j����0y��fn�F8���,��5���~��X��u뛁��)xA��լ{���|��b�^#��L�	U��������zi2�RV��nG��bqˮT��	`]+���Q�{���-ۚ�x���������m]BN����˶X-WVԛ���^5��M!��Rdԋ5��E�^pKQ�p zZS��>E!�M���R>x:;�\�UBZm�j�}�+�M&�f�u�%֒R����5�c1M�!VVS%���ovL]n2�\S�JD��W�@e�����3D�m��2�U���(�_�
���"\F�	��`����h�	ID;ǹ��wMא%�L�2QUEK�Y��Z�k{�yG�X ͨ
ԥϐ�����;n�C�N/�%�}�]O��]I1�����L0��X 愨J>�^.o�dY�B"�!`Uj��C>cX!�9b6��v����ǳ�������1,�&F�z�t�XN��>��G�6�35%�i|���L�5�o�;Rf��2��*������,ӕ��%�2>��P�ˑ��������/͝��9Jxl�Ui7*l^*%��!4��ia�$��aB�r��ڍ�#�_�h
�c�o5��~'�|�c�tCBPVY�ɠY���#ǸE��N�GG�]mDE+rJ�VH~�C�!^�M$!�@����յ�ci2�';Ԍ��2 T��ȭ����`����}B{X�K8LM* �B�H�C�q�Z�El�Ccq#]J�C��E���>H�̌t�B��"���I��]�N羒�rlST �3ۂKXa}Wg�FY�bR�=x3Ak��f'ԛ0��dkgZ���sƜ�bh0�x��=
���X��c�(�K\�xg0:u���q>-�g�鎵I�,�&q2|O~c>M��+�&���q�A��Bx�@�d��p�W��Ks�ο�����+T1~"�_Wb�u��rC�H�('�i�厘nm�~@åv�ze��6�距?r�-�?���꩹4�7��/����s���a�ˀ���_�w]fַQH�W0V��D�*���8����n�����Js#v�ߢ��n�~�^��aF#047������m�h��O�`6a)di��l7���;����Du��Φ�Ԉ�/k�W�Feە��I�jδY��x<e���Š@=��G���G{n����tg����:r��n�1~āV������+��~�oF�+�O6қZs6EZy�!�O��1 ���z����4����gu�C��c&w>�Qh��-d�XuaZVmAAj�������4z�;Q_�Rh�!Ք���vM]��F� ����� &��u�����E��V��V)F5��Iqg�<,'��:T���=�oZӋ+;1��� x�ID�	|o�>|��i�]�G����T�G�od��09v��I���z����@">�B"7iE����D����|T���V���F:�M�Hmͧhz����|��m�O�'W�HBMrD��HA�ZֱG�M<\%� ���C��3R�+�u�y�yz�����]0^"���ǌ�p��)e���f92�����9�U��j�Hҥ�TN��1��ߦαJ���=Ŭ@�y���6��m2��*Mi�l|���f�l8��,[�-u��Y�u�I�� ���Q� 2��.X�Ea<*�vF�����%=���u?QC����9�:�T
%I6��c�s[���ҙ�e�q��篤g���$/G����xӫ��S	��"Ҿ�r�bq��c��N3�J��9jR�q,=�"� _�T�>�2���4r��Z띃�:�S�0FTy����m���[VB�+m�O�m�o��PPz�i�q0F��F���Plt*��OA'�� ~:�9h��G�{�_�+�+�p��X�O\Dq���!E2`�S�+}��Q�ZP�G����,Y�k�v�����0�_5�;�\u��*~KTL�9x{V.����6?6�������ӽR����V��\��i�on������6-���מ.4p������34ok%*!�h$8��ŭ���$�����e�ffn�#�1���Q��{�G���x���ze��i׺�ֺ�\�-O��2|`�<C�{�6܉�#�� ݖ&U���nf� �t�~�&�䜲TM��͞I�!��M<v[sJѫ��JwCJ9�֥����{��{�ڥ��p��������(���a�	�3[h��z����|#�APn5Rb��+�����ð-*C�_�)>�謫�M��s!�!,��W�	C�o�]��Ki�KґeS���Kkn�+#ʛi��ˎ�/��	���]��r��	����?�
@O�����GS^�bhq�#3��e�r�]�����a�A�1_�8b�Ü�7s����2��&�ꦞn"�k��ު
���>e	h���̩�頊X��N0��+>}�7��#FY�%��.�������ZLvD4�7���W]{�?4�,��G>��)�"�P��L�90I|t3@�=��hL}�iK�qd�dG`/�$�Lݝŏ	~u��*�	���B�g��n��O?�a���W�6N`V~Ŗ�,}��3�"�����N�0
�t���`a=�@�%+H�)��F�^��bhE\dQ�6�X5���x���ctq���o��v�\���q��ẃ��P��c�޴pvb��7zۈJ �I$DDZ������bI�D���vG�K�G�U��'�\��S��<ja�N]y�Tu�t�X��.,�G����Z����T����C�5v�	XL�B��a�P���nm޸�w1P�l��ʲ�"3���Ajt��AO��[�Bu�t�-��g(��J�+��8�Q����& �ԴM}��s�S8�W=hB���'+�k�"�&��t7}���j�ǭL�J���9B�������	2�d��X�~�=N}�̇|K9q�|:I^�)-C{�5�M��ը��Aj@���0i��
6�w�����s����FC^ǻ뭛�k�F+7Q8NS$Ь#�11�[Iw��ǎ8-������l�������J�@[��:@�	6��~h�PHG�C�p��cf{�`c6��}2;}`�<ǝ�↦3;��o��Mr(3��Ǝ��kXI�[�G�v,ѫ�>>�Cp^ShrP���Y�0vH���(��.q �֠�-�*t��1����[t}�价���u0�.Sa��X����B���-�B��Y�.{Dg��_眭wTi�;�U��5��M��Վ�i�$�w"���Y2p�J&v5�Ճ_6T\��BP�cն���q��LQʹogN�O�4ğ���Dg�x'_b�B�p\7QW�����Tsjd��j�n��w�e/��$�Ւ����:	?�A�@�c%�V;��=�����}�"J=Oq <����Z/\��r�'�ж�BB<&{Sb��L�����"sD��Y���y`���r��_qBm.����S�E���rb�irp�kf�ʇ*���uD�my��p��X�ή8\�<�ݿ�rM�&G�U�z|\�7���39Rdf���l���:f�>�]8@.�YCXiy~�ن
1��1�F`���x����OB�؁}hg��;��Ǐ�W"'�9\_�n�f�S�Zr��N�jL��}�� C5S>�z1���i.*Ź��`�9�q�nI�����}hF���㴿�i;���Y�S�����Y��^_n��m/�30_��"7�6˦�}���35a�1�bɰ}�(��c3�/{�X-�(�Ʋ�T� պ��3���&�z!�^s6��Ɖu��"�*  L�@��Ԑ+�+��v<cV���v�z��Y�+F��It�`m�=���ܨ?�%�)&��rE��s�W���N�\��!.�ʉn�0������R�(H[}�sn%�q� 8s���I�/5����6ʯg9�6/�.Lf�,U?6��zg����G+�ZY���ٳKD�]Ʀ��r� D0rX�Ռ6�D� t��Ew��-�'�No���������xЩɩ�!��̙+4X�5=b�2t0��t�c$P&O�5������~;�2M.y��u�V�G��h}��/�/@8%��ݱ
Xku"�HvI�y7�R�ہT�o� �����ZA��L�d�$9�r��c���%5"/@��+��/<�8�e繊6���8����hz�f��������9�X[:��eC����m�SRy�M�Pl``��qUwA� Uc����
�nn�MGI/�)�����k��A[�H݌7��PlQ� �]<�M��#UӹQ��/~~��(x���uw���~H����T�R�%p*r�/��f��jԺ\;6�a&��W+�ٗ�3�����X?HPvc��y���(Jh���mgC)����P�L�bMӀ�V���A��"���
��نF�cC/�\��wͺs��|���쿱����ɌaI��I�P89�}��Hy�лb��6離���Jk�&�Ϭt��RTW6����ܟ�٠5SK�R�e���iė�Z�+CL�_�߁ D�w��j{�l���UW���U23R_�0os����D#J��T�F���_���#��C���!�@��Ʉ�9Nj�M͎�͌ˉ�6���� g�ޑ���*�͈9�J����"�&e��i5~K�j�ȿ;,3���.�g�\]S���X�S��//���1����7���=��s��R�A��ۀg�Ȫ�,QEy�D��9F��K<�&0�׍f�F�_�D2�4�� '�W����Jj�y�5�G�H�'��]�?�͉�*&���u�I�M"n3Y��}pQzC����0֯���l��IW�p��D�]q�!��X�������	 ��s���[����;z'�i8�8�Hm��D4���Δ�}y�ҥ�s|wD���9A���I�;����8-F}L�����#�;��JWC�l���\W}h.�����:����C��+�$G���:,n"`�0[�>�E�9"-��x���l�� ��젫��~����R{i\�حH�1b���em	6�z��0b",1u[�	L�Ra����SC |�����k�
1ǽ��~iJ�v+���8G������:twd�E��vdA4:t}�$N(P�߮�#��>p,%����*�!��r&M�ƻ�ї�^P��^�B�S�h	4��%��2`��7�U��$_����`��e	(M:w} >�	1'�e_Gs���A�V�����G��Q O@��*u3��ʦ��B�<��l�aC,���p���&��ҵ~�윚nP���W� ���G�R��'qi�8�n���i�La	d�V+\@z/�yn��@��q;*t�k95�ox
L�u��(����O�i���Ǘ�Y6 @����xP6�@�c��с������f5�Ԃ��^�8n���b��1v���2c��h�pӔ��[�z�7�dkk�k�eBށ����i�w��9?=@&Z�;$����N0����c?����o^4?}t|t7���v
��<�/I"9|@�6B���āpmΖ�:\�����y��z�52�/c�ԭ'f����`�0�p����-fq�E߷�]����`5�I�T�;{8��Hɲ�ӽ�x�5��K$AF�����R�4���u;Q�?��\��M
-��8�}5ȿS���0#W��, �	&��sC`��4��5�}r't1��f$�����^�4�V+:���o�^*q��Bخ4H]CX�X%�p
&��G ��m�ڛ�^X�Ӌ<�ϊ������Ƃ��(����M,�ua	���]Է�S���bD!+J߽m��qW��E�y�_��Nd�L�[D�m� �$eSv8���p�6Z������>��P#;L�Ͳt_ϫx������j����C30ո�U$M����"	rs��	���~v8�q���S��iL"�$�y�{A��Cqn�ɜ�=tV�tQ�/�,�sfZ���<H��e3m�%"���.?�ć�f]���O|�\?���9�n��MdM߷��%��B����h%�4f�ڹ��:VN,-��ϭ,O�YX|�W|7��"^��=Vn�D[(��o�sS��P��{@��)/�
�����B�r�}>���+9}�Dߌt��k�X��6���ST+�ӫ3 U�������df���o洹�6V-�� ������e�.�o!4�f\I�C-n)�Ep�/�$A��B_�K^2쯰s�b��Ϳb�)|Ҧ
��>��B�{���0$��~�,�L�
S�Q!�r���(����F��#T:����S����l�K)�K=�Ŷ�J�Sdblt�Rm��A*f�t�B�;�co���=]�s!��DT@�%����>�,8�;Nɑ{?��lV�O��Pu��zyA<yC<a��,-���Q �2��y��]�ztѝ\�qT�}�7��O7	�������v#"M]�㴚��j|�x����+�S߳��b.Q�p���e}W\���J��\p��:[�`�l/�9{LE�����
\��Y=�ۣ���U+�J�=l}��$��=!��4�vס�?���)5�X������9��&s�>��&%6��ݩ����%���G�5���f�7�Mbl�rBi�c{&=/8�:�#:}�[l-_��'�؝��
�-}�F�Q��#N}�4����	�O�(�N�uE1u��HY3�S������B�8驡�p��s�Ft(��k#��;,��A5����?��oGM>x�}U����M�����ghT���4��e���C�蜄�u���v]�G�a|?Z]Y�=֝�^��;t���gc���D�k�ʉU`��H��hlg��jҼ����&, g�P�|f���^M�P�k�u��
�'ʎA\X]��5�6vw%��4*��f����p����vB�i8��G5�K��q��Q6�G�
,��l4��rl�|e\#������X8f�I��;��Bڮ�`�֛�z�{��qڗ�am�m��`=���s��
"p$&M�=�	�Wy&�q�,zߝLK}����4_)�H;H�u�2{ڋ��訉��+�p}��]&$���4�a�rr���zD0� ��ؚ��%��t�u��̉�C�E���{bjЊ���Z�<�2�3%m;�R��.X��K���MJhfN{e��M5h��;��h
���AyM���{�t"�<��l��p��j
�Q�l[����م���$:oYU���<���Mi(��C��Z��a��P�Q��������}}� 9�$4<Fy�>�t_a&[�&�&��u_z�@�g�K��� �b�5@��T��C�ƲI���C��]��|בreq� �s�/��	7�@��w�E�$�h�ӉH���&��ٰ""�>�0#� ���e1�H�-���,���$m�����s^�+����	�`�2ʈ!7���8��x��u��H�Bn���|h��~BO�'7�����9N��3��_s'}��!̸�V\�,��ۮ�\H�s�Q"����7�r.��]�t��NU)Mt��l7fC�z�����e�L�S#X��H�y��V�)��Z��Ğ�	d����dҙ��^[�cd�'�����gfew��"`�2��s�j@�)(7��_�����˦��w�D!��D�Q�tE�T�������m�!��vC�ަ}�+ؼZ-�0ς����O���F5���澦G^'����l���)e�tF޸L�W���-���U��[n��O��|A��b�p}wZ$>��`���/�w�v����l�P"����m���dc�{�؉Q�8WzEy�o�����č��('aG�#;e��ŕ����%@�Ԯ���;��4��*�T�}���nZ�+/�?��܁?�0��_N�����*FC�?f�6�@�Ǉ���\ױ��$���?\��+1֩���-F�b����Ȫ�.���a�Y���4Ob��?��H�����qG��Y��,���kwW��M�)4��r�7q�Dio�If�1b!q�x�Ÿ9��N�C���d��Tr�,P�0JDf�������tn'�~J�-F�ő�c�Q���2�$�{(s�w� �ߛd��<y&G���uZE�-ʰ��k�Zh]��ԫd��Ŕ?qG�nS��ܟ�fi󁺐��l{yy��^�� �M/��!{C��|�a��dL5��%�rX�ۚj�����Ȅb�F��8��Rƶ�bi �����P^�D!���l�*f��LHm���V3�F	��g�|�R�JO��t��S!Vڿ^�L�m%w��"KY%N�W��Z��H��Դ����v����n����ƌ_"3�>�ϢmM��s�)�cAya���aJ9�K�F�
�1�U7X.5�\sn���}��+N��v������@~��:,
��KaTԋN���V�3$�=�H�.
�6�K����3lٌ�;2�!��
�48v��_�jj��ҊE[�"����]mX�Z��T�������Xa���q�E�c��`�UW�SWV�qTA�'�DzA��P��F��|=�O,'�Ы�6Ѝ&B!@3ja�I�6(��f
�e�����M ���9<��b����%-�x2V���dSF���'o�2{��0z���3�y�|y�u�|�����s�����/ř��$��.������ء��2�w>�{�"�6�
$� J.�Q�)\:�@���|��={�2�%Y"�Z�s�Q{I�QI҆�܆���6<�Ǝ;�h!�|�N8����=l ��艜n�SM�,�*��]�]�VX��㨯\
��(nڌ�?}��V3BQ�4d,�W�s����?cɝ�‪J����-S��pW��zaSt:��8��s���#� �I�c��_^�}^���;��Y�f���ء]����~��d�0Z(�����W���0?�A�Lw7���_�%%�.�ۆ���پ��7]Jk]W4^I�m�!LF���]�WT�Q1��k���pZ2)N)�	j�0ОS�`�Zw���_<+J �J0~�X�|~�䓨;	�<�G�]z��
�@Z���N-s,�}V	�M���s�x��x��`'�3U�-�pŤAԽϮۆ_��V��J&A���@�-�:�RV�l[�>�8j���1%bî���ZL<�|��Pٵ7
�M}d(�D!?������o���=0y�@d�<n��.(=#LVK��HEF�V`��!(�I�;�9��{�y�N����Q��m���I%8,Ղi`̨��`�@���Sq�u���ڣ;�z�J�)O��o�qߨ@[�cK���_�:�x�-�q��cqT��h6#x�#�Ѣxa�\����ZV�����z:����� �
�7z�`(��+�N:��=�n�{%8bĈ-s����?��7�W����'���i��X)����ha�%o��K��ᯪ�_��t��ȸV^ڋ���6�8G�{�|j�t������t��[w�_��)Z�E��h5�xk�N��@�eC�(��{�#�kOc%�#߸�_t*��0n��;�V�A*;Z���`z����{��!��0X8A��N��cŧ��tE���e�0��� Z��8�T&m���Z��v3`�@wT��X93*��:2<��m~|�4o/�1����ƿ��vn�E�^��3/��o�5���J}��l����dBS����"�6�X����X��$*%��������qp��h	|��@��� Aҁ�h����]�4wf��Gax���cGC�Q%D1_��Sq�����qP��p[@�����Zl����i�6�\�\p>���#�{�s��8�gOl�rPlfh`��⭎U���?�j[X��X4�.��AQ�hg�����8%�戕�IKbL�n;1������o>Q��Z��'����jO̗��[��Y����H'�q��5
qʃ�(%(A� �m��է�:�C0�#��J�.|��)�ܫ'65�b��A��Z���&`�6\��TOڡ�9x�F.
�/���>�ۯ���w�x��+��oh�6_���л�A�@����B�0E�=��Vg���Q����=�B�p��8�ow7�}�Zk� �xR�1/��i�GS`nY���77f,t�1S����k��ȳ��7f߃u����E��TT�r�4z�`ڨ_�̶-��1@�}�����`t�-�"�~.=���Nb醭���+;!y�<:��9�=�$�@f��Vi��L�a���� ��S(���b�7�aqP�b�F,��)��A���`!0�؜�c�E�ñ��e��v�g0��3\����-y��gq�M7���Њ>��t;�%o������8]�̑ @g����1����0�ܳ��ݣ��o?*Ry>��+�={�������vh�mm��}��L�c��\�C�_�W��k���·��APQ��P���Hڲx�f��)Hf�e%
����Qf[3��0c:w��\7��U�cT��$0a���1�Α |ݐ���-���=,y�]�:Ik��B,^�>�4*GO��=��R.�)8zL�a��N�b7���|G���F�5���¦-���,�^5���0F��t2¢Mq닯!��P�D͋+�P�o�}4�:�o[�����`�sء3f,4�z:`ˎ���5�b��gᛷ=��.�����^�lժ��۷�8��Pq��q��5�_�ϼ0y(�P[��'�E��uh)���b���gWʹF�'�ߑ�!d�3�(��ʸ���2
c�,���QcI���}q%x n��:�b�L��9݂��`����٧���*�5+���q��ç���Ǽ{�E�FK�!2,�w삞C������^]�[��M��O�цN��*���ab�=�d�v�H$��?vvh������7�^����o���k����	�a�a����"_B�pq�p��%xi�:����|�U��6b���5�:���+�evC��F���0�gu��-/��ښp��	�أ64gq�^�ڡ'<DZH�.Df�wa�b���/Zض�_t:��� n��
p-X1��]�b|�YT����?���~Hy1�;Cc$��\	�����0�{5,ؒ Z�HX�����k����<%ov�.�<���	0죒(�`�U嶵���i�	�GL��1�a��|�퍍���?�t|��GPݥDőDbWA����rɚ��w��1�0�oO�V���$l��	EY�o���dgiO�vt�Ec�l��V"hk����X3�)��a�&����ɓp��7�,�F��U�X�G�3�0@d&��ۜ '~�0&��Z����9�릐���j4Uٷ�¯��-�X�&�\!��`�qK��
v��>��t&�}��2����S��W`�@p���544|�_�l�'����.���h	^\��B���&�jV�t6qef�sd���-g6d�E �²���3� -�����0��+�6���y���Z>-��f 4���P�P=V���Hdv��u����܍[��]t�ҵ���c��ex��gQ;r
���_�v��1A�uڐ���Z��%i`b�����iA5i�6$���d��xe�[Ht�=Q��,+���m�
�q�b#4�F�'HbA�Y��9Cǎ���.-;����f݈a矆�o}���$��=����1}IӨ�-y��"�(��W��>��;w���=ܴ���^�U�M�4�W���	Ua�qV"�BŖ���Ȉ<��	gL�	��)�`������{�X�a�p�7`��a8�[a�2x��M		N���*�3WʪİC����IuE�;��3�o���0ӆE�����;�턚�$�Va�Rz#
Dfҕ&
D4oH;�G���A���ط��7,���[���_544���A��W �q�a0.����1.5�� �H���<�Hd�l*�D!��e�2�c=��X�!
��U����D�
&�R2A�S�"ur6u�l�s }.��Z�k.>��%n��Jt��.9t�2F)=��QS��G��K�R~����(�2��$T  *d*:��f�`�����Vc���^:���I"$���N`�J�P$ h"q���m-~z�t��ᨣ�c���][w	?�4\~ۓ��RA�\Ha]�9F m��qx�X�1\�@���yq�aT��H%�A�쀜I(���%$�8�2�>TK2Y���8c�L�L�#ƌ��(ۡ�bS���7\�[��������穚!!�4;`�����/��]��U�;d�Wa��Q1��n�PSY��d���+���4�R3�T,o% ;T���Q�'�I�#��ǭ,W��o,Ry>y,Eᒉȗp��H�}���j-�G*��|8VG@�aS0�:PuE�t22�П���_�	r��*�Vg����_��{$���E����0*��Rf�B�D��o��/����߃;f�:�։���������!�����@S���#�)Q�B*�@'9��P��h ��J��������u��̄��f�5NJ��W�bC�6(M�ɏQi��al_�1ذ3fL��1�a����m��o}�0W�~ze5��HH��)�H%�q�`ܞ�ﱤ���T�����c�0D����K΄):P�������FL rYO2��S/xm8u����8|� �9&ցF-�Ə��^�[����Ν��&������v�Ja�B>g�d��v��ug�����V(])�b��dBu$-E���#P��N1���O�A\�D�^�c$��~�z�ٞǹr|=?쵏y�e�Dy�.��~Z����؟���U��ZB-�!dn�]H���K��+���[O����av�'$P*H���5�L.��������"|���ɸ��KD��*�:��%�[-��SJZm%H��#׸7�<����[nB��:i��L�a�F�����w�Q�䁧a��BX!;[i�ZP'���/4u�)��،��k�	���҄kA��',x����"�v�X! ��>���KW#_�D+Ȫ�W\[���8o��I|�1���(��H'Rغu����q��.���%����,�@`*(���%�C�&���+d�F� ᐓ�`� �05R����m�JNXL	+��� �8N��<c|���Q�dƫ�7nF�n��³O�GCGaz�ޒ#I�
�$��n�]�q��F�{�L�K��q��/'
��p���V��9z`0��Nѕ٫m)p�Yl�T��y�s,:���#G���P��?%����2����1���+�� �@CCÙ��T���$i�XH�7wQJ&lh܊����������ۡ�d���P��ψ�5R9p��qD<%	���ao��.U8�\��(-���=F`�P,�f3HקE��}k!��5v�~vZ�z�d3�<�:�|������o��
e_"�N�	�~_q`%-8NP뒵����l����7�����4�Є�걲M��x[�R3�67�U���e�W]�'VB�e�(8E��������"��{������ϵ®1�4�m)��(l`^E��/��,�����
�s!2�#��	�詷����B@ 2��:L�w|$���V4��\x���	|�K_D��n�K��mx�չp2��͙gA_�u��\�AaF�H����:
V�z����Y�\�C\yZ��ϑu�� $�)#��W��(	M7�{�.WU����)���$'����B/"H�R,�U/
*�$��G)�B�"J�D5!	���S���ö́��������<O8	��g�:������B̆߻����֭���_�7,~�(��i'XV52�y�#RZa�zOY��o�z%������+�U+𾃠.ޗ�	VO�A��D� �� ���ŕ2�p�=ؐm��6��&��ۚU��
�nI��\U	��1��+ ���)|LX�!�b@d�֯��M��Z1s@fN�"A�L�n.�g���eq��>6Y��������A&��G�/��C#J0X�a��Ą02���}G��c��`$ #]�Ǎ׶i13F�׍�$ŮM��䰽1:ӈ��G ���V���Pü��`]7��xn_�^srv^ڏ%�Gڬfj��I-��	B����T�la���SF�an `G�Z#�B�ٚ�I�6�=X�	�͢T(��L�׋o�q<�=Û�sN�h��>���{�)���G0���O��i����֬�SML����
����Iu�(u��n��d���P2�	�	��/D#>'�l�Z�a�7*��9�����g�|	~��hniCU���)��Nu|�+U^}v�
l^���\~��o�J�=��A�������Nᓤ�'��_�2~z�����&�-��Z�!C���U۞U ��
�����|5�%�pEK(	1��i�h��n�?�ćq嗾��y��"���%�(����ٯ����(.�����Do"L2p�V��x>�9���2�FU��� ȿg�����8R��fA*+r��	E�@r�F5hAZLݯ,�M���.̾��>BBo�J���s�x��(�9�P|��फoF�9吒�C�>%#�Q4`�.x`�$�1�V����8�cU�QI4�"(����V������<��6al\�+N;�/ᤃ����#���DG��C��F��}�a�������
�-񘥣��t^W��	ܬ@�����C�A�.+F%�a˛�OY	כ��ω|y H��cCf��xn�[8���Ai���0	ӧM��
ؖO�i�x���U�+��yկZ_���;j��h)"� ��f*��$^���CSc�y�y�V�lO��y�5�G`0��V>��jJ�>��?<|�!�D��lJ��*F=!�:9��#�W4��u�X�t�)X�ĳ8m�}0}���S��Jk����d�E9w�B�n�2؝����@ojF��ȶ!U:E��{+"1lلM�;��K;�.@�+f :BS��,n�l)	k:���p�
�����~�7��;�ô)� ��vr�T-�����1�9��o~�)8�]u�0�غ?� &�F î�IU��rg�z��l��$QV�Lyg�K0�{`r��	���ba���k�����I0�9��G#ߐ&����)߀rX��W^B�w�ĩ���_��	,��&�#��S�4iʖ�-(����*[ʔ~pT�����B�|�3�c�MH���E��!D�����Y_A�#��=�Aɲќ�	Y���ue[�_���J�,R�)�؁+����Vo`{W�RZ���/�Z�D�� #���� �^_��6�"�b���³�_�F�E�>��6	" 2�MfrՇA���̔4����N��棛Pĝ"�J8����q��̣��������afu������&R"���p�<�����}#v���]��y=�����^�( �59*��lǚ��X�qS��N���n�W,QC��6o��p�ణZ��	퉓v���/�;OĤ�G�dE�<h+��!l��ٵ1����/இ�>���^\����Yx�.�8��k2G�a��-��5JB4��DM��SF�L��8�3m��y��2��F6�cƈQ8��]� �:�<et#Fxhȷ�T�:-b�T�pL/�����l�}޹����q�W��PB�)K�
�R[f��NS�(�
�Ê	�:*��cYg�R-^�)	L}Z�CO9��}�چ�O;//Y��Ρ(�дT�156(APb�H
�cv��U�t}��
�� 7U+�Γ���+�F�%k��[��]}=�>�4x ֐��[3��;�ڊ�'��Z+ �|Ê�������:�����}���_��]�a��I�1(Yx�� ,��6���|�I��=�fs潀�.�2>|��hlo�ŏ~%_C��zH���Z�O�>nQ�� ����Z�>��V
1n��k    IDAT������/c�)Si�D��鮍4��D!�F^fu��	��a>N?��8o�hn�ɽ�^����H�������V?�j�-�[2����5�s}���n|��L�:m<"��KEJ�h�cT+^�T���E�����W�Ơ�c�B	(�y%,Q:�k�r�1�B�/��Z	�:���7"�������kphX}���䁸�G��|�ԏc�����M�V#$!j-K<V��d�-}q����J��ob�+�W�ݬ����,d���tM�%��4��X���l��7�a���u�����a�&l�R�cu�S87"
�klQ.��7��I	�(e�5M'	4ۖ?�}%6m��ދ5K�b��1R����7�9�鎆��vV����@^����{����[�0cw��hik���7�EǗ�����Ȋ��M�hU�"���������d��"�"T���Ï��s0|�P4u��
ʊ����#H(� �:8��}�i�X)�ů�u@'N:���w 5uU��X۱5Z��(F��J�6�,��U\��"\W���Ѝg�|
�?�'����=�N�T`�c�y/��cDe�b;����X���f}���0a�x�z��AoR�3��g{V�2 �0_�גm��R�lH[\ذ$OU"<��Sx��?����G�r��|���ж��:n��տ���g�W���rì�J|Ͷ&���P�Z��J"@&FR�~(�u�P��W9zP ��
�6?��������F� �	7AV�Re�m�͚l����k�0Bjph�@�]|�B��T-��M"�I���9���|�+V�0�ZzJ�@Ά�XH�H_�:6j����![t�M(�q���e4����*46�hJ4HdCW�`UG����b���0B.�E��c����O� ۅ�bO0��$�����פ��6�% 	AĬ�5���K� �	x����@��/�@q��B�m��kl�#��8�G(����~� �d(s �Ţ�/	+�ςZ;�^���|B��MP!��@	|֡�	:�V	.	<��LC��,���� �}v��U�+�>���
���2#5��hg&�?5׳����"Myt�l���6L���o�&s@�=���X�R�r=7����q�)CY�DB�[:UxղL�XB�Ñ�(��pu��)�`�a()Y�tHoL��2]\4��n@���\֬��b/,��h������������r�%@G�sb�-`FoO-�c�Ф�a!2�j\�-I������YaH�T.�C����!zKU��R�v��IH����� ��><��J�U٘:�芘r�V�!���،�0�k45�B�π1S2�3l����"3�um��%91`�k"�RV�
�D�ms�d��9�D|g�3���T<�Xc�����3.RV��1N�<y��w���>��������V�}Ao�dy&Ěr��L�'Y��)���I��*
��m�gFՊ��J��xEب�����j��"K 1%�J��`:��x�V����ViYzr����Ԕ���G$��*�Eh��R�Mh���I���F�~I��6�k���U��%�����WASK3��>�B��2�T��F�`��A�	#QD�"X�0طX�	B-�lK��S27�l	J5Dޢf���TM
Re,U��a(椬�0`��
{e��#c*����K�N�E�D�µ�h�7,m�x� ���Ħa��(���aU��oZr�I��f��*]]|P�]� ֵ��(9��K�!=e��c[ڡu|7+^���
��
�� (���/����u��6^9��d�q�f���)� ����8�r�B�f�̟RՊ�h��ʫ�bBe
�2�ch!��TLm/�2���[��$?��>�o�I{��TR�H�R�x(bg�S$2w#(}��Q(�`)Q�ۜ�w���SsG�D����JPB��ʉG�Q�U�F۬���3���_g^�&���bY�K89T�H%dTm��V�co3T)�����&E�%H;�:/d����ɚ��G���u�3�6����g�!LVd^���F�+>~.4=E��'�{�2�5LS�&�*5����%��-�8��e���dÚ��j���H=z�Ԑ��.^����[�����{� Xߒ�+����V�`WW�v�M�͏�إ)�8�[U������j�2��� �y���,�W�ƚ������Z�<�ڟ��?��������uP59��M	��ͳ�F#א a%Š�v�	��X�d�Ib�e������B�Qh�&s��Oo{�ֺj[J:��x���-h�a2y9��z6B�H�"�.o��H�a�(n�6V" �鸚Mn��Ųuk�j�e���f��U[��S����ޠ�k�~�z��B�mokG���ј�J+���s.�$EDhpr�s�@�T�lX-҇����
h5 -�իW��c[.k���Z�ow jB�i!�����fy-�����0v�h�L�V��p�%�?� ��t�n��Ϯ���^�����^4����T��Mag]two�؛J_Q6jFz��8��S0z�q*%��?��ڙ5��T�̛U�Vm;֖�l�X"����jp�-YΧ���;w.���K�0u�D45f�W�r�A�rHu%Ó�a&ѐ�,h�&������	Ӧ༏��ɓ'���`U�EĨ�S�<g��ږ3@�۫آ�sj�'(:U�I����%o�ߺ�,��]&OD&��Kj�����D���d�� &���^A����w��	;�\S��ԣj4��
)�ـr7�	3o?��)ןmI(۳E�ǋ�=�?�����0q���זAw��+R�JOEy��(yHjη",��J%lش�6v���.��]�a��!��핖'_��]��T�[�:8ݼ�҂�y�|��?�Y��$xk�R�{����λ1~�D8�+�9�I��;�I���u��[Z�z�غx_A��C�A�kU<��x�~E�a�b%��،��z;F��5��֭��Tm��� aBOI�x�W�ÿ�,�H%!���yw�!�����~���>�'�z��e�(��J���#KX�� �4�6�����}X�r5�癧1q�Xt��Z��FY[�I�7E�%h��*��_A��-@��Fn��w��aH�������N��Q��АUC5#iο�� |�D�J^	�\����<�0	]_�b|�C��fe.��*�<Q@������=�Ȥ�df���m���10�XڍO~�lZ���D���i���h��'�L\����E/�֮�q�)'�>�ז�P*��	Li
/T$�D��V����$� #d]�#Ă�zh�z]�0`�`hÆ!ܴ�]x!����0j�D����T���g���� ��+W���
l��Z�QJ�6����%6Wն"+?�k��+bơ��?��\W�n�Z��檔��&W�9S�zJ���?�U!z,iBm�9e"�"$�;�0���>�4�.m��<~$L=��Z2��l射<+�B���h��=O���&���<�7V.CSG�2Sd��� /5��8�Qp6W�j�Q4�$��ϱ|1�&lж��Q��fh��ɧbz��c�;��+��`��D4��0�W:b>}OΝ�����~p�x}�&d�ҫ���U3V��DU����TlUM���[Y��W�N��E�x�¸�RX��Ow4܀KϹ O��!���O�H����$K�D�����P<�,V=�<Zښ�o\�y�yM��LF�B�:%L�~T7@�pҘk���Z[�s]��B�TSD\F*I��j{r�Vm�߶q�e_AۉG�G?�>>{ٷ0v��0��Z��w
3�z��wD�`��}6��U�+����FWW�vN�W��$��VE$oP"AF"���J ��<�0�}|Z� Q�v�fY�i
ն\մX�ؖ��;���}�����'�%��uu��w�=d"�ո�#�a��cR{+���3�b��7	Bvƀ�p�.x��{��q��B_Ά�ڈ�uP��0Sy�V��ˍ6�ꇄ�/�K"*��R�bj�t���I/	�mʠ��[��;,��e8e�=pԔ�a6`�)��CSh���<�b���sϿ�W�m��(��w�m������1֐a۔��OL� �)Y �D�����)�X]��,ͷ���т���e����p�.�p�>;ㄽ?��]� )��$����$�b�S/`ɟ���MM����Q��+����R�F%ʧA��d�N�fb���|}CĢS��8�vr!$�D4�d��2tm�&	�_��{N��]?��_���47u�4\�h���3��-?��J�m=�'�W`����V�w̚5��"aE��
C6Ze�E�d���S���k����kz���(99$���X�Tw�nhԼEU�����6l�1薥W`�b)˫�m�2�L�ҙ�������?�?�v;����ƘA�j�J�a��^|���q��@����?�Qk;ҖF�z�JȊ̈́�e�Y�Ѡ�D�X*%��S���*&��H'2'��O�?�	Y �!�>���fFP-Y�+>}&J/��#����fL�f&(<!�hi�7���׿ۅ�?|����Do.�y��Nl���y[��W�ܕ�WKuj&��9,IEd��5G�j�uUJ���\��n.<�0��٘2h �������Q ��u}�����e�\��������-`s&Z�Ȱ��Sq=�ڙd*S��jVf|mI~���5�qe��A. �0�����$��\�	�|�4�<�x�FŸ�;�q��5��Z��?K��'��;lo�_���h�
���;gϞ}��A3���E��\A����Zty���'�G�܎O~��0G^�l�@T�@"n$�j�&m��ș���������J�@?/V8j�(a�$�$��R0?��	�rfhç�#-{�:E�6A�����ѝ8��_c�������I��mO��� �+&\;#)��rGd��M����O"��*�����L��A�$�z7�_k� kT."� ��U��ܓ�S�aЯ���N+����᭸��xJ}��f�-�JN`HhR6�ZH�l�SN�*0�. U-�<��t�Kۖ��j�'���1��°9$�w�*\���p����KO<�ּ���gcI�^Z���^F�س�����1�y�/ZB�M�������#[���L��)�sA�Vu�t
��a��U-��h��i�}V�����ـ?-y_��\{�����?F�7k!kJ�^�I�R��UR}v�
lvuu�5k֬����A��J1�
�o��o�ǿ�3gⲟ����m��Y◜8$���BoI��T>��i������JV�ѩ΋6ϑ��E��L���K}$+��M|�{�^_+M��[�Pڄ���3����}�m�;�")P�m�)��hSV���4Z�q�'H��'��j�1�!��J�-�k�����e#���J^EH'�1已�ub����-眎G��9���m4�Y���$ �8~���V����u�XtG)R+�$֑O1�'[���
iO�ċԔ�E�A|�c_T�������	*�ַW�oڄ	�ŜZM��M+^å?��<��;
�Ǐ�_*¶�B\z饹�z�a�~�9�c=ܜ/������N�QR�xd󳡤,�D�<̺`��rn�y�F���&�[!E�_���#���,�d����8�o ى1Ӧcܤ]6W����;I����������;Z���믿���/�����B��){3�P��y�7�g�.ăs_Ě�<n���HZ"�8����EORDR��d6U#��Ԛ�Z7�oh�*.Gp�J�Х�!a{�-���4�Tz�@Oԋ������9g��B�׾������)R��h~��;�>s_|���v�CoERf��s�$����4A� �]�S�x���1	���k���O�m�e!d`�Ê0�&l�Fk)�8��\��+�렯^���p2�<�G�{�i�2~"�R(��%���Y�~�?�Q|��w�8M�P.3�Ɇ������PWf "	��L�I�1�8�AZ�Ԙ��!$�$��[5���>���#�p��G��'�;&&>3S'�E���C�Fv��[��uc�`���6�(�%�NN���#IG������3"H�����I�� 5:��u���mI�TQ≼��@�	�ىqk]�gb�3OEӈ1�<mZ5�W�ۭb'����X��������+��V`�@����Y�f���@P��W��14AP%���?g�B�e�[�S��mO�����<MqN���y�ϥ��b5Gf(�JD]���R=-c)I��k�{��S�$���4��*I�$���=�.^�k/8/�p���7��т������^��<���{��nA��p6�p	�6��bTBO􁖞S�&i�����G�y�P���T�L�4�g3T�H�U�7C��u�1�ۧ�t�5��V/ŵ�� �7v�2	���?��5��7��=N=������� ���s��r� ��4��Z�T�I��d-�����\>�2]a�rH)���g�%-ª�hM桓KQ|Ћc��{�:�9�L�E� �(쁟\6׌���q7��̀z5�e%(���C���CA�Q&�E%�P����TD/3mU%v�����4�*�8�ѐsQ��D�j��B�&�o>��y<v9�8�;G`��o&�ԈL���?k��Ap��m��W���ւ�/f͚u��AiYJS�_Mo��[�k`μy��%x�/��g�E��!sNE�c:�3$1C�Ch��44�\ijD+}0C��N�5�x;	!�w��`eoKz{Q��c�E��H�4,Ĭ��FRFy�b��3���7܌k.��Ç��؍\����q�4=�8��h�2����(fѦc�kR�FB��2���U0�_;&��	m�m2�z����d�z ���ˣP� I���c�I�Z�d���>�������C�.^���S��,�5�W�_�s��uL��9������}�g3�H#"2O���P����YA��
�b��41c�$�X#-���t�r���C����5)	Jը���ڃ<�K�'��u�=�`ό���`�]&����Jb�^Sp�W�k�nا�?�,݆R1 �ag�,��i-�/�Cw����x�Ћ\G���F��qP*�a��Ux�O�cӲhji�Kp,�J+<	M݅:x+����ñ��φ�9;O�.m���|R�ൃBu��w��՟T_�w�[��]wݽ�g�>n{�����$U�)_J>��G���>�'���b�?1Zs;T���sGC����H�٨��9N�>���D�\�F��"���T-~lc�_E�W��~X�#�5X��\���Ȋ��b�B��+����N�3�܂�/�2���&���e�y��h��>���A�),C�.'��R#尯����ʵS�8���`lk;2B,�f��Ҭ�?�X�_<�g��~��2V^Z��?! ��ӄ��P���Y��~�W�㰃�Ì�Sj��^�f-Οu%��y�x�h�%n1&[��R�.�{��I?UJ28�,�x��7S;;�	�ϔ�fe� W�����w�p��᳽h��e6!ٯq,���2�ΠЍ�����V��G��Sw�5�5�ӹ����[�ĵ�w����BM�F�2S�>er/��Dp�RV�"�O,]���*:v�	�dRq`��^��� g��&k��$�r��h	c4��5*#6�oc�݌������=�8�a�4m���Ζ�DGU���?�z%�������+��V`�@���뗳f�:v{��S�}Y�	����>��jy��g���70/��'��l���e�e�E�g��JZ�B����c�F� I=��O����f2��5���KV��E����(��&#��Ķ! H_P�`�r5�8�d<}�-��ҋ1��S�^Sॗ��_�MS��~�0��#�Fl�*�2U�*��u�kc�5ڸ�&v���nɒ�x�U��F���ڡ5g��K�񛹯�q�p6VD�[�f���?��ԄȒ�]��q�W�����������a�z|z֕����q��w�y�(ĉ	[��1�o��uW��+p$*A��p��8l�`4&1^]�Z�o&�4��wJ    IDAT;��Օ �/^��^[�\���G��%�&��c�pE���AQ_m{���A!�8({e��t\��ٸv���w� ��#		������18�"kX(��|=.��4�B/���y/����H7�8l ����_['����{�it�6mS\h�ڈM��3@�c]�`�QGc�3�@f�L���۠�����^���믿���/���d�.�|ؖ����y�
���4����ۅJq
��0:��S��"�;��(^Im�p�E;�(A��G���I�)�$��z5�<�d<{�-�����S��j��+���3�E���R<��B�knF�(|p��8xd?X����ޅ�m02F��i+&�6��g.�S�:_����g��K[�6+C~%@�1�DrA?�0���Ǟy��[��"TV��Y��FE�|��CY����f9�@4�l���d.�6� %��bi�Ԍ�[���=��~=>v�`A:,��[��/�ƴ�\��[%���Nu�m�v'ۮ	'O��ɶmkrM�lL�m���<_�������ڏ���Z���<�|�L<�k!�!�q|P���8īH����)T�S�g*���>�j@���� t����l����?�+���Zd+��~��s�Y�����aV��A�8�ukl�qh��D�t���1���ã^�|~���W\?^��N�I����҂����+F稧?�������}ǥ��������ma��'��*_^�H�KK{4�lq�v�ߔ>�W�xI|ql�&�ԧ �?M��n���0槄�q�\�8$�(e��h�)���hjO��85Ά'����|q!ï���:�P��탰a�c(V&t��8U$P<wƎoO�b���&ӭ_�����W(x�����t;U�����C�З��"�a.��I��u��(Ҝ{�>w�I0<� Z�!
2Bb@q9v3W�	�>��""��,�U�x�~Ո�v����ٰi���lq�G���s��`[���|<3����4�3�#�(+(K�'���6���Mzuz��s��w�ڣo�y���.����m�"<*�щd=�}���:����(+!�?/U�ȸ�
J�H8������dw��@�9��W�,�j�o�(Ue)'��,�L���,k��4�e�r��O�n�MP�H L��X(�@)��N7��13*�R�������_�����H%�f����G��]��v5����H����",m� �0-+��тi]�H���vG<������ie!vz�Qxo7x��r�pd�`��4�-��kssQ]+p���z�ʳV�xgVx�eNccg��n&�;�Q3B+<�
tΕ��P�1Y&��ѷ����_��1�|C�T.�'�h��6K�0=�y�Fy��C�'����rc���n��w�������%P��w�A��R��g�-��Z��e_�?�r���D6�^|m�譽;GYVh<5�����]�9-���������'�����:?������JNB�*$��-XЕ��B LRx�i ����FEr����6�{X�����z�Uі{��+-#�Ə�hČ��b��������E	�X�eRR�;�K �L���c ~d����$����){c"f�$Yr�N�09�9�I�����]���Ё�P�RB�^�X�Cs�1I �Ӯ���Q�d�ȗTi�.B���O[q.�q�B�ﲕr��/|������=��yjY�<j�&e&'s���i��Z���� c^���x�_!�)<O�������u�^v}��I�G���jHq�0��e�R�:��oy�9��|k��Q[_o<�'�Ώ���@����H�)'U�/.2:��H({�Dv�',�Ts��?snѽ��а-6���7q�Rwpkۑ��$v����;�r�:I�'���WT&��e�z���:|l�P�����G篛=(�28 �P���f��{���hVRL� �5e$�����)���h[͜��$��C�DI�V������⻝�E	r�������~6�Y%u?����1	��(�(I�`� o� �J��֣�9��9�3�7�?�?�z�������p�������.b�f�ɾݞKV?�}J����Ο!k��\��w��!������^|d��	ڃ�I� r#;Ƞ��Qx��e��A~ŋ-h�q�,�[,!�9�!�p��¸���xF�������EO^2O��7X��W.׸���µ$�2�x��zN�.��`60�1K(�Ym��
�*7x7��57Al�&��]/~�~�d7��i)!�Cem�6O*G��$����iKPA�<�,8$+R�6�u��*0��/��0��{8����q��X�+�9k��[�J ;ŷ$��i��L�`�>��ۋ�F ��~�z�w5�E��*�z��٣��5���
�MA�%pÄnJ��n��̎���G��}d�>�~7����������X�0s�	R~��S��UJSd���˭
�J�k޳XQ�PQL�'п�z���]G�_� �c�N�H�^���v_x�H��%|�Fܫ�*�������W�vz��GzN��f� !k�{x"�W`V};ĥ�?�+�#]�.�w;�̄��1jЂN+�]l���[!	�����Ŏ��h��¢5�Tk�2:�x��h!w�*��J���|7�<>�3G�j�}bX��>�(\E�������	J4F�#���ש�c��(I��D��DA�������ͪ�?<C2�\�E�GR�ȝ�{9sj�R���FR"5c��(�~<�J��hH��酄��G~����0 ��%yZ���B�pz�oŶ���@�3%���	��3���o�z�')lv�a�b�[���'��f��� sa�){�����F�uo���q>���z���*����(�~���w��2���E�<�k3�
��G��B��LT�gC�fk'��$���Ƣ(Hd�����k,
S��Y�� � �DA4}����&�U�t_��]���DW�d���%c���v���Si�Q��P�^)�4Ovh��uIꘄ�;�H�N8
/�:^�3׍f�|��b���}�U����|ԀT-����#�I
^Z2���8���{�8�(*�r��6nO�6���v�0�3�R�@37;��*����b�#@�J��Q�	��V��&�/��%� B�tڧ�x}���N�lX_q'j_V<xGz�@4��Z!���.�D�vY9���ZD���ce��BL'�<1���xҬZ���_Pb�B�4Ǌ�&-,2!� ��	�x�����يmyC;"����lzB�L\y=��,<�V#ƛbO S�΃	�#�xΛ���c��g��)�0��X���hǳ�42T;%Ԋ_ �O	kh8-,GW�˟I�8"#aw3��1�r1�}�����B�W;�n�l��n�/����8o@�9�>�*/�.��O��G5�沔Dw�б�� 2��/�Ɵ3�~/�f]��S���Ey6�P�8E
""Hz����
>l��'9��v^������z��S�n��my#)�:��F��y����tw#!{�(vV���.ߟjN�]n^JN���YߟT�KM6ȍZ����Lئ�KEc�3t��3�!{�F���+zxi�{��vGXY���X梹̅��p��Z��t�1� PK�*��4-Y�����a@�i����!y7s�p��6�4�Iz)=�IZ����%��9�T�E�հ8�Hd�{���E����ޜ�Ј�ޅ��~�O�^u��
�%*����>m�g� �үl����G�ob�d�9�Պ���؁�Y�A�W8��@�u1�e�T�h�d�F*�U�7��~> P�$�)��Odhx�t�),c>;���K��1�����^a)������2����g����|'��We�?��:M���N ���6���2��.K�Y��0ėͼ�FD!�ӑ$xS���Hy��"�l@=���
��<i��\S�0'�"�è�#���XPEV��F;`o���Q���}%0b~��m��� �RX����"�"˒�L���X$��k>3��(QOih�҈��	vF��W��;��<m�������_{���v_O�nގ�����]�J�0|PH=��>OM/���ْ��~}`3^���ˑ���>��e�+T��W� ;�1j�I*q�M�I�O�/�{�W[cM2:��'j�c�a���Ӥש�����Cr�f	3ęPg�ߌ���m�Rg�	-�5u���:J׌��o�Q$�P�������߲k�80H4�����"E�aNAQ��=��)
�&�L��{S�_����7¢N�"+��vjVtR%�t�L��%t�\H#�r�sf�L�D��4`XMw`������<�c��׉��Fq1�e3�φy�HyT��{e�D������!��h)|{@w��T�?P��]��;����영
�e�N�j���R. ���(c�+ ���9��)+���M׶H�9f�UC�ܴ)�O)�������əK���k���{��Z�Qd�Һ4�,M�]&�e�f�v�A�^�;~蒲9'��xԸ�9/Ӏ�j-�{�jo�ѯ�n��T`�}W�{�J�I�GA� 
�!� b[ےő����Ղ�
6���Ea嫁�0��;����S��f����r�}�#��24��}f'�]�P"Tԍ�Z�V�8;�:{��8~ӻ[L��}���t!a�2��]��>���/gR��,rHX������^��'�F���bg3��m}�N�Y|U�����fo�g#��?��*z��^b����b���)<2(})����ӻc�i&Fv���y0x�����=�&�ë��nr֑��qjF�X���@E�I����V$�I��%�z�a��/� �w�JiY���P�@yd�y�n�qn�n�et���{M��	DǷ:��a��{��BP5. Cm�f��a��n�&e�L�0S�2��^9L�^�w�U�����zY7�e>kR���zBC�cޞ'����,O+P����
e�2s_��e�������l�gX�=��˵C�:[���_�I�� �l3�
qu�Aeྐྵ/X���lq�(�w���U6W����=hN�� ��Y�G�%7�۝���}l�{��ʑS�|��U��y!8�/�I[F9\.e�ހ2��2�y�#��;#�Y���X{�Au�7���}Zk5�e���5Ʊ]�>�4D�l��`R���:��2��|ʰJ��+�z��5C�{�����J��0"qpM@!*wܣ3t3!���	:]g�O�����?���w���WB r�9Kv��`x ���H��������>��7<J�ΙݻMY��r6I$}��X����3�72�����B5�T�M{C���Ԥ�A!�_�3�Ѯ��Ӑ���� �qnT��;���Y����2����_��O_�a��_�ò���o3X;q�Qd�!����[�����\�JL�a�g-���ޯ�E�7Q�'K��9�6Y�<�1b4�`z�3s�j��oyʹAC���2����vE��_-�>�:��6������ο/�	�d�����Ճ�"MVY^c�r)誇����ܖ�MpL�a�RE�Q����Vf�Y?�i��1_,�B��fV��Y���2:م�K:��u�V�g�I�>m��?A�9���[N��v�e?�.Df̮�pm�@�J���D��`ܗ[g{���}�f�?(Bd�$�Oj=g�e0N�����O�N���Pvc<�Ճ��vp�V%eF�F��O3�|;4���BO���1p�4?�FZ��@7]+�u������|��έg?�(�z��ل?Q31� ����u����3g��o�d�,�9K���z%�����L��1�3�x����X�n���p6�k��~���'qv�i���ՋQͰA��˴N ;��q�5�x��v��[�2�lNk��y�r�8!������ś�L��)U���N=��%c-(Xggu}q'�D�C
��u����`��:�Q�2��Ig�g�%��0X��JCV2��[����y�A��U��;_�2�=21��j�O��'�K��ڷ�:3 �SD/O"�H���R�I�ℸǉD+�y30���^F�p���J���o���<����v�qz�OÓ$���Rvd`���	[r��K�+���(˕{�͘Qr~a�4q������ሢ�-�����Г�M͈��p�����Ѧن�tٰ[+͐��ݴ9V��L�j4�^!�e}�ϕt��
�����,SL��I''�g�g��D]��oZ��E�y �nK7�A�@@���$C�\EX���t�i�\gr�.��O�(�x`yh�o����y�r;�}NB	�!��;�OC�C�j�͊�ǌ��4��BC�V����P��J��i�Q�tA 33��#�I�{�[pq�!�7�+�D�r�:�o�u9a�b������?7d��_�s��p�!��ڤ����[�oo�m۳�K�+(́M�� f�֠��/��U�~9^ft�Dhj,�~-�D'�erZ��ֈr1,�H�{���)�@<�}�7%�����k(���#��g&�1�<}3���T�^1�
���~�V=f�9�-6�����Y&Hw��7tP16��X��X�gϦo���<�:��hJ���@�u4Lԍ��`ȩ�1�5uv�-�zi?ϊ]A,�"W^��U�H�5��7�k����x�t�?������!!�Hk���Z�7�+����&@�	�4�������C
�υ�	���a0I�88-�7JV#�F5���&�vt��a�_s��3��8q3��OÐ�"�WZ�K�;�y?��ɪ�w�6w�t��zE��LpAh��� -V�����ef���7���7Q�S����01D�IZsXy7�U86��t6��4����ljU�`Ĳ�4�^�-�×��E��F�9m3�6ʩ1u>���q��aZ�a��`۞[���g��g#�]��ǝ�����>G�=2k�lwrH�9�	X��d�<���&�y�ђ2�q&,v������4���e]�`���%z�xtH�)1fd��}�!�!�8ި[]�G�t�H�>�0�{.�r3Z8dگ��D�)!���3�f$X]�aH�D4:l����-/�"��}�O��(6N��t13�l�o�j��jX��c����<��L)��x�}��B�+l��[��|��ћ�Gb{��5 �7R�m�Wo�����#��C-�r�� �	�ꌭ�L�QKv�ʪ��l�-�V����T�,o��4��B!�ȥ�,^���s�����a�<�;G��1���E��5��w�/�3���{��ʿ��T���o���h� ������uL@�~$�$�p)�6!ޜ��f���~�<��������\J����?5ZD!exf�$��Yge�V��{Б���|2�6�����K?(�=���ĹV	��3ï����Χ�Z-��~~��*6�g��6j��:����T>Xy�q�+dƦ�
j�����Iv0oĉ��QE�Ͱ��a�Q5�WG�0Ħ} �3iS��`��}{޸R�8��C7�=�H��M��\h�F}��eXTn@Oa���P1�D�����y �G�fX���#�#_ϼ�e�fs�Q�R;r6���7�/��+��E�"N�@l���] �.�ѩ������ �_9�dW�"��yÂ����J~�>�w^y�����5jyKV[%�ɩh�0-�$ءi���o�`�)����'�\c]�&�������0��1C�<���&�]]�S<�9v<���o(�L���'�|�X@�s�4L�<k�s�f�߷������7^���h�n�p"g�p~0�F��t�&C��FC6��٧��R�M��M��ɭ�����5��R���Qk�����;^��u�W|iRg����l$�H�e`����i��R�1�c-�]ȥ��gy�^�T��U��������?�7�g*HB-:_�MUA�Ը�i;aӹ���)���q6cb��]#�L�� �	�!�SD�n�����'�,գ��w!Wr�r���v�ݓ�2K`Dv-&�]���C􁼻07� �ԆI,#�wm��.�,��:��/����<~�J�Ǆ�+��@M(s8��ߨ�(V���Rs�G�e�1|1����hP�9=����%9���Y�"L���մD���2� �b��_"�˸��1s�;�Ҝ�o�Zo6��bCQ�"�3)��;���Х"�
=�|-6<���;�r��L[Z�1�����4�/���C�D���n�:귞Y�Ő���oe���������vG"7WF�g��=��nۏ�ЫGm��'�Q9���*��?����;�Ka����~�7_�k��5�H�KU�ƒd�	d@3��(!�����E�����3�O�� ��djf�n�r#o��R��o5: ����;��n���V�I��cr��T������=��i�|�Ha�M�P�#��}c���e	��p�	�R	{�so~C��F2�[�2�/n�eYpX`#�O��������8�y���\����7�]EE�����"OKEE�*M���~��g!��C�P�� �������t���VpNr��@4��z�~��~���ģ���)�H�ow�r,�y��EI�Pِ�3���ͨf�:o/�����ER����<U��&A��m�2ώ(Ӭ�h=F��o�7� +V���!��l ^lc�7
�ۗa5C��~q�'u��h'��L�b�ՠyU2C�T"����l.6"�W��e�^�e�(ea�{�/�c!�vm�e0>7[>�#�3��$oO��kTn�^�7+$,�����ょ*���$C&����s-7BJ��̌*蠷��f�}��F�d.�i�l^�%n��gg8���w������������J���Or4�ں��׷u�qC�@�-�\�T���v�R6ϡI�OOf-(x��Z��6�@���l�C�ϛEbO�W��d�]��P�� �y����݋X�j�&Zm�n���o�S4�N���%�4�Q_����e��1�n���ub��$��Y^�0��%n��^�B.���}�o\��N�7�/*�u���cg9b�� ��e��VkBWr�����|D�9-�+��P�b�Ǚ�ȿ� 	Cp�xY�tA�����^g��ź۴�31�(V�c1��h1T�4oix��ƿw�侹b3x�e�� ��G�UY�����#�-�m�E[
=0C+wĝ�8Ȏ��ks�i3���QE�}��OM_��B�oB���a���HB��p��X��Ҥ�X$�j�y��k�0���x���u
�Td�zQ�])%��Z���;��[H�C�n�
���,�V�H�'�{��(��7������9M�t��ޘ��i����U�P|��C�����F�<n֥��K��/�#.�[&��Zs0\PY۝º�y>=̱���{��(�~��;��ͪ����}R�U&<�O>��K�CHzӚ���n�H�ͦ�4IP���wY�*)�L����/��(+�,=�ٻxv�A2$�T�.?$i5 ��:�ȸ����ig�dח�\C� oӃ��#���ĳ0�C�hBQ�Kx�K�9��%��5F ��p(u���`͝�T܂��雁:b�w�����IK��vTZ⪗�N-c���������ٳQ��}\��ڛ$lk!�*�ħh��+!�,M��%�Z�կW�Giu��
yD�vWM�GT�c}��9��'[$_�NH$>)IB�4H���C� Z���$�E|�j�=a�K;��Hc> ������v��:D揚y߷�0l������pP�KR_ �ÁWy�VyE8`ЀtL��C������g�����-�G�O߷o�j�}к�w�):;d��~�;�.=��)�(8@�hX��S�"1�$@�X��\�Q�I׆+�J�N#����ٟ�\�X��T	`f�LWm�����'�L��듶��\��9"0�\�6<Yuċ2^�a%g���,��p�V��]b/<�>��SZ��d7Yר��t��EQ�ۖ��ԝ+�m9Y� Z7G����qE-�/����)B���8O_\J��T���Ց^ebG�x��J�H
H� 	fAy��:>��/�����*B�۵��c��PI�����Z� �0�{������-���WQ2)Y�_r��k]�pO�ԚAo�DX��]E�l�#(!�=BԦb}Ƈ�����e��h��4=~��~^S�����K!�v���^�IH�s �S��r@&���ƥ�ΜU>s�Uq1���ԉ�WDJ��(�����|��eNu�f�3��>:��g���1��߃ݼ*�<�q�0A�8@��vL�= �A�	
F�"�
����;2¨cz��3T��"I��X H����>6��L�H�*�V��ͥ�/�����{���l˚���G/�bϕ>��2)6;���_fh�\).%KK���l�&CU�Ӥm.S�	 ���V�A{B�T(�t[��t�*߭�O����m��v��,UUld(�=��6�x��-�Eΐ�^tr$�h��0"�f�����ے���+��8��򶪽d �JI��r�j��5��-����d�Q<�n8��=��*6��]��Q@�H��v�U��E!E�Bd���=�f�y��j�֓B�/�0��q�4��/�ٞw�[p��i����=��W��_���Ɲ�a�<9K���^����鰈�^�$>y�����U�/��� �>0ͮ��R�+Fzy}������]�m�Gלt}��N��D���u��t���*����M��ԫ���$
!����H�D����m}�	�g��,��΍��6���kj��U�j���P�R�Z/���P��ٲ�r��ڲv� �	5K�M�
=8�!I��+���HūN��dI�n��<W���v�����+*�����P��󻘔��V���^�t�Iy)�1>��F�st��[���^��?S���dc��}v�������e�#jP�F�À��!���p3a���6[/d(y�Dh���`hTR��"$�G�.7�_��N,�V�~}������	����y_Q��$Y�˷+��2d�e-�f��ϗ�{�˕{W���F�F-���GB����R�U�UԦ~��i��d� FF^a���;�^�\��Xci�ym��_�_���{���P�R�6M����!�L�16�CY���`>&�g�29��*5ʧ�2�N����h ����4-�}P`vė��
�rj���A<7��x�N�?F�O�P�k���Ak��3\��#Q�7����-��-�Eq3�d�1.͠[�YLU9I��R�٠��ϰу2�L���|,y�D����F��d��r�I>��U�;[�Ɨ`z�6@\?�E��6�6v?����kXd��gB���m�7�7�h�8ນ7Q��R��N{!� !l-�F�
�4j�d�Ka�^N\�T�ɩ��s�S���� S�G@"�(V_K����b:��Ǒ~�	z�2�((GE�B_(U;.�E�#8�9$6r��c�x/J�x=v�j5و�S"���֥y�hն��Ѧ��c��d�Cyi���t�ΤԠ%��c�uxc�]��Q`p3�L���T��x
='*p<m�1+���DK'#�yx�W�.�Dzޮ�`�d���I��b���Z��R��t��qr��(�4�=��T��\�q[Q�R��z*J0��`����H��R������lO�L���ֿ�r4�$OPZ%�Q'�oF ��*Q�B��K������5�/�Z�v���d3x�,I��j�c_e[R��%1�P��J²�C�]����c�&�M$5��F=�`˪�A 8�*��H2C��6�W�D��?h8���p׹���QXB�`[��5Z)��)0�!k�L�ל���c��:P^���e��sC5abcڶ�VQ�p�bBSL�]J��ԣt�)`��Ш��L�8uι���^��3X��7Q��a�s_?l�}?�8Q�1��w>�]^:'o���WS9��J�nK}P 3
�@�������uqWr A��6`}�tH&j�u�f���U֩yz3B��w��=��>$��;���E�47}��m�]b�d����X�]�� �Nٷ4��Ǉsu��qm�Q�� �犊
4DNo�FsW�	!���"n��<d-)��-�	&v�OI,��ְ*M��aK�2z�8���Q�b;b6t`����z����0{Ww��<5Î�ȯ����e,��f#�Q��;,�w��4���g�������@��aH�D�<��lnR������.OS�ҳT���%'Lk��>�k즴�j���Ԩ�c\)��!�
��a���n������W�~���.E mM�vL�_���[�n2��U%�GD�+`����a��@���O)�	���]|�*T5�������8�͒�J�^؉B2s����� �mr�����h�nv6�C�z�,�j%}t�B `jj�v���_����̐D
�$Na���?��S��K��7�')�kR�`O2�������+̎�9�VzW�#�����o�����R\=�$����5���{ H�c�5�{��7�6�(�ف@C�i'{
C��RT|!5Y�֘{�J��1N%B��}� ��A�s5Zkv��l�J�U�4�����f���/��ͮ
ս���HD:>�fZ�7Dp�I�*q�v]gQ_�k�K���"J��oI<{�fҥ]��) ��`�q�R���S�������j����ȶ��6?��n�Bݛ�ҝИ��oXe=/�g�z]c���l���Cl��޾J��t��K���M_6�>_P��A��j��X<lv ��m������t��,�l����"K��B�#5�Mp9�^�*����-p�Ԋ+��$��c���r�L�Jj�r�H��æ��4UY��m��\�_h� q
:�b����p�pW63��f���hM��8V-����&���+�	�#8���S�};_Y��U%*��R�cy1�R��A�0��8q8GK�v�$��T�i�Q��R���$l�I?yK�5�Gz2�������KɹȌ3�"}�<�����j���7Df�	P�q.�p_3n��Թy^��!ea�52��W�!���y3�H��'L���A�O[����h��#�=u�~��+�6��tN���Q3z�<!��PZrCݺBUv0@�tVP:h�4�+�A|�m��RQ��A�mLGk��������2��3�N�C�i�|*@4y�aJ��s�FG!"���N����$%^r�GQ�=]�Z<(~z"m�R&I��<�`��0G���-�l�k!�?|ބ�p�gP�wN"މ�;[[+�'
<�� �[�� �@�sR���D�eʮרވ3u\6�w�HHǤz���p_�s���ؑp?��%�(��3��I�A^Zۭ�F_�Z2��-&pM�z�z)_���tc琹�{A*`�����i��D�_��".���ۮ�&�&#�eG2i
�G�5ń�����V�����~Rg��K[�Lp�;���U;��� .�3�?��f��4f#d�!�Rub�l=�=P]�	H���LE�б���vw؆l�Yr;wj�2;M<�iu?v#m1|	l�)jo�������w0rA
,�rntI�v�Q)��z٭��i�����J�����ȐJ�z�Sp��!\�k$h��)�b����;~�rqH�Z�+��?��+��F�Q����@X.Y _���G�+�$mB�|�%�y8Th��_p�]x]�ޛV#�o����^"���#����E{��������RV6k�+�އ$�������P�x3����n�BK�ODbW	�jy�3?�J�1V�b}�gz6�!����������SЎT,�r�R�����W~W	�b`t�lN�$��=������Q�`�,��%��K���X���r��2�J /�	K\��~��]�\Q�E�\�� N�O7�z�ݜx�Ɔ�8��iTF>K���ӌ0�v�� �U3���Cs�a��i�KB���;$������)�t�.�U�9wC��F=�H�/Tԅ5{%ρ6�^��x��tWf .�$�9ڏ���L�u��n���!'̣�+te����@Sm�%)�2��Z� 6��e�^�����	�i�KnD��(�����c��g�6����L�O���s�ߓ�����^ +� 1:a���F�hM�fv�����n+����f�n�֏�&B���?�;���iŹw�%Gʫ>���o_"m�/�W����PbSu���Wd��ѭ�K牐�n�	_���Hl��Z�DG�p��@tx��&Ǡ��.F��mS�9l��F��x��zpS�6g��o#�-PI�1=�hU�%�Ac[j�m��41��%�S��R"]�b��xc$E�����:Y��xZp	���_[��P�B����j5�����_=6=&^Y8H}g�ߓ�hX��;Đ�I2�K�p���J�I�]:�9��5a\�w;�/](�W�8��MX�Y�}���s��Kt$T��+"��P�}h"i�z��}\����1��ެ�]I����M�~u��L��3J#"m�Vb���PY���2 ��n���et��%/��C�D*�	��#�4�{�zm��mW@��RJo��]�{J����D{8??W���?^�yo��������f
��u�5aPu&b+�{q0cj�7��*LL�ʛ�q[;�E]��.�����n�%���~��% �O>�vۧt�B�I�,��iRsJ�E���Q��p1���wm�/�|��@� �� A�i]��@�MS�o���3���� �s���1_$@sD9�+g˱�1i2hZ�x�*�j�*��HK\�P��mM�jM�YZ����HCh������-%qi�5E�ve�"�YI�$\w��1
"�)Ѭ�(3��6��_�(�}taܩ��N�Fn�R�j/?\��L�k��4�i`�p&K5�L"�&��搎-�	��I,>m��3�j���;y�uq��XeA�5_��҉��n{c!��	�'~[�/#�+UY|f����3�c���X� Iw�5�}2����sy8�_�dD8q���\�����N�A�=&X%�/�R��v5���c�n�~�&���ȿ6R��D��@D칕J�9�� >T��#]g�����V��7���{B��EA�;�'���[����`d�}����"?�rlܚT��p8/E�=�w�k�|tE���̂^38�n�*>ͮK-<�� �M�q��r��-Y�/�O�d�4��Q6.hD�>��<�e�����QQW��噜���C,ؼ�R����:_7t�l���ܫt���HIӠ"��*m�КF8�ݒJ_�Un��2Lv�"\�����y�Bx9�ӣ��Y%��b��lY,�}�[������e�7��A�S����3j��E_�[�͹���'Ib�.1P�6k�aW�ՃG�e��u�tĬg߳�����B���y�2�k��]���`����,^��h�N�8��Am�S�>\q
?e�ЊL�f��|�ۀ��r63�i� Dy&YM�a�ԅj��}��1��$Pِ1�Xss%����pl��Ml�fn�'���!cxNB��'i<���g�H'������3TPh���R���!�
C��; Ή��Wjc����2���Bc���� �G�i���+~��/+'���ݯ��0�41�B�XI���M�P�[X�>J�͘�0UzOl뤴�_I�u�F����*�i��X�����H�Wc��z'�����^�pi�`�/�]_,�ER汶�_�GH
;j/�W2��VIP+"��ԷV�r4��(E����v&�Q;mQ0����@=�ӆܰ�]D�m�')�c�t��H�1T;���r�מ��{���b�r}���V-;zG��d�������r�M�P>Ri�]+1}�$R��kǚя��y�`r�X�_��F����
]y���0�6j{3r��©?�\�Hz}!�^+M5��_/U��U�xr=�o�J��5�˄i0����zA�ؽ�v�K��v��&��&���ny�3���k��~2����W#ׇr;�� {�n��v�z��p<���O
�ƕ���M��O�h�;��XtPJ|v:l��'v��KE!�����zٵ�Jr�)����>��V�f�25�ӷ�QE�9C��c�n�hC�Lc���u^A�`�=��:�I ���zl�s_��^�}O�!2�̏$W��X*w�,��R�!��NH��O�F1�J��n�K�K��k5o�� Z�C4��VAKV)!c�M�W���-�n��CM0W�˷���*NX���$n����n-�vB�u+��r�"B|�"���C	;/牪[�M���a�A$�S
J�S��` +�%����=@��(�R�XJ��eON�.�/���?f] �U��0+�����
����u��l���	���G}�#N��c����k�@�e&8�,�w�-TD���6�,�\��C#��t�!���IJ.�-M�VX��6]6T�����X9��SѮJ����l�)��	�L�,��2�T!�����������}�a�_��^\  �X�����(o�ҧ�D�����&��u��C���M/b�C1X����&�7�9K���Qێ����i̺��^Qsx�U
>h�@|_
l�!Ör��a�J�@�FQ�����w�;���.���R��uS�����@�M�ՙ���c⛢+a�h'�N���Ķm۶m۶�LlM��mLl���u�Z���{UW�ڻ{WS��/]��]T�Z�$1$�=�]J@�K�L�����S�l��x�E)���a�#/D	F�ƞvY��t'c�E�c!J,�U;�f�u���x_ur:���}�9��F9�_��>[k��5�� <M�tR���f���|�jM�܊�5p>�+���톨�E9�K���K4٢��'����u3q��7�����4qeU'��B"�(����ɛ�"�r��ݓ^]:aɝm#�]M�aK���)��[@�J��O+���X+�K��E�G� ���@n���FWX3E����x��o�~�L����ϋ�CQ�>��zl�K�T
'	�_����W�����P�5 ��z����9	)���j�.��jS*@�1��eᶅ�GF~��B�%���t�\jLT��Fo�e�=z�"?D�� _*����X�Ip�k��\(-=�J�ۉ���%��%l&�_z���hZ�at�}r�Yn�����MP78��H�?6�B5ܸRZKz�L�Hali�����a4P��ڂ� ���BĹO|��)�7���I����ȸ8״�*P��cW�
ʮ��9^�_����L&߫3��ehc
ި������� ����^�%�W@�I�[b*'�AI#K'�������>޵%�!�uH�Z)(�ZaU	�Ɗ/�\z���)$eC������L	O'f���)J�= ~z��ل��'dgH��"�e�S�;���-�$nAD��u4�֑���et1u����Ⱥ�� �c�5����cCV��WЯ ��X�9�`9���z��g/��_{E�����8H&,������	�E1.��5���	�hy��y���}`���%�R+)X4W�N!2�PI0A�o^��5�����o��b��ንL�7������3p�h!�;A5-
�I�n��r���.�0c���ώ��������~L�b�<��%;R�7h,�9)8��\�ö��B-�z?�8�a���Po�B���U�D���E0�qN�:���񈦰�
�#F��Lip�U�g�D;�x�UW}9ְ�E&#{ew;�x�V+ȑ"?l����F��P�f@�8A�Zy��͕�$�DiBF+5�R"��/�\���t*�5	�r��D���.yu��F�2�@6C�`1D�[��Z�ؒT��F�Z@�KKJ Hx�4�y����87�-�HC�ph�Ȑ-N�40�x���x�%L���TP�f!ݣ��}�Eق6�����p�O�$��<��}�w���|�g�B��|[`��<��0A#�Ŗx�T�=��a3�8���</VQ����_$Q2����;X���J�2��sq,���Y狞O�����̰����^f�L�Q��1zl�A?�
 ��v��5-F�۟������\��}��w��������@��|0�R��T��;%4Kt���"dE0�ǿ�Ո��}�9�����dC�������R7�򟐪���I�j^�{�����,�R�V�;�E��ؽO��ïO�b��3Y�J�J�������)��
�r��*V��3L����K����"á�n�g����T,��J,�d�=\\v�'w�A�b�ݯ�r#�x?F0� �(*��}g�N��C�YمcO3Gb�h����M����je��cr��( $�_�����T�B����*��YΉLa؁�4���Ϳ'�W�8mH�!�F@��#�[}���(����Yё��a�\m(�d��!��U?�Zz�B$���aL���0cCpkw1,��2�����Uo���UD�������sX #U�7���N��-|61/F�\������1���z��=�A�St0�v��ԊL�$�<��N�g�����ٜ��k�Rٜ�Gf��y�y�5��WT%��(�˔v⸽#n[jD�r*��4��ޖWL2GQҝ=
���Y�9�j���{M	�/<�?�6e�}��Y���o�i������|ΩT��J0O"�l�p_�d��5�SIϧ����t���
41�����W��ڕ1[*+CpE^^����xCc�
��Beʰ!C#�u`EH��ɪ��P�{M���@���s>�*3Z�9h"-�5�}ZM=k;��f��@>�EZ,�G�2����l�&}d�@O8��\1|�Ćܶ_������d������2l7,\��4��0x�������j�_OG��n��RB�*A}��Y��`��A�BB+��v��w��q/�9GO�te�
��`�7�l�ڑ��5_jv�]W��;
�*$�� �L)Y�,v0$���+���ٍ�>�^N�9���
�r�G%21���S���=��!$�'��FCD�m9�|�q��� ���>�������"C&`sm� ��A�����v-$�o1<Fʹ!?��ͱ�J+U�\�y`}��5� ��[������/�ӿ
��7]H�ۮD���-�@�����	��M�6cI�O{4A�ˌo�;�^=+�?�dz�1��+����d�j{�}�lU�1��z4�����(�� \�O4{��L�(\����0����;�!�'=�n�{�|s9�N�� |k]�;z�B��I�"	�U4y�����`N����̭��܎�	��=�j�E̲׌��=���>Pn�9�q]2����(u�bQq/�*A�'3JQI�HZ���T��F��BX��vS�۬ F��Y>ϊ����n�u���-�W u�M�9a�X�`��&�-�����-xM!ᱡ+��Q��g�읱���rvz�_���mϗx!��	O ��j��d��T����G���v�)�/��h]tE.Sz�[V�mh,6,U(���)��x�dI"As��I	h,?�XI��t,!��}bp3�N<ߪ��M�>z'��\��}���QM��68����5��O�d359�t��0���G�ꛏ��" �v��yp-Б���Q�r4a�Z#o-��y3h}@��,�F�	���\�c?[}��r�H]'l����G]�(u�IN���.k1�p�A;�$��pFz�X*����uw��u'T�v���DW\)���:�˥uĺ��ࢡh�7
V�ťD�dWZ�-,�Ce���M#*�����R2G��k�h�����Wߤ����a�*�FD4Z�j��WC�98� #��n�Yr��'�(?H0dl��_���mu=�!�q|�,���=(�0A�Z��9����!����,D��̹�����w{�p����. ��Z`�?�D��%�Z��Y�H���g��I�I�!kA���+��u�O�
�ģB�]��Dc��`�d�#����r���c�|��L"�;P�_����4ti���{o�v�������\/�d3��ɃsC���rp탴S��~{}�����ٮYEZ�&g���� ���Wϧ����N77?��覞_�:��I�E����@b�5N����Oa-~p�G��5����u���2#e���n��`ZP���rpWX)�p��@#&T�Qfa�F�`6̂L�MbJ8����m\��k���"(��D:�C�R>�.M���x�(��
T�0ԭ~ ��vQt�õY��v!��aɜ�;�uP������}g��XAMC`w�̂�^��t<�&��8>0�n6�J0J#�Ā��)[R@�tc+z�Zp���4�2:�)8J�O���2ޗMp~�3���]�ֱ>-��n��@�w���ϒ�t;b���	Iwo���T�'����	��x�ω�b�b����p܍7��Ih�=�A츈�eX�!����u�f8�ބ�m%`qR��1�(;0��H������9��+��A��S>�
�{a/b�V5����"����Z�)���<x�m`1)�5��+96�6�?�|��ϪO���S�cF!��X}�� "���
���Q"�jgx�͂��L���g4z+���9K��,�̖�_��Y�n)��"B�1�ޡ�f�vv�Q]$������z
�j�0)2�hjf�C�z��5Xi��rfH�2.���3w>"X��%e���r�����J@dj�4�.�"VD�z�6��$��~s�sm6+��o�<���mċ���L�+���.cAI'��tVN�0�]b��^�����R��5�(��=W���(v��^;�$��UŪ���{���X`��`Rm��[�
B;�%���v�m��ׂ�:�2a��}����}t��~Zb��T��:4D|A�d(r�FX��F�s"�-P�,���|v('xA}(�C$8�h�Yhq	�j�br�)��YTѹ���j\�!@��j^�5�ی��v�
�(�= ��p�x��tL�wNQ�`��n,g�}U?��Q�p�)N�X6�8K#{�`?U��8u�n',?ד+�bI�G�W� �G�����K�+�����<�Ö�����w��hY�NW��]�h=�CL��m�ە^=�u��U�E}7!����B��f�-K�ߚ�����������/���+V��ac��
a�3�&W�!a JSa�1�F�5Mϳ�	�=��TU7z�ۃ=�����*V�TVV	CGҧ�58���^S�������1���M�e����IZ�~�xvFxyW1�#�$[}��D�!r��J1�a��Q���n'*��^p1b��s�q������Yw}i��'���FD�6�M�\]�M.!����a��F"�A���0*��M�u��ۦ�I���V����0$L�����V�mN^�a�bL�q�P�}-8�y*2���^@�٠Dɡ��`�+���ѱ݀�-�jlag>�"'���0�rW2F��0��]"qI��x#> ���H�뜰����@����Ex�ħI���M�ť��n0��^��@>�ٗ���O%g�1'$��2)3)٦Yw�3����?� �<V����^�'!���m+��$��D���|�E��$�����7���w<�iw�Tٌ�f�> 2�Q/D��`z���o�I�=dϯH��F���e����zs����G��m���	�FF�ޅ5]D9G�*>�[�:��/���tW&�\�V`0!ݨ���ކ��kh�)~e_}�_��L�C:3_|N��o?z���͕�`]�IO�I���^t�:H�./��hg����-*c��<L��D��6�(8�U�"Z�+N��������t5If��/�����a�T������a+׽�wA���?����Rᦣ"���~Mf�Ó��E�(4��&�5,��`�Y��o�c���n9X��\�X>�Ն���Lw�
��?z�k�E�_dQ뤏��sq!`�F�nߛa�0�J@�X��約����St����zK�O��� ��6}}G�4�r�_m^��d2�GCٰ�S4r�_��������w���pY������2���E����v�þwU�_�H M����R��p'1��Z@Ph����+x������Ð����?�/3d�E�p�z_(y�&�w��ǧF�g�J��/V}�XK�i��+o#�չW�J%��M ���]7�IN��X>���SbR�d5#���ds�jq3��<��8�l+4���&�ˮꛉ�W���BsU��6�hk'��B�.�/j�&�2V������8$N�������gu�WOK@���F�-Ɩ�DP�|V����|��\��P��r���I\ǥS����(�5��y#����(�tъ�j��h��!��:�� ���L��ݘ2�'���'��Y��p�X�b�ǌZQ-�bDw��
u��3$�L������������Dm�-����P��W%���V�P�;t`vє,c�ȡ���Aħ�ʔ����tfe�2���;�s=�>���@��_��������_�w�c�2qlw;��$?/�Ѽ�� ��j�W濉Cx��a��B���t��(�1�3�z������&�����|_�խlL� �-Daf�C�bla,���dW��,Y�~j���<l����ui��Q]o6 El�/[�s���F|�	�q)F�
E��9ڭ���vA��O7��ܓ��ĭ.ag�SH���|)�$r|�6a�Y.8��&,��z���w��U��T9dr�\G1+�4?&�i��R�@-rl�NfbwK^�_�\W�R5�2`|:,��?�=nGN�� l%�]t'��;�2\%�� ưe��+�In���~+�9������V�_��:�G�s�Ѝ�l6g8��B�"1B�����!�B��8��ۛ���-�s����ipU2x3�� _��ciQ2`Q��sqB^��N.q�Q<�ۑ�'~{�~Ŷ��S�8}�B$�$n��^/x�}ghK�Z�-Wqc�_�Bse�&Q��F[҂�!�P�!ŧ��>c��h4a�v�*E>����O�$��$ڑp��UсPٿ;v�7�)\��_�cN����u�&�~ A:2�F�U �v;�	3��矣B���s�3m��N���$��_m١$$�evd��0At��(W�P%¨�?�/�H�$[���`=a��f0�Q)Uܛ���e�b
�X]��rҬ�K�DB��k;L�4�j"�,5@8o�+V���B�%�IX���{XiS��/��������A�!����>#��7c�˗p����!͈�����m��d�^<�K�ׁWQ5|��1A�21�X��¹��Z����oX6#/0m��k�/hU�Q��(��E�A<��,�JJ�R��9>fO�j�$��*�:���v�&����f�2�PrXDB���F�;��B5�E�2��?p���&>hL6}��p�e�Ag�f>���4����P���^�gf��.�d�o;���泽��-��}���N�AyJɾ��±.�KrO��E\�br��a�(l�yvCQ#�����Ɉ�p#9`a�R�Dʰ��Zū�P`ൌ-���vh�-qnc���
+]�����'��T�x��˒��;�����E�d�dG
���q��rC�W=�~��EН���]V�b�0��<&�^yL@��G�.�0u�W�l8��W��/T�!�6�"݂#jko���v��.�ߒ~��c���_zdRl)����L8*I|�?fY�l;Bo%{�a��<�*0�u����B��tr}��O�pG{��T�au?��] �u�mk��m�"�sA�ooo�;��_�w�)껳u�~���3�����W}�n��E?��T���t橂&�����SM�)�
pA�p+����o���*�> 1n�-3I6%#�AH[�`���b��o��7�H���<W�3�^�Ə�z���湶�\RNF�*��5e�h��csʴkr�~��R�ٱ���^��C����K*UK�D�m���Nt~�g�?�3���F/)�fk:�'8�P1�m��w&9l�X��{*�[�j���D�A��j��V%��Π����!y�9�p�}�#��7�4�������^
����K�w��4j��l��C�+U��
Y{tz�K ���P<�GV\�+�\��Hpx��n qb��,��p�e����-��o��A�6oc���2V��kF&ڏ�Jά�?�M.[�1@��1��PG^��5:bF�UG�_���!4fr�>��g��I�E�H9+\�XKQʝ!9J��g����-��0�� m�ȷ�����T���2�\6�m���Z0u����B�Y��0)�73{2��f�����zm%t�fق��^	�@������>��"��o��!�x�C4��b�ُRiˬ�|����9�ݴ�X�ގ�\ߜSg��Xʆ��䜑5�����ke8Y����[�B��{	k�Ð��ʀ��'0��~��x�$x�U�ߥ4U	�c43cs,�cqo;F_�~���������}�0���{��g��F�DH�M��!��Z���ptƠ"~/��	\>���}��9���Y/v��A%]bR��#X#t6n`x����T7n{q�rc���$S�0��m#Ialus��
�F���{���Ũt��B��|R0�8���b"��?��,������+}�������|i	Z�^7����ۢ�B�2�{q�p��Sᐚ&�Bg��d��/��*N�&��^$����d��	%�\	bU����7���m�
�E93E(� .x^�K������^].i��z}/����F����9,v��%ad87��`�C-�7Kx;��W�0���ic$�Dh�_!-÷y�x��~�N������ݘTP`�	�������\�[ls��x�s�0�r2z����57/S�[�m��WH�.���U�P2�蟖x���nb��!�@�6mr.ߊ�)����&�1I�M��Y��6�Ǔ���g���lc��j��r����_3��NTv������M�,aɨ�(6�w����/BH��R���$��g��en4�$��̅�z��(��=�����|��2 �p�_���N��g�k�
����f���e2\�D,{T�$�q��e��b��,�y���m���UРD�7�:_;`�����,m*����P�Zd���;5�dQ��8$zZ _��3���f�C>J�eH�;���7���ӷkJ�GF1��x�����P).�yE/@[�T3 �k���'��N���=�B�h��fкQ�n(-d�?A~���#w\M�(��9y�F�����M+�f �L�[��\����?��Bc�߈6��>QD�� �Y���E�8����^h�:�G�.3�Sjl^�k�<pٝ!n�Ի��}`�\�a9��$�����)�.:����I�εZa�z��,����ۻ|����/���h����!���V�`���ʚ���+��Ub�c���ǣ�w��@oISŨ�b����l�	U$!V��S�����$�NG$L���|��<U1,�=i�b(br��$����MBBP)�J�`��v"먷]�+�=�IH- ��xnQf�1�|�[@��A��7�����bJ�/�Y;�]�c"g�^�qV������v�ڃ�!��珄3|a���4�]�E�%��H1FE�,�|�"Ã��ͣl�@]儭��Ʉ��IW����8��Eِ�}N��V)~h�B��X}�mQ�i���y�Ho{�!q�j�*�d��;-�`5�@��jا�X�/7�B~\��\U��������N�?A~:���� ���{B���p@��՞[%�`*�2J�S��G�(6��l=�*!� .��d��͋.��,�)���<??�b��c���ɇ��� lf��Ki�UwF�PeO{cy�ac�%*J����3���#H��L�#���-�v��"��D)�2O�hE~�ӄM}Al�ր�Dj��뒚 w:�����aˁ��Q�W!=V�#ŏ����[YBڛ�P�ҷO�:�C��	��{~>=�R��7�g������uiq��g�r�����܌����rA���:4XlVo�&7%��m&������N�~�s��Ȫ�l�CR�m�W��J���>2�o"����l���ٖ�$
$�u�Y��Ot�4��W��X� P{��3���iRB��L���4�̧�5`���*�I��ƒf���1����i�mv���
�>l�t���p����r{$����J��~V���c�7W[K<z�h�ǉ.$�m��_#g`���q�g�~�\���	��d�C;���ZD_m����Z �NbY���$�6�D_Hs�5t���
�#������ɗLW~�r/9���y���;�?_	�$f��)a��{�3�@�w+2�+ʎ�؊#B�`���	�U~� �m\���TU�9��o0v�]�Aqc��Z�Y��n�P�C�}�Q�<;:'M/�e�.�H�X������߂��@H��E� �I�?�;҉�fN{�W촁8�a*��F"���<@�F:Is�|��aX&U���B�|W�=c�@�D����Ց���땝G4a��-�zm>��O����f����.G���
�����S��bҦ������V*(�SV�/H�SBX?)�D+�*q }� q�@�h�����ja㚂��H(,���v'8>v�pޗt��
�����d*�گnc��M�8j�o�9`겖���5S�H�/��hK��G,�	};�vĠ-�ed  �a���1܅&��6�{<*m1�����
��B�H���Ÿ�(�vP[0Tp���ih }�Z��;���P�v1�w�]��֝�oXE���pr�n8 ����X�bnf��E[�>،
[��$���	�Ah�Nj=�QJ�"�F�U�^<^%x�In�^z
̀B����C���	,y�EQ��u�	��Z]u�<؆�h��' ��\5|BǶ	�hidK;��@�T�����UJ_�?�TZ�<I��Uiag�ВKG6�Zk�C��u����m����R�V�&�P[�y{`��������sy���D U���e������I\D��C�%x)]�I���LTYT%�!��x��l�F/�@[A`">�%������.p��n��g��6!98;��񧿷/��C�`�F:'zGI��Q��Չ��˅]H��%� �aaHW�J!��8J�Jz:��
���9l^�8�p��W��}���r�5�^�\�����y׸�1��a/
/F���X��g{ʱ{!Y���z�P,V�i�p�f����^�T= ;j}��|�$����;ZZ��V���׌s��x|�����{c;�M1��O��O�ʃ�/n\�R$���]1C�E��Žq~�ؘK���(��E�1`/E����m	B��Dgr�%�W����O�xs�1 \�N���}�r���s��w��>�=g��5JW�ᅓghT��ߛp��}����?�[Z��\���_������y����Z��FS���H�%L���r��J����z"�~|^�,�`f	���#�G��n�T���fs�,%���C�N']1l!�V����}q���Ry��u��G�7;L�ѯh����wJ��>,��z	�R�2����V�{Ge���x�`74���f4�5�|R��.UQ5-��VkC:���g�C/���rb0�~�U|ߨ�+��x>Њ��x���瞦�R�D���� ���g�+�f?૮�����"���hj�H�)���W�6��=�+�CQR\�1�J�8ܩoL���@��\*���#o�7_˙���71]O̶H�S�԰K������V��y�A�	�c�}��l@�B�zOY�4�p�Y��'��O�	���qCH��'�����,��gP� qg˰�|q5z��H���fa�]'"S'}NX��A��������Ƶ���t�+D�I�]Ah�@33��%'z�l�a��B��-r���x�μ� �_���I�;��~6+�f�Q߂�8&V,`���pJ����Q�4#�a	�1`cݫ�-p�����
�se_T�#Kǝh7����iۣ����w�����^�.=��`;���o}w�ǽ1b8���� ��?���ͨ�AMR���dV�9M�W��~��aB���'7L%�џ�z�ʔq�餉Գ��x6�߿�w����a�8zY�h��5�`�y6�BG��C�,��U���1�]��58<]}c8�
��\���2s'\�!��aq�᳻nO�.½��1�N�Q/V� ��4�Ƹ���wF��J�?8B��l���d��f�ђ2�*��J����A����p(����:�@��|�VM�b���NP�� ���+a��`0!�Y�ؘzus�ͩ�������#���@O�V������@zMd�4С9C����&h��A����MS7�Pɢ�ۼ7Y�`�����m�����b-�����xE�F�w�$o���{����gZ�W'VR0��I��`�8�����C��K@:�S��hv�U6�b����Rm�
�4\��$9�Q�F6�E(�\�y׸&[:���C�sE�������� w\ܲ��x1��e�K�1���4w�+�O������Z��XQ��E�R��9��pRz��Q�42lB���$��$�a��V�Q��Y��^���'�1�,��ȉ�9���0�ä%EA�[׷9U�y�V*]Yi#04�ӹ'��4{�P���{��`R��`��U���j~&L�Dva�$8�UJ���93�j�w��=~t/A^}{���8�o���_���Ӣ/�`�
ܥ���˝�#z�_~�RH�P{��g�9g�J��ҡ��wI��AR.q�\�0�]q3��:��ѥ?�V�N)���~���1�AV�H�j��������T1%�b�� �(�}���X���c���Ү��Ө6���W�=߽�X�[1%�T��nx��얙����~�?�8���*pw����FM��PEM�Mj�ȹ]��U>�@_j����������y���@�*������%�؉�ʌ":��6\	Di_ޜ�o7�G�R�U�������k��(QE�dP%*�`�}�<��E�����hkb��*�`���|�gyu���C��z���sv������u��AfX�1��s!5�I|��Nt����N'���C�E̚T�au�`��
�b���~z���ԮbX�r*��lL�����qme��j�f����>��k�h��d�
ErX!��� F	��7�-+�1r�"�[�]bW�L�ڮ����q�+j������ZeM��HM�>�f��\�ؓ�������b[>j��4*��΂!�����+t����c��8�F=0P�eEe���;�WUU=����ڸ�S�����-��=	�N s3s�O�萚?��YT1�:@�sjd���#y��[S�&��\��yN��R�A]@V�d��(S�Qbz��!���i������3�wOK��#��Ju��>O�(b������i�"T���Ea^f�覷=�	L��?vqǙ�
��P���N�XH��*�H���<5D�e���-pl�vؽϑ��C���/��:��f�
,��Ÿ�\ؙ�C�]�(B��H:ϟ_�#.�(a��� y?�g��l��r���3�@�MSx�"�.����2|h�>��	b���K(@]�KyV��1FfymF���,�f���ۏY�[x9�sJ���|���?�W�� _��Q�eF��qq�M=%�,��>��:O�L���
iF�y�LGU��0h�A]�]z(�SjT���"=j`�j��{v�zp2I̊��� �VC�m6�@��x(QT.�&'O0Ģ4m<�X�?�g���o��*��*	Q<�,�$7�RmI�q�F�Eᷰ�H XKP=�n]%>f�t�^g'��*.RR��%��iҊ��`��b�拏|�i���3�%�x�^^�V���G���)1[b���h�Cv"�<��¾=�6�i�>r+yv.6gæ�_h���g��4(J �)�`�a蘗�v���_P�i�L�#��K��o�O����|�f�9�D�Vi�jM%_4��і�)��֮ӽsi��xؑ:��D��-���+Ȧ!�(d�x�	��H78Tvś�`�
�$f��ެo�E��r�����}�&4Iᣣ��!��<���&Sr4i�$U�4u�}@(h�EN:]lڋ^�Y~)H�""���m���!{:�?]�ވ�QkK�Ru��Y!��<�G���y����Z��գS�C=�&c��-�����2���O�o�<��=Q�rE�9Bγ�� ���v�z���
��}����?�e��F�b\s2��.�o(j��>k(+��c0�il�3��%$0T�&�9 Rw7�i8#(P�N/F�t1�mT�"��Sg�;̀���j���?�� &�!�
��U8���ܒ��}%�� �`67-T*#��:z������^xa��@ ׾��=�MS�ݶ�<&����w��8MRi��t�[�W����{�}=�#)t�i}���ǫy*�U���Ӓ5�4QP4�g��E\[�6?\��%�J5��S�BFj��ޅuP�)�N!r!�����6��t�^4�
�L+�J��
�&�@�D|��������X8�ý��f"%���ƺ�����t��&�<��5���tKW��K+��@m���b�c:iZ^���qv��)��L���ZN�4IJPJ���o��ҞnV'U�)xZYK;l�`yI�0}d�:�%sI�2��$d��;Ѳ���Y)]���W�g�up��d!�n5'NƣT�O�V� >W�����yq�>�l��1~��S�ߧ�~>Z�?s�-����g���z�G,��+1�wFz��I~�ף���B��J��)Ѧ��ԸZ�Vh*�zՏ@(䞞��������+w���r7ŉ���������U*6�Z��l��+���%���M)�b#�������
vu��Yw�Z�ed�����&LuM��49֊�O�;�訝gV���U�C�1X�]	�C�^3�5M���>x�c���c�I'�� nZSV�%բ�ȏC������k��b�}\F�+'K.Q 'h"lP��w+4��ّ��)�� ��N��΋�'`6���vZ?04[-<W�	��h����oJx�==Uxŧ�������{5�y���6�!*
�ì��� Q���ﺨ���3l a�/L�4]�Ӻ��E��Ŭ���b��������05�A$$�mi�� ��f��k���t&˲�Q� ؝0g0��c�âW�s`������	S�`��cS��$@y���.ؕb��؂�Aҵ[���L�b.�vҀ���;����J�T%<R��P����������U�Ы�+���^�����	��i-�f��S|����˧�
��z.	{��ث<b�g��.4��!PE�H����=`7��.����H%5�	�ְ-u%_<�l���=��BL+�O�G��q�����y�ʦ�x;W�|j�|�ا��y�}�|��<ۅ����q�E��<QPW/��R.38�}���+�x�~=LV8P9��4��<JU�c��1���F�Q������i��_���*~1wC_�P|_éΗ�cU�ڞQ��ǚ�~���&
I?�K��HRC��3��l�g�Y�e9%I��vX��i�L>��]Y���J��8]椱q���Sk;�}^���`Ee f���$�T!Y�l���H����j�;�2�36̧t��w|�'|�xA�K�ps�;�����
�u�0	�Xߧ!3N��!kӆƖ����gH������:Z:(�E�^'�+���P�4�`C�[_'s_l���ا5A:1�pMQ��C��v�}U8�F�~B�C�T��.зU��;� "�8�i{��`�ŵ����z�q�������� ���~�Z"�y,�eڜ�������k�.�;�L7 �qb��w�����`4����q��Gf�A�����|"���FM��٩��89;pm�N�N��g�O�(U<��$�;�7��� ϸ�s5�p|�*��j���¼�VOW��j2;"�:)�t-����K6&��5�=�AU�@��ЋH���8�c�qT.�&���]��Phۓ\w�y8+���uҸ��0�U�Mb;�L�|��~*��A��.a��t�� P�=HBo��֥��GH��E�ڌm��W�G�d3V�qm��x��UXR!�~fRR�+�"G��j���l��Y���},��Jy57�����y���p�AM��l8��({�����s����|��/�K�z5ܸt��~uu�,�#T�:��M�dYJyF��
�Li��Q��<�K�����e�hS��s�̲;�+N�e��MS��"�]!F)�/Y����ho�M?���4	�ڤPBz![׳3<�F��]�.u��E�6tp�h"�ф��%��qU�hh	���vR����Z:Y�hd��j�nMO���ȓ��q��d���SS}>��U��aΝ���ز�hݎ�F�ZM�]�/���+��A��A :�����U7���g}��.Rm�`�h[ X����g�� �t}4k��b�ߗ���E���?G������g�\��
��2��w��<,��שּׂu����9����C�Xk<�a�!��;������k����
%�p��"#��݌&-p�� Ym�������A�c���\P�c�'��A$�7x]�����W���^br�G��R��@\6,��u	4�3j�`�2.7�f�;lh�] �f��8�6�#'i��4�
���s�~��V�ħ%�vv;�"q��VԊ�䶁[P��~N*�vK�9��[y�y����a���ʇ(��o)ip@J)G�$D�FB���!�A��;���f`��;�<���<��?�̷=��k�^���>h�`��ML�Hj�k�QBfv�F4�o�g���1O��>Ҩ*��� �R�)x�+p9��S.m��ּ�u��v�����(�����'dk��	b�r��m Ϳov�o;���{x4݌����(��o���޷kTb�x��ۑ��M�/?���^�;���
s��-��ZvJ�����k���E�g�[���g�0�b,��;�K���?�oq�(�x1Σ��0$�SŰ���Ν�c���"�S%���q��Y�Ԡ p�.��T�����d� x�i�<�v�yg���5�_��	�Ŵ������њ���o*!�2��YNC�~�k���Y쮙q���	Q����V���}"��1�"��_%5�y���S�ʡ�w���9�;�w0&&5��(把��@峵�{IH�gz���/�~ �-+��t_mXT5-�c!��W}��їasa���I��9�q�+�޲�p��j�_m�*-wf"���tH�Γe$Ap���1�H��/~G�������@bi���y����6����ZL-�n��H���GM�,;�en�/~���v�aW�tęt��[i��|�V���3������Yk�h^���f�T)�rS���xl��3'�YG��:�,a�	��2:hy�|ʠb�W����k�^S���0ް'�t�ܡ�^�Y�f�UF�Y0<��QL��ǌ�u�2w�j:��x"�(|n�?|����C���z�)�GQ.�b��a25s�e:���oM�?��+`�(HyfF<�={�~���{a)źV���p�����iك×�������W^;�2��;� "�X�k�ə�A�u�c�4G,�2��#b�hŽ��R�1Ox ,i3:�NEY�!!�}�zȦ&�c�Z�ǯ2�	^��w�9.y]���*�?�֯<�`J���O������JE?�Y�2���~��{_��(3�_�d
?D�+��4x�O	�@b}��ϰ�e�T+G=�K�#@�'�-ii('Z�}�?�ـܜ��3����C��|��
QsZ�X�������H�p���b�S��1��7!����=��bP��%_�����Th/��0��AL�*#��]�.>������R��"'��-pR}{P��כ����? K��z�Y�.j���5a&'˹�-o�>�}@u���w�+$�� H�֯�8�
�B�7�Ae6��<�.`���>�s7�S����B
KD]��||#�d����Zn��3�py��)��v�za$��r�R�*�'��1�ҳ"}�_�\�M�����:�~+�)��/]��1"%�mw���#�勎�8��rp� !59�E�v0���^�V�V�l�7s���qWM|�����y��4���z;�boAQ�x*�����jĶ��Q�<����~b�PaD��gI�	�ү�������P���W�',&;%�L����>��?p��K��?OlfI��ʠ�_v���e��7["\�m�'p{e�~ټ%(��U�<�I"&a�v=���r����L6ߍ��a(���������T�̇�}�6�î"�H#t�NS12��G,��CsY��D�ӌi2�K��%��~��e��G�[����;����Ê��������6	[�Yv���5�ĺ��	�s��;	�,��% ��%*�YF�*���?�сg�>=(������վ���IJ�I���(M��@������JX�yuޝ�FԨ�8�*\�v�|(3P{Q�B1,}��O͇RM�b6��>��hxm�)�o�2�.���nF�/�����btj��rW�i�i�%=���[{���3����z^�NI�;�m��"�xO�6q9����8{.ɦ���s��bU�Ys�w�H������ݖ'��j�Зx�����srD�_��ޯ��l�LU᭩GBC��4�`5��a���]�ߧ�-��K���7}�K����ླྀb6!�X	����[ؒH���"��AE��]2�V~1��KuQ$���O'`��/Dra��4#7~�M��o��9Κ��l>js�)E S���,3?�1c��)߶�M=F�G`���Pt��j�@���sz��'��@�9�!�]��F����$M���Q ��k�9�:!�AVt�f��,�x����<fw��֡j.8�ƃ�a�˨tmit�=m�2�<�5�s�Q�����}�nyY��Jphc4{z��[�Y�Ɍ��t�|U\Klm��F�63�]p(��Qy�����o�S��m&4G�!����+|���`��[��t���F:��R�=v@-yֽ�qj�ud~�"UA������`j-i��߸K�xV���!\[��:Q'�x	ת8{�f���s�m���͙�U�M㐦<p:�r���������.���f��<�7u�w��ك~�%��I(�5��37mg��8�M������6�~�R0�t&�!,��kp[��Dl?��l}�gu�ҮyY�Y�)}��b������;�G;H�8{$���.�IK����m��>KT��w�ށZ�^�[�X��OD�鶋 a#֤? �7dn���쫻u�/�'i�������m`�(��P*7��T����uUu�։���{ F�o� V��{m���я'�Y�r5�6!�_��+N�J�'��7��L�t�{H��DQm������ww�Wؖ��8�H*���m�?"qKd����L9sl�v��s��<��"ZQ�z� ��[��膐��{�p ��4����>Xh�rvrb�k�piZ�e|9�h�j�fx7e?Uzw.�&�|4U�\����`�Z�[E���M^z1���]�=�o�{.�3q�S݇��A���"����!�`�~���K��� �eɦM
�&Co��+
xӰb�<��:��\��ܠR>b�p��yҙ���]��U���a=ISX�ӫVQ7��0��2خ�S�0����?����H�>]z-qˏn��и�|���4��D�%iV���X����n���m�_�
+�e(0%%=R���f&��O�Z/ٓOٓӧ������}���f��X���蔦OK���)��@��jj�=:3}��P����^��U�}�-a�b"h��(:YP<.�ڏ�����[�����]:A7��o~�X����t~Cv�pb�������B{�D���Ł�j �=q򠭗ϡGGO 4�v��ă`�=���`DA�r�jW�hI-ᤔ0US�*^K+X+q8����H�)g-EE(��*�?�MG���-7�V]z���ў���򁡤K��U�S�Hb�S}���2R��f��[R_
^~.����a�
~�ޣ x]��؏2����	�Qy|o�'-MM���@ߢuWژ#��|o��d�\�4�um�oH����:����g\ߗ��4�n�b�q��}�k�w�~�*a7KOGETq��G���VK�?��AҾ������f"U]����ڝ�V܅`s$m�ϓR�j]�^���2����*䯴)1g�T{�,嗳�	V�2�H���?L߯��# 9KM*lͱ �?97?�x��1���]�E~::F�3=�7�l�Pa��>��=�}�㛍_S3�V�WՑ u��?y$a���:�����3!��R��s�����>|g�b]�Y/xMi��ăP�^��[ʚ�r��!�����&����U�����I6o��EÎ�9BPj���ti`�zݚQ9���33���2=/�9�*��g�7׵I��B{ӝ�H�H��D(s���)]��ZO��U=��������82��	����ׇ�v/C�%|֒�,i+�g;�s:��L)�Q&����p_d����&Qi��!�{�w�{�SO�*0�>�������� $����rh���9�K$�������I��R^Y�t/40���%1��knN�S�����M�皮�ȩ>�.�,�Y|�ӢG|&x  � �:�y���ڄ`=�xs�PJ�&-��=����}�=T���C6�Xm�&��a ��� ":����o,��(���~�T�Z�CF�J|�9�����%���F�q|��ͽ����=��I��#v�Ϧ��+�2O��ZP�iЊ J�����B��}�Q[��7��0w0:��T���_���,��( &}
�DҢB���
Cz׀�LM�?9a�����Z�D����P���"d�%�T��=��FT��m�QxOCC��5��#x��-`�n��^��B���f�K�)��G�S4�O �����W�P!%(D:��[����TQ����)�"�'�ӏ:m搔��5�=��F˛���+c�$4�H\"��F=ƌ�E�P�ݗ�ޥ����r���L_?0�`;� r�#�M�PEe^u���g0 ��jJ�y(�fb(t��yG�ڜ�����3���EW��ɞ��"r��A^�����0�l�QL�۶G�j+�E�Td��Ņ>����`�3Z y�(bG㈨��|���sqT2RU�P��佌?fY����X��$(�t}�uG�Y�0�ҙ�JI!��Gr�<�L��j�� ��;��B,��]����g���җ�D%���s����y8��l�$����q���^����4�r�4��W��:N�o�#T�\�'��mwv��u�Cj�L����@�0�@�nD|��� B�,��Gκ�V�)�'�/E
L�g�l>��ە����Ҭ�)YrB�t�|v�T���+/��>�>��_��}�C�̟�kV�8ݶ��<��nn�TcB�}s#&��g�v��&s~CW)unjn�m�y� r#���)�K�M�z�T�%9�rf���0::�3N�ej���G�����-���c����N���$����ק\M�J�[�煶�H�Og 1$��Z�Ej�a�]�z)(ϣ;�a�RT8�Jsӏ�8�(��}����� ����H�&�x����)�EݳCȍ6�Oǥb3���	��!�0?�#J)řSKD�-�B��1����ڻ_i �s�p/�����L���n���G�&�`0��W�鏧
U���B3�p�v�ݨ ,�sc���u4�dɡ� �EH����Z�<�d�� ţ�4�ϔ����PY����2�	"�u��ʠ
v�k_lF2 Jm��R0�pP�2C�M�|gmkM93R�O����``!�a!�"
�4PK��B;A	3t�X��"8�W��m�H�R�Ng�se���6'�z�Q��+�`�i�rC�r��B�$���j9��8n�����"�v��k/'V����U��4|���F����u�ym��R7jگdCsv��h��&1��?���k�W�aHf�d�S ����"���U�!JH�Ӛ9���
�`J�5I��H����KT�9v��?��qI ���bC�r�!��G�/��C� iwa�-���������ͨ����%����՘��Nɶ���mE�u�1RK��b���vފ�C'sVnv�ĕ"1�sq>�0������?H��ݦ6�����&��y�Yd7�*�� �� �J�h�J@6��1�5�S��L,JAѨ����.�s^$�S��z!�CTC"X}j0h�k@�.�@T�[. 8U�(�s��2��1�L�eӧ�ə�r��%'h�X˾ȋ_<$�?�֎j��c�(H�69$�S�xAE�):p��?�9��oi��q��UuI��3R	���������_U�U3����LeBh����'b�:[^	���~V�w=�/����)Y���d�j:L7��.S|��xI�G�F�?���^c�밥���,�,U�s�ڒOH�ȶw1�_Z��;�)�a<�ef���m﬍�&���<��7�.+���n���?����pj���A��"��")1BxM˧&^��f�-v���@	 m�a��m�7�6}^��ie~w����q��Y�C���·�v�L*uE��S��h����!�$L޷&p�
�-$ykU���] E��k&�d�e�o�Dq���U�<�:��K�(�N����$��Zi�۞���F����{>cDd� ؤd�����\-��]`HM��ؘ|��}3I�ev799�F�!�Ph#@;�T\�F:�Ȃ}衻�M��\�)��ʋ�������������z:�veq�L��̵��5���R�I���0�����rQeӈ*C�����X1�<E�1eҐ�G��=�7� ��P[�����S[���`_ kV���*��f2Y�\b3<�Iʚ�R�/�p;�I�Xw
Fd��s8o��҂[�Ιaw�ȼQ����'gf�B|��2.�i��8G�X�.i�yd~��쭗6)�xgƹT�C�;ZQ��S\����,�a�+3@�o|\������TY�K��R�?0)���/�T:���v.�.�\~,Z|4��O�ɥ����JV�l�����+Ҡ������[A�8[���[���,\I��	�O�p��1Ϝ�^5�yQ9�ﳯ1��/{�qon���ʃP�	d���ydNS�Y�VM�{u$��B�.�E���g�VJ-O4��R(=���t�����o9���-v>3Nv| \؊����.⵫��̐*�
G�Sb���ٞ�������͆R'4��G �i������eם
\�[W����팟>�#�hŀ�5����蔎-U��8����j�9_sm��p��lr�i��W0��g�v���h0;3�#�D%�l�F�b��z����G�8
�*(�
f8A�I�Yu]\�Rs��c�lt���N�W�o/O&J4��w.���N�=�W-g*��Z3y�_�Qد/ T�ĥ#��L�Ld��J�n�j�G���l�1P?fW>�LDOa�d�}�����X6�K���_3<`��Hy��OMt�_��ʧ�AHߗ�9�B���Z�:i��yV��8�V��,wO��s����e�B�gffZ="oxxP��60!��k���u��O�c�EAZ�
{�V��]I�m���q��.�x���ZGX�$)b�T��D��{��OR9��*���2<ݥ +Z0}C=����%��z,����]7���R)o�<:>�����d�H{U��*C��Wb�9���P��(�)h�"��fh�LSu�+�'��n�OR��7/-&JKS=��A�crb���2SB������%�iWNys[7~�U�W����2�*�kO}-Ο�R/_�iG�x���>�9]�
��5��K��M"�aΕWmb9�R֍��kG�I7�:NO��:���W�g�K�D��8��TP��^�:��F��	47ѷ@�=������0�z1m ��.��p[UkX	نE5I��ݞ8@�#�Yv��D*���l��~��ɼB��ж��<@D�7�sy���I�3��$c|٪�=�"dw9��
X�H ��ƫOΪ*ڴ�D��ܸ���ӽ����3��Ѹ�����T�m�ѿ���?vj0�!3j�w2����bKčj�L�$)2��.�صc�&0L8�R�������+`qz8�D��� ���*T�ݠ�i���]�����ץ���zا[UQ00(�)c�H��JUe8��+���X���|)KŻ���q}�`��q�Mƍf��A���Ř�u�Ut'�C���� <�0
��U^i��z��9���?;��p�]\�X���O+�y{:��(Z�᭝H��S�݉/1��j
��=0������t��͛���Jȼ��kQ�x���2]^�33E�ŕ.wK��y@��ۍ�R�-�������u��.�y u�~�>�e�S�1��fe�xx8h9۶_���s�1��\r��}�I�~�S���+��c+���>We5������ �B�����r�ei�>�]�
����4��J�y^�Fjo���z��%�P���7���s��gס>7���..�&�A�*�]���t���4�W��������|a��؇v��V 0(�^���G+C�y��X}&_0���(gV�	=\F�6>��'^��p��U��Y!\��g�'lY���d4�b=*�pþ���V����g�dd��� �M���^�U���H�g9T]���Y���!?u)���?���;9G='�FTr:Ds܁ڸ�"���	�|kiiiׁ˳�ͦ�\︥p�����p%x1m�z�Er<�5�,Fu�jt�p�C����L�5i�$��W�yT��C��[�u�!q�5�I:_�>��n�Vi~|�
����M�s,�Xt�R/�����E���K�R
��aC�h���l1BZ4&(��A����y����yQ����� ��t&F����@���=G��g��
����/��\�!L��m5�}��h����[�vF��U�F��q�M�("Q���$�}�1FD}
r.�W�/�@�i:3'G3X3(|!��sܔ+��.)���?  :����y$.-4�MדT=�:�_(/�E;���
mCg�(�7��xo�?j?I~��.dUVH��*@$��WHa�+�ԐzQ�␑2�4}Zni���މdf�����B^|���w7�ӕ� )����D��Q�Bx�������%�_�-y,>H�M��t{Z�V0��~,��|�]C?�м[�4�^��r��L s�d��$\N\
U�dvn.q94\M�)V��v�\��S%�<�I�We!B�/��� ~�͹� �k�]6
�&Q��7���i��_��>lG�nh{ۼ���~[-�݀!t�PF���F�s��֕V��8|��O ˺����MV������(�rp(���e��</�>�sk���o���������A����*�4u>o�A�N�����=:ry���m��B7s*�$�ě`X @�`6rn �3��5�k��#MLm�9,�� ��ai����$@�_'�?�l���Jk�~�(��W/��@*�v�ܷ�b������kQt�Y����_90���pN��feIJ��F2�w,7�-
^�YI]Z
g}��T��K
HA ��a�a�h#!M��/�JK=�o�'�
��9���V_��!��Hi�#s�=�d��%r�>x\�d65=�2��e�������9��"QN2 �*++�.}i����4㢋է"#����űs��ʘ��R�f��{ "�s&T��qH�g��GQ<������Ь��T��f����Y�/K�V�w��B��]"��K��$�uG1�<�����X���¡� �9�LC^�7[IY�����y/�r�L�� xؐ����hv|F�q��G�V��d4~ʎeC�B�N�^�۳�J8��_��8~'e���4�������l͜g1¤�2�VM]�j�DT��n#qI4�)ɪ�b�2��=Oy�a��f� ��,�%��UQ(4�}��R�/Ȍ��^�(R�OP���2L&��o��+���H�|q�In����k�edڧw�s/�%/�K��o�U�̤�������2|�/?7�����ۼ���ʈ[�#�j�h����ð:���{O�rs~t֍+�p(&�»68�ky1:}��617[����|�`��j�g�'ܰ�7�f��K����B�Z�m#�CQQ�
r�� �dW�5�y�������I�H+5�tݦ���\Wz��aQ�{͢ی�_k��ʶs�����y��&��g�hLz����c�q�x;l	-'�	V�ۉ��*���=+):n�-iI�)�y�{*A|�KRJJqk=n�@�ǧZͧz��:�j�Âӷ뒹k�Wv�ӿ'��/����*�^�� x��N+��7~7_���Q��(���E���M,�K��-S:���#�ߢ���uD��� �y�������M;�>��h`{����,Y2�.ƙ�˪�˭���� �lr�+cR9/�!�Ŧ��I��\�å����f�Z�.�l��O���%ƅ�V��n}-��;��x��u���x�ۼQf���2��}��-Mq��QXT�pQ�p�77�#�-������	j�.%��*�M�[췷W�TYY6X����dc�+5c
bb n�q��{U+B�%?��Z����������������dD��ĉ�lb>n��\�z���j��X�}���͜��T>����C��׌#�T��8C��`ș�2��q����d�Ϸ����W�$�!r:%�g�7�;.����/�zD��A����np~D�� W��I���Q%��0��6`o�e{T��m���2)G�QGiqR�k���+��i�&�U��c&K��r�w�s�5/�����|ށ��=pY3޵?\p�?�l�w\Z�y����)�B"#|*�����}N�{�϶���'�
�}5��*�ƌ:)�cp��sԁE�=;��y�GX��ZO�+�v,b,F���˥5ܩ�؎"9}i��^���p#9J@Sl-���i�7(:��E�߼�!�_Ҥ��0}���lM���Ѱ�i�iN�,�Տd5�� ���޷�� �6��8x[��/�/f��m��WO�G~�F�p��<a�1Kow��Bi�S�(�;w}�p�E-"{��m̦YI-%i���ݎ��Zn��|,21Q�y�������jF��6Ȁ;�����4�?[!7]�eeuy�A�Ui��ve<&�KN~#��O��d�j�\++p�S�G�R�;���P6t�_WN�9���(�߱���<��	�NU{<��3]D#����)�[��k��3��K�z�q�˗B����0�M�|���!��t$�y�s[�����
�M\/��6��|#��)� ����!ܦ��^&�* ��
ɵ.<��d�	��J�?��-)�F6����0�7B��g���9"y��N�wu��;�űb7���P�_�r�U����c���P�:������`_�E�s�����k���(���Tn��VU|���L%8,�p��Q�V\"dE*�c��X���H�.�ܠ���Jo���,�)�����}���������x<�~�����0y��2�=�ϥe>ywI�����l7����t�nљ`&v�Q�.-�*>����Ә��[S����ׂ�7WWSPƋ������w&{�9\4yQ��r�b-U�����"�6���y�D��O_�%^E���`N.����3�W�Kbm��?�q��I��qm-n��h
�R�a�c]w�)V:�]��j�J.?�g�Lq�$�ύ�?�#�4����@��m��&�Uw�uB�M$�K��ʕ=�{Ӈ�z.k �A�=�g����>��յM�s�cI�����%��b���)E���VM�V������X��bW"8ު	"p}�hE! �;n�SY�/�~�P9T�5�=�%ѕE|�Z�sҋ�po�A`���nR��"VJ��h��5�D@C0f��ÑY��	b��9�R޿�7���Zn~���Sc��Կ�5D@<CM�?��4O�S{�P0+�5Lz$��"����<L5�E��C�H�D=��:S�aj�|O�_���qdc6� tT��ԙ|㮿��ރh{O���_1��_1��_1��_1��_1���G�{a�B�u�=_�G�����x�;C��PK   �<�X/yR�c  ^  /   images/d2af519c-c065-45b5-bffd-6bf239de2b90.png^��PNG

   IHDR   d   P   �	��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]	l��gw��c};��ΈU��ф#H�4�� �U�R����HU�V�z� �rD4��F��\���І�p8�Rb0�41���X������lf{vv����>�g��f�����������*�8ˏY&�d�xY���/�m\�BQ�6��#���a< )���������������~��f���rݟ���M�s���Ȳ���x= �IaB�� Zl�ۗ��������p�I���zV��ˊ������۷��v��/����,���$1�#L[ 	����t�ҥK���_����Y@NN�;wn�RRR�_s�â�Ͳ�e�[,>�7�AI�5DĐ�ˢ����I�&��2�M��	b���j����͇��cg��3,����r�x@c�0!W�\�[vG�p8���/���#�)��Qr��>��3L�9�e�OX6�FN�^(�1G����:joooHKK���"����.ܻ�e1�wYv��(�S/��t����P�������;D\I�Y��;,+YvRT���h�p�Ȼ�������Ғ3x�`b����M	��*�?�4�@�!�R�?x;��������/4A>��E�Yǲ�4W�{��(�ۉ	2n�8:~��~XŁ�Q��UWW�C��������Y^e��
&c�MFyy9�]��� e޼yqՏ�#)S��kg%���㏗s�=m���Ɋ+����
?o.?g3s��qLA��À�"V�k_�n]\�8�OI	���a��ڵk�9+2d9�N�&�|ʔ)t���)��@��<�zۇd)R�)���d�x���F�O��dgg��W2�T[[K���b�-�b�O�>B`�[�{������p�}RC&�6�gXo{�!��
b6o�L'N�S�N�p�]�}���Ni1w-�u ��ѣ�\�������h�ر4|�p��ʢ�S�Ү]���=�R��`8�)1���㡊�
�Ng�QSSC^�W([|���)4!H�"�T��u��bK�)wYY� %�� ���w������1		qdCo�B�p��R���L�'O�dXq;x�~��i6l�p�S���t����DEU#�)���y�2��SK��י �`\o���bU��1���@q� �Sc�����̌���A�Pt�K���7n�nJ�S ��Յb��[dS��o��f�q�V�Q��2(���]l}�4Q_?F�~l��=�������F���u8�)ܛ����R�2-�W�^d���is�uD�NXCC��5e6�u�LG+=9t�;؅����j������)/�y}����D�?蠃��G��M�L{��P�/�f�Iv[����-���p��N+�n A�&��y+')A�ج]J_�p�-�c\	N
̘1��/_N�������e��	VBA.�qd�̙��~I)h�v% [�Jo_�25ys�R���ug;=��h�����=[(1\���TO-���������tQ/+��2���Y�q,��!���l�U�������dy��V�WLt9����'��IA�0`�Ha�]�d	m߾�������`�cdn/��M�0!|��W�
f$�G�|���B�����a�r��.QN���E��S�e�l�t�(��9?�f�n$���,��4�jNO��"t$-�����A
Z<�pa�c�ܹsE9b\Z=������D2n��Ѱ���RЪ�����\A{/L�*�B߻<>l!�*զ)��qd�����.�a�7wO��n�f�=�<����nR'F���@�$��R��"�����/:yP<�-V�.�0ta �3���j-]����nѢ�lXHt�bq�C5����
�B�c�X݋Z|Y�V�T�����3�x� @]){��$�]`�� ��E"CF�v���`�޹�yp[pu�`�)�6�:�.�f����.�d@y(3[Ay�禋Q'��]U_	i�aAqA��ߣ�=�v~83"�{�V�,��1	]�p9P0������"�Bl!dVp] ���*�!��9���6_F�֔��Q�^�}(<�Z(�X'\n8}M��(
�Ҭ�4��2a!p;��mA�1z��gg �
��X#�fʰZ�Y�xϛ���1	ٸq#Z��髊1&��D�(n1&V�n��L�����Q���ƾUg�I��Ç�Q0��p�BJ��;!2�����X �C�Dn��ʕ+A�ZZZ�$J���28�T�y�f�}�>~ժUaRt%n0��TX�c<^!�,�IQ�u�����%�@�#�MT� ˈ�E'����6�=��z��B0�٤�H�L�w����!��	h����A���'�ǃ�	��SIH$�	뉢����!	��A�9�SS̰x�bw�@�u�������8����.��$���Y�9s����e˖)2�Jʃ>�zNN�M��֬"yܬHH�oD�F(�E�`�A[˒��e@�1;(1	n�[E�#�$����4���0xXPP�̟?_]�z���z%)2�?�p�\J�\��G��`���eI��X ����;��Z�;�x!ř� eŊ����ۡ[�СC�"p��c�xԨQʢE��M�6��d�HpV*^�q�UB?7�|������*���4�u$?PLՑ����<v��1hXb�q�̙1�����o�6��i)=�f�4к�:����yx?oڂ�0�����{����z<�=�-2#\�F�H�{���z	�~l����gY���O��h�uf0c�����>eVl}>�d��K�,ccU��P?z��k�Neǉ'�<�	E2vt����Ԏ��[�n5�V��$!�!:
����$B�/	I!��=ѧJY�"m9^,�!	Ijk{y��?��Kښa/��.*bJ�$$EX�tӫ���XxlK�dXb����t30��fڲs�ӣ�ZX�f	o�MZ/^ZH�C���늟���w�ÂD��&��$����38�MXXC��XK{5bU��O�諟It'0�T�vMu0Ȫ X����/�~¿"��t;LQ��'+}ݠ|>5�4��e?�v�߰%���?|饗���nX��,"-��;8��,{YvKBR��_+��wi.��1b�|IH
�ي��������_=�3�A��,��|��Q�\IH7C�)��+W�~��XO�e&��4ik�1�=����nF�UX�h�ol#�k��W�he�g����-$`��0���RFZF��F�e-���PW�`�ΨQ�^����>Â5��(�|6*<,	I�m�ǌ�>��e�|������,��V����ǉ�H�B���z�����_��V�B�0�.�|�4��$|��9IH
�q!n|���k�}bj�UB���9�X��]g�0�����V	��=�Y��D"��Κ�7�,dYb�|����$)�d@wm�����0)O��)B��fA���u�u��l��"��`���N���x�]?�~���&�e�_w:�x�$$�|��#G�|�ԩSq������A8c    IEND�B`�PK   ��XMi��.� w� /   images/d9f6b7e6-de48-4348-9514-eb3e948015b7.jpg�gTSk�.���Ki"��eD����!�IX��Dz'RCQZh���!���P�P�{g��>g���k|��7��?sf澯�~�2��̣��l��;��v�׋������ɓgN���sܜ��89�/q^���y��>���._������wE��������ވ��]��!�'�|�̙��v��3�W�8Ą�]��! vML�_F��U���b��BW���]��v�O�_�O쪤(ߵ�G-lO��:9u����N\<v�Ʀ�o.�<�o��~;~��)�������Ա�'~�u�h��܉cl�/������5����?����x�����LiL��F⺛cAq/������ٌD��?r�|�=��-��>��"�"�KASE�w̉#0�Jb#�1Ӭ�o�
�%�Җ����ҹm����ٞ����_u�t���^��/�T!f=e	���(����:�g��ۍ�#��%�W�mS�x}�?�'|L���?m"�)�_�����]��5�U��\,x?��[V{. �SW���P���Ը4[2��XGPh��ȸ���qc��w�l�?�����9��\x�����imH+M�q�s�߸r��P1����l�ט����JEtl:}�];�g��U�����Ԩ0��1�Y�P�X���Z�Ӷlv;�jK��t+ŉz���_�ݣe����%w}�1��Zk�&����vC���-Қ�_�Zf � 6��,U��R����c���>�c��{�E���z$�O��cr:��r}����?4��1��a|���?CG�cl�n�4a��|-2�ʿ�2ʯg��l��w��+Ȣ��UR�)���OY"�mQ�eKQ=�K�2��	���ѓ�?8�31a`h��������V���N+��_7�o�����k��	|>��AX�#����-����!,��~�^%5�u�ﱗ,�`A�͉��0�g�|�B9no�"� e�$f�Th:PՇe���)1E��GыҔ��W<�Ҩ������{q��I���dd����J���-�/鞰,�]��{+^)i����
�~�oh\�A8j�
3�t�o��!��k��9s���{�hM����`=��� �+��Zcv߁IyC�p��jLk/�e}9�w��:�jK2�k�4��|�^��t�ľ\i������R���l�<aRC25�b[F^���+5�Mx��!�Y���A��#����UrQ�'#[��L����o��ևؼF�#�P̾�A����F�Ζ��D�E��\zS��#}����u�_3Ⱥ�j�-^I+��7��{ƻ���q_Q����5�lT���Ů�_����^ǡ�R�R �Q�-b����
O������1KWև��B)��:�PS*~i�_kgjs}%#��(����R�-�~7v�h��+��C�K��a���<�`�����2�`1��l�`��y��<�y�q�=�in��T������%}��Ev8x�7�O:-&��YIP��E�U6d�6�Qnl�H�m��V���ܽ;�3�����"�|�nz(�G0+�W�<�w�
�וY1���"��3�Ϝ��/��ԽX�h��/	6!�^i��wq%{X�7.uGlv��&�TM���@��q�E��jty,D|�2b��D[�����%\h3��p��R���u�eYآ�	�P��11�SZ��������W��my��� kW�SPN���Y�rzr��� �����
�䀚���t@������_��m�Ő�(l9]���1���m�i�.��!����V�'����i2�<�SR��&���ҭhG@#��uu)����e��/�g��}:v��P �6��W��t�:e��e)�5��Bs��p@k-YJ���4��/��Ӓ�)2�|՛��r5�LS���c͋�u��Zde,��*=PS�]�Ұ}�C�4�]񳷘���*�Ū�2�=+7�T<Xv�e�vp�&HX�3���//�%�k���3��'�q���<�����S�&�}�S��dm��/����!��-�|k(HkQ�٣��7�<�D�D�R��3���^�ƚ��W�&����Y�2q"̤�3�:���֮���ub������
�<��du��m^�_��g�˳Z�[;��xCf��c�b���{^{2�U=Ճصt�~%�ì�@
M|k���ge�y�}��
��>�r\o�Пږ�	l
T�O�h���.Z��f��6������JD�Wf�����D�򬬵��'є�n�0˒�^"����N�Z"����q��_��Hx�1�i������Ka����q����'���v2d�R >&�]�!1O�,�����{Q�&�P���n��у�G���Ac��#���D�Z��K������)M�ʳx����u�����Y+N��~�WFyҏ�@�!Hd��S,��J�hĖaB���.��~����X�4Qf'�)O2�{�,�v��>^al)-U�V}K�?�mk8Oor�nÏ�y������;����$ׅ�291ܹ�B�+�먡'�(�vAQ�2&��Tz��m�:N�K���Iթ�s��]�$)�v���c��I]��v����g�dҋ�S.�'����pD6��j-I���jM��kMs-��ዸ�x�h(��a ��;S�R����V,&/;0Q�3�O?D-�3..��2��_�J�h������h�?D���#wǥ6�'�y�@$�Z茢9�V�4.9���~"�m��N�ˈ��T���^�r`��=�/��;@�M�YE�����2���(�{�@��CV�n�[������`�ʩ��+����Gn.��P[W"]���`�2O��c{P�(g���P��֬�\�m�U��щ.������d|�����1���}\A��:�A�$OX�����;��JJ�U����Ph'�	F��;#J��a��6_L�����L����92^��tP���0��fTo7i�D�g^؇sh�{�����oϺ�<ƃ��֖$�}S7�m��6L������t�����Q�����k����S3ޑ�풅S�i8�v�
{PW!6W[�<{g�\��38���im?3�-q?����RE����N�Eӕo%G��9�>&D��o�kT\��
���l�.ӝ��K/�26��N��4�!�D�G�pKg���w�$2.�ǈ�w�8J�]��aA�A�e�����>����A9t	��aԯ�2]�4�� 2+s^Pw�m�2ELI���9�:�r�;�1���p�Q�X���!���z�M6��Cނ�a�!+�$�S]��>��ra�'����t@���Jb�nxRݨ�	&���E��jҡ\0�����V�+2S:��5����>�-3�d����	��~sm���{O�4���d��~�ۙh�l�� ��~�Ͼ�[���O~r�A����K�w��i8Q5�ϣl��q�v[]�{-#| pZV	~}�H^U�p��mт�m����߁�����g���tj`�� �è�z�[�y?a}�=�M6���1v*XX�&%;��Uko�b�j-ͻ�>�}p3+�1���(�iFW|�����l��~I��K��N�dY5T(:*Oz��vV�{r?�T>@�����,��/��<i5�[�`��a�hz�F���ل���-F��Z�-��e�����F	��I�J�PC����c�5K*��ﷇ��ې!�e�#ȉƉ�N��O�:��R�bI�(2�n6����Y���&Q4_�z�����yϱ�"��x*=Q�
N})W��-l���6���A� ���%t]Ѓ�yV�+���T1���)͍4��ϡ�c�Y[|qf<C
W�h/[�j����pOV0�U�:�R>/�IkGh�1�]-u��d�	M�.#����(�6ĭ�mb��a��Z6��^Gli��e勇�5轉��X�-@i'���~�li~��Q�J�Z�`��c^�[@�>T_�w�� �w�9��'�tk����&ۮFj�߻1>��v�s*�#�¾�Jq��u�W#c���v�����2������U�+bTR9������|�A+v���6H�캦�p++>�!�YY�gyi�a���}E(A�E�Dg���9j&�7��Ylt�X <c�kc�Ōr��J��@L��W�ւUR���rJ֛���-'z�)1�5}����1�EP�z�������:�ۢ��f�����Z2qR5�z0%��Cl2�_�e>���^eGq���y�:�>x�d�����M��Ӕ�}����ӦMvB�!�$o�Ӂ���_5�u�<Ɵ���A��2��zb����؍HSHԂ,��[��}LW��M��������ʵ�i�͙��w�X6m�Ց�U3��U'�����̽�W��ka�#�'D�-�+���C�|�k�I%1�O�<���#��a���.�J����f�r�"�)�CvJ�ſ�Z��XT���x�t�]��nN ���,�/��e�c��'�Ւ��M6o����i����>U{���%��%�؊��-zeQ:�Qt焌����y>=�*1��ҩ�&v�/��)����GK��{sΔ[�Ǖ��I���/�d�4�a�?���FJ�SF��=����,�2(eh���&a�aq#x�o���mN�@v�X5·��B��|{5�A��6G��r�s��b�N�m�P[���3�Y���mV7�$0/�#F�)�%UJt��j#�7���0z���D�G�����'����� ��=�QZ�:(���W){˗�_�ɦhy| �C�������b�"�Of�Gy����*��)\�}ǊI�$n[TgՔ4#�w�/�<�������&Āp����\�g�n���j��!���T���BɂԟL��x|֣��~����${wSYq.�4s����=p�&8�
R��k�_x
GS��0z^�k�*[{iI�GEL��K�C�V*h�喊���ݳ�rk���s*�C�8�]�P�'�E�c'^H+�G+Ou�.�?��# �wsr�IZ�e�,���a�GKiUJ�kv��C�8U�`��9��&���W��b��D� >~UYڟ���(�f���jUQ�#"m����P��j�i���t���m��]������6ѵ�����	�s-����ZA�����G����3���w�/�TD�F�����ؙ��Y&I��
9������>�ݿ��zu�Ua�Q;���������+��q�Nu����S�k���m1[�踰�Az�/�����w�����|q�N���Ao���t�r��� ���|+[e���ե`�E�>]6�0y��5ק���B�HY;̇֏���f��
*���noy��[��!�F�Wh`$ڹ�ga&6��A3�[��S�n3Hƚ2��Y�Re�-�:��e�-'L&z��7������n4S`�P���ڗ��CK-��i�Y.��L}�~[ߨ�T����O����f�P�#6����޹��me����lj�3�4O��d]�r�36�5A@E0�F�P|�v��6`�{9��,u�@՞�F��ټ��>�蔻S<J����ˢFՎ�|@��+#��WS7n!܋�!�kS�IuBMn�5|�݉Z=���h����Ru.u ������<�,����Y�I똛��,�YEȏ�U�f�b3&�g�_"���}BH���hz��|-:)�������'Վ"����{�e%�
�n�%=�8��=��ꅧ�^9����1�Zi�/ȕ�=�+E�*�o�O���f���^���O?S-8�X֚ ���nɫ)\�l�[��K	�#2^�6��X�h����������:j:�Gl� _�����e%+H74��Y�^t���2;׆e�HU���G=_��i���z�u��߀�A5���>P���6	��JK/�(~1���UjʣCE�6���g���[�E�j�Yr���������ݔ5!s�c�7(-Fe���W�v�-/M(�k0�i'�Sy���*�3} YTekC�d)8��:�
����$����C�Z�����C�u���橒��8��&_��N���S�?��u�@��u%ֳ^��QL�u'����:�YO�b����Ï[5�}��k����f��g��j���|gߠ\_]���������XS��\Tv�~i3A��}���MYUTV�����=�vKD�J�	�c]_8�s�������������L��l�������D�����K����1���쵏���c�7�tu/[X�7s���?��
��V斃O��A�
�����a�	����G+���ƒ��`���u�Cm�m�y+�v�:ng�]�J��a�|�Et����蒬�̟ۉ��-�1�\zx3�"W�����F�ǲ��_-����m��M�-!��p�A1��}��#�����4��Q��,T���.�Y�����w��������!��S�����O���Ͱ��f�t��U�s�jr/d�x2�[�Z��5�����r1��hK�EPiD�3��ɠ|�ʏΒ_�pU�a��SmC��b`_UW��^��Gl�ͺ���oK���L�'�RQɆm.>#R��
ok��P����H�C����'�H�T^=W�q2�$�ϳ�|#�i��#ZΜ�`���c�O$��F���x$�=q�k�
��G�TX�-o�&�/�X�,#����bj�t棬�P�#{���C���fV%�rXE*�ߘ�xW ���e<.d���x��@YT"N��N.���������pf˝&�[N#0���������<���WU��q�I1����35�+��(/��D��_y��<%}w.��,�%5/\A�vK���(��~56�a<\��\P6�h�!w>u]R2�םٳ��w}Vg�+G�$� ڨ��F�E읮��o����?���n�͛�ߢ>����z~�a��|1��D�*�I[o�%�6J�=r�[y�X�Z��ɞ���r�Oz�7�ì�žy���<�+�i�3�,�GE�X��Grߛ����P�����"1�y�e��d���X ;�|�}��ˡQ���0��D�N"��f��������l!�ߝ���|?*~�qѯ�=1����x���A[��$�i�H�oO�,���"�?�-�eAR�N=��Um��,���*~'�'�˙7��S3����3�|u즋'��S��c?���_lIK7M�?|��t*�S��{-����w|l^�	������?�$���3��!��[��MF��V1}��^_0���ۜ�D�����2eym���ˑ�Vk�v���Z���q�z��\(lDՠ$w���Ƞ����7f�R�;������4�E�<��I8pۭ�٘�	LTsbBA/���^��Ш�p��T^V��-,�.&7�k԰��5�о܃,��pax0��R���.e(�Ϻ��|r7x�Ң����tK������p?�=G~�u
)���띚���v�D���{.ه��,H.hB��y-Uq2���9������T�+���z~x�!��-��,D�͏�vz��1�Xddڈ�+@e;�	l'Gp7���s����rJb���6�� �w9DE��6��k�Kl�!/{��F�mM����o%�qͧL�>�-�͟��#�&��%,t�v���F�y��<��������%E�HU%���U)�9^�a�:jG�FAUƄ�S��8g�S�e�#�W������9�|�ڇTz���ԝsDJ���v�� ^eឌ"�2w���5��r�'fʢ�n��oQѹ��IM7���,�0_nn�dm�Cј��1���fĪ��$�~�>M98ŋ���4�-+d�3Ugr�5�w���F_�Ǘ�|�b�4�K���sz]
�����f�x��H�c6�[j.x]�M<�S뾣�U/�4��Z:
ڻ(�TmՍ�� ��1YO���+� �ґn%�4���(,TS�.��V��jP�|ň����|��ӡ^��x�kD<��)�#Nxc���K�TT$'�]X�u�_S���?.G]��� o��^u@?���}��$��?`�/����y���a�w���o��u{z�w�M��w,x��Y�N����Zk�R1��C\��E��[�ut��x�^��`����œ�7� ;9��V��B��Єv�������c��t-��?�-n������R��sұ)^��Q>^�yW�c>���p�M���8jp
>�;9�de�.��_���uT��Rld	��˦���,~JY6����3]���#��!<�ڔ?j#�<4}�2����;lW���4oՏDcI��缃�*y����s:/�����3�B�Hq��?H�,*�SJd"/.򴦸;���"D�2z�o������_�)��*�����0�`�t��	-6�倌X�n�j1��Ѭ���N����b�u-��5�?����ec�.��W ������Ӯ��ky���X�:=�\`n���|Tg����)2�2�U�x��:�x[��˶ڡ�M9b���[x��\�``�5$�(�L��׺M\ɢ��	�.���q������)؊��%Gv�S|���A�~���@癓�`��bH�%z~g䀪��4�@��L+B�X?a;�Ԙ��6��07�gf��Z}L���0Z�}a7�:�K��#%�i���.O�K,{J%'n�(:��x�����Mrb������x~;���3R���q"'�E�V�=�1NF%�!���Kځ2��/wMě�I�0-K$�@{��oA��9���p�)�Gu�Ԍ��:O˲�=���-�6+/�����g�w��Y�)��l�����pAI�jJ�}��N��;��M�\��_�ۺ�(��0~c��^�e���T�L��i���9}���`��i��q������)�܉��$����� �+N0����竞�k:��e���]"6C3���2[w����w]Œ ��X lڀO|~*1�����`�/�Q]R�"�w�􈍔��S���l�5�>Ժԛqo�J�����Y6��?���Y���ꎿł��*����&͖ޗi�(���]�S������ܯT𫐉���t��׽D=�?�|����5F[��M(��F�%��;����{���(�W]��5�FF�5���,�W���H3K����6���L�P��շ�iLg#}�*O�g���ک�a�|��b��n�X�_9A=�2��HU�{6�GD��7ߙ�-bK�~��[=��G�J-�Цv[g�7��&�_�\�Y.gt���A�A ���T�D��<���Tٮm ܽ��O�{٧�V�
�>��xERZ�#�1���z����Uܡ1�����9�[V�o��z���1�#�B�����\o�w��g��a���SF�Ĩ1�Oc�&����-j>�fg�S������}Q��7мN��[���R�`r���q,�W��R^��
,�����]U�!���|�Kfĸ���4�&r����n�oG>5���<	�^k.��\g��{�,�V7���jm��O��?Xd{_q2�+���T����iτ�n���.�E�0g��[�$���K��ܗJDJ��]Te1q��}���D��(��l�TIтG7�������TC�y�s�����H1�=�`lc���D��-�ek��U�OM=����6��)�*��P.�$��<�������t���+p��)��|LPee*�1��>V�s�S^5Y��ܛ�-�/��1� `I��tu����hsb�>����8�����fHH���"_�ub���aM��f/�|�QcnD�%��2^騪��^�����(vꍟ��g7�S��q�E?!���g�������6�C���}x,قFv���!��Q�8Zz<1���U`����#�Um��1��q��)؏-�{���N�˘	�!��pJ朴˄����\z�e�^M�عSށ{~��伄�%�l�b:|ۧi#� y}U���lD��S=bKm�S�$ ����洺0J�t-�K�h��[�o�~�x���3���h/b�w��6鯹e�"!��VXI�ڎ���N5��BK�NW8�Jǖɤ_璏������$2��W��`'bX��ܦ�0��F�a��L8�r�]�h��Z�)|���}���O��S�q�L`��ww��sx�.0��@��94b��N��A��������F�	JH�'�e̼�[��J���`�������J�<�G��^E c�2��|�s�.�a��]�#��d��욟��`N��0�C���j7���oi�`��!\��iJ��;_F�E�ڨU�v�o�9��*��*v�E����|���bM�c���~h ";5��i���W�,�߽XH7�5��ڗB����@�[i�VΟ^C.��k0q�h�U��������f��}Rݑ��X�<�W�����ه�i+�Iv�JJ�mf���[��C���>���}=��?�W�V��y`cp��� ���#�(nhz���h�L�;\)�U��0��4�*�\�"�2B�t�y$��,:�mL?���8�G!۸[|e�=��n��/�T��C죠vO�c)�nJ� ���5f��)\<d�DV#��3j��+�}ZT��JCD�'�kڭ�$�Q>xMh2�N�z�3y���Ѱy�%�X��B}5G��5Px�RR�\0�����,� k=��xUN�O��`c�FZ=��{P|��o��4u]stE����=���vg��^�� o�&�Y�c�y<� ���ݶ����%0Ry+[tW��q�����b"�1IM��dTc@?��xb��������7���9"zuH�K�T�*
q�ઝx�������K��"o�!g2��NF�5jD��ۻ�j@�ھ�9����@���9��+4�vM�+��kqiT�U��z���)�=m��e[��h��Ra_9����/�zn�����Y� 2}��~�]�)G�}�X�@�9�:c޲���7ËN�O�7��ߧ�7��[T��%��a�������^��͕�Z�g�q��[e���B>���:�Enm��\�,�FL?��V���ߤ�M/�����dmI�9�����-*�h��
����J���!��0�D�pï��h<;ٹ�������U�d�8x�#"v=�Vsg�5�޴�޷�c�
��2]j�K�;~�V�S ��dx����=ܜ����r=l���2j�`U+�+U
t&���U���;���\�A[Q�F����-�pe���K�M8Sӕ����[!p{99M4�/���g=O����E��A�����֍%�	�`1��
��~9�ͫΊ�޹+�؁>����G�i�/1Y�e�ѱ��-	�ਸ�6��H��Q��]K;���o����Z����Y����_d�r��f�s��W��=��@n���$���rWL��rYd���ͷSל�.V�O��?�8�5{���*u.�ze��@�����L#*S�X��? �c{�s�m���B�*�֋�{9���կPV�h:���ڌa=Ƙ�K���b	���7��	�����A"�j��z{�9H7K�����Y
��*ɂ�|�>��V�Ͳ��OH^MA3�<j��-xp��!�Dak����Aa�8��%j��pD��v6W�~��H��y��i%����,tU<v�F��e���OZj��L>,��r(��Z��]Vԁh�fѝw�b�*����=�"��ĳh,)x
CRzn}��|v�+y-"�����%��,�3��%w6q���|�l�h�E]�O*�����)�^�Y�V^p	+Џ��/�k�98=����I�!U)u�"`K�d��M%N!���%�����G�/u-,�7��>Q�M�����^�m��e�*�QC)�w��*����_�Ԥ��>����AV�������>�!A^��]�g蛮u��������*�ϥ��J-�P�L[���3�_*'V/�k�l�=y:{�~�աjj��eR��5�\���%��)<�2␅$E4�CQ�-�@��#tX
x{(z{ǶyĦ�d��kt�M&�7���V\ի9��dݕ&`̉a��.�Ϣ���^c!0��&�ҺJꦾ�L���iPY{�U9��Y2�j-����yɌ'�7�#BL'|����u:�P|�ծ�Y�>�)*9Ň��qPS��w�����p��}��ۧ6�����'时��WΊ��;�z沪˪B�5�Kʮ'!�)��FA�	wy�	w4�Ĺ����c����#?���%��I(TA~�߈��f��R9	[qa���� pQ$�+�hI���0��Ç�f�y�Υ���Z`i7�����Ċ�����FK8�եj�H'��5�JQ����������h��Ё��ȶ���� נ�~pH�z�1��2I7�r���\�5����,���6m�s�&�C"�6�_��n�x��z()X]�3c�$��
$l������IG�b�����N̳�ز!`O��3�r����`�����u/�q�f��X��%�~�|�ur�>z�,F���{/�u�j��9on���B^~��~��oɈ��+k�>��EQ��L�b �q�c7r��:���Pf���J$�Ϟ����y,3*3x���|�~�zܫ���?�\�~ȝ��I}�i���N\9�0�)�sm荈�C�Za0O�cD���7Xl�o[Zs�exi�"��/-}��b�$w�ԆMJO���;#�&���zBLT���(��{��1|�ʌ#��χ<^N�����^�3����A�c�q,�'���\3�I���'U�犙�u�k6�_lL>��)�D���<���;q��]���#agĺ��^C��C�Y }A����2��.	�&����R�9-0[�z�1������+UgoS��c^���j�$��2���J8�y�d%mj�଑xUF�ŝ�0>� U�>csC1��_a�:;���⩧����`2�|�C(��驴��1灕���I)<.Lӄ�:�fL2�՟��	��9��{�wPf�z�&��a|ؤ��G'��-�����P���U��֭,�&�]]QK����ۏ���dKQ�gn���Y�:�kl���զD���H�]��y�Yَ7�l�{Ó|�X�G"�Xc\�T,ر�����ȶ��SEbĮ��8������~��/����ǲ����)A�۳���V���]���>��A�������M"�{ktQ,]thǽ��'�Q��}�ҿ����o�h��%��E+�p�s�})X�Ԏ�J��s�P�g�cȏ'����$IG����&�V���<y��
�?�г�؂o�n}E�6A:���@��./�T"xYe��3ٛ��@BD���?S��4�=�Y�\�*�u��87�E\��d:�zT�o?]�Z��d�l�zY���4�B����űڕ�}��FR�Z�d��~5���}������_O$��0q��c�?6�B�eq��.~zK!��v$�x����;��y���,,�`�@�E]~bjm�������RI����O�^�M?�K\����Ҩ11�L�)���rb���\W���E���'µ����&�~b|yTjQ7�JY/`D��SI_��%W�լ�޾�j��y�F��l����{�1u@X���J�inM���jm��eV�1�A�<��=�U�\�;���~vR��K.j�5�\��-/��6��{��v5��m�b�D����P]�h������N��pX>g�Źd��^����]]����D�9��6���ŭ&��BV���qogr��)�2E4�}a!��9ֽO��*�&�v�O�#���FV(��
�����`)����&ᐩrul�V�pR����@��^���f�zZi��ʬh�t�`+V4CxW�]=��+]N�+3���/%3!Q���y�a���p������?���J�V{�(���നϴ���Zv��K7�T;e6w�q�ߢ����1 BQg��C��c�-ZС`�a���Om�}��+ҷ~7�9PM`��<�;����%s�0p���9�1?�9���Eb��1:��Y3�!��t�����[LߤyxR��p�!�H9�;�W���ͥ����x�WMzݴ��< 3���\��ďю}�XAp'����m���\�y~R��c]�O=os��o���x#OV�s����) 4eȏ��u>�_��ilfp�U_>!w[ꦶ������u�P�z`P��#*�|�3A�f�k�21喌���.�O���#�!�b~�	N��G��-@;Z�k ��k��m|+�r�Ũk��m�%���r��i�������w�v��1q��k�͔32��/�W��������~�+�߮V=�mN��jkߢNn��o�;��?�'�e��C��p?@@�^]f�uRCM�� \�a�疃Uu}�P:�^��_��ͩHդ�ꐽ1�#���'�dټ�
'n�|�[��r��V��y�7eR<<ᲈN��abZ�*.�zX)���4R����ՋK�W�2LmKΕo$��-5�s)��W9J�&]|�>αZQЎ�%�ĮF'9�Y��$��<�rXw>u���v\�֪��M��f�M�Q��p�VFv*et?�\Ji�^�����.�pc��_ۭ�3�����o��>�J��F&7%�{���@�V���m�䕜�7�ΞD7ˡ���Q�y�_]o�^�X��y:�UŦ�y�ܣ�j�=�{�8W��kT���/�]�eX��S�C��,���������tg����40�/č[�d'yubb�/_ߑ���}5�K�9Tߖ�iKE��i���K�6���P���}M��#6�U|��0k�1�g��:ګMCd;������5��qn���0�w��~���4�N�)��=)w?�x#�x���A�O�GD�oEc����;�vN���R8���̑�}�������e0go~6�L�L"��)gV�a�t��~��.5�`��.�5�ljQ5T�d]c��%�ll�'G��P�P�L3�ҋj�9b�6���,�1vST������z柑ɫ�V׼��in��	v,��o]�X�w���{��3h	�[4�v�Y�М��:J����'F���&~�Օ?f��N���l�
}�j��WE`Ԑ���_���ll����O�X�'@{A����ViZ��� /��,`��5�������)�M۱�WOݲ�CSw�bO��݁�;C6 ��ɑ�����.���3й,Î���B+�'&)�R�;Nhcƞ}��O�S�1������t�i8�������1�{[�������b�U-7�����,'G���o7 H�(��ղa�ڗ�SU~Z�������d�n�=����� �����:���`����`�첃w�a��w��	:��U�,�٩c,��#����2r����-$T���t!Jz�Xnm�ܮ�2��ը����O��ȧ�t�Ѵ��x:���-�B�ٜ�1Q��bއ�B���C�`�ܼ�����h	3��<�[�'�R���־�����9e��Ǽ8<�������x��#$g1�ȿk������A_3׮�� ���ԫA�$�V�M`�4f�ؔ��K��v}q�0���1�1�8b� %��l�=�{.��U%/BlzGQ�N��>-�J�6ݚ�a���>U���-)k����ӵ4~��7A��Ot��7e���FK�@��	��ּ�?��p�Y��Oֵ���}:!���!�
@{!L+�t��Cs/8ky���4/ޙ��Eizڃ0M�YT���S��W�	�.���:�������Hq2�'�{��b��jB��S���i/���4!>�=W�s�߀�~[Z�B�yv0��(VU[A�̍yz��;zP3|'B6Wvl�o�ه@)��Q�?��q�[�ɸ�s����jJ�[Ï��j@�dU�ډ'��v3�ʓ:�˞�4t�n~x��7x��rp�8���Xc��xQ���v���!��t0PxY��M��CBtC!��ͫ���������9���r��%�����F����Ƅ��B4�B��A�C�_,��3��`��>�=���tt >�s���)윈�R��AJ��0��[�}����,�輞��ڋn��{��6
�&~���Q�%��x��U^�&0��b@�'����w�86TS9$b��;�S��i���^�2k��h)�|�$�m]� þ7ʯ��&�ء����]�v�k�On�1��Ebȍ_�f�
�[�����?�V��{�"��Q�~FAt?H����E$+��"�s֬�m�Y���ۄ��k)�- !V�h�z�� �0c�g!_Ӵ�����̓2���)��O�	���5��'��%�F�.�w�N��x�M�{�1h+�_;m�� ����0R���gx�&��p����o�Kw}���}2�e�F"C���쳲֮h��** 2����2:��õ����@�K����߬r���j.j��k��/��?-#Q��hm�����f�3�2:z��)��Tׅ�"Mz�&��$����E��(E�.!�PBIB��D_iBPDz(*BBQQ@@���3ƹ���}��Xc���5�Sn�k�������/��)��˟W)���9Q��U������ ����w޵ I�뙙�T��w�
�l��	��xy��:���!�9&F&FfFF���"��������eucA�kP��ޑ�B&QW`¦�p�����������s��?,'����o��]~�gu!e9�"hT����U�H��������(�N����Ԩ9ټ���*��מ6N�O���s�������-{W�K���!��x9���b�:C.�;�=1������\��	l���� Z��j���9p���Η�d��u��Np�҈�O����XAu�R[;�βuH��NJ����^yi�]Y��m*T�\C<�O-�rK�o���m�L��ϲ�~�'�YS�񲾽n��Ŗ��>��Q��sϢG��>��3��^�_��_�3>��y	�G}D{�˅�~	�ƍع�{Xö뾾�K��/v�7�.��>ro�����U6�//r��_z�d�+跞�����럫?ۈ!C	`獪���ੲ$--Y���ru�	��1�r>e��\��lj�`O�ט�Z�w�N}��c r�`���j��+])?��4�T�~����\�&�F��8F�Q������ͧ�$�g��-8����D|0�R��~6<�\(�,)?�)+�>�rM^���zjC7�`�s�:�i�h�_:Ǌ�i��"s6����gs�kX�<Ua7�f����h��ø�i��r�{m�ne$�2���؞�ٲ���tHSbQ�	��R�:w!y��h��㮳���;-Օ�l/<m^zp����G�#O�TFސ�E�
y�Ð8���J��pE/;��@kj�]����.fO S��+b�慇�\u�LW�=���U��m&�sH������. ��Pw�[<	~5���s�P��.沁���G߼�6����Rd��Q�W�����=����T�-ƴ%�1(w��b�)��qitR%�?[�8��:h�HB�a�y9�pߛ�Wnk�;�{����ʭ^���+��9O� fz��i���7$~Y"���-a
h�L>��~������
S���Ã7�|�?���F[�Tl�۰�.�o�.���:Ś��!F|��dϜl@�k�����!uB���d�'�#�ȑ�sd�ׯ�[�T�:IcĖ�����% ��ϐ��~6���� ��/M�n�w��9�}��5߾���?M��h��O�e��+\M���3�vd�+j�ս���4Kd�~�$�ЌЪ�Dm!��,�5ER�9m�
|�k�譊(�9�k-���4YY<��׮X�7���@?  � C�Y
Y
y� nt��ݛq[�MN�
��*�{.�Fs��~!���i|V�cx^A�rǬ��؏�C'��m�K%Le4.sH�=׀C�%2
_	���zc�e��8^I	G_s}I�-����3�Hi�D� ���o �t%F�uB��ݎP��Cgt�Z}��h\G3~�L�E�Z�aD~���ǹ��̳3�^�p�@4�< n��[���m��d:�㱿�U0Oj�"�k��������z�����G���O�����t��_� ���_laҬ�7ZA"�{u�%Oo��<�.aq��;։8��7���䃻��"��B�/Q��g��w���r�i��n#�	˪�Je���Gمq��z�N�$��棇�};�K����m�����1���D<�Mc�_5�rl�!�2�2
YP
I�;�W���o�o3�{�g�k>7�{�B���\\�S�ݞ�%Y�6�N��Fw ��� ��Y��d`�$����{B��O!� O�� ܭ��ԸY���ݣ�[6-ĩ�R{L���Е>���("�@3��a�\[=����|y��i;��)Ys:�9�&;+�d�b(�2O��A�>�!�`b+����Ͳ̏�Q%�"WU��eB��ڱ�`�g{�EH�]Cv��d���������/F��2�W����]c�Q�
g�ӥa)
>b����v����I9�?��E�����x7�FF� �M��M�P,�l����Z|����}���m��kҚ<�믰�o8�}��<^��ZҀ~��c�:�8�`�NL��0�iT����\r~ƱO(��	k�~e��r�ɺ3�6y�����o_C�3��&18���e�����Pj��} ^Z�"ߢ�-����{p01�gUs�LyVc�~KH�� ��SM	�9��C�u+����+K�fY�Z�]P'��P���`�E�*1>�3�l�E4+^wH�a�����Pk�2��Z��T�5�S=�Nm�s�ɵ��Ga\���{>����9~��+��z��@�b����R�\w���(��^s�YS�]nS��=	����$8�O� t��O�_9��M��e�˖�}���f'G�{��'��$={�2א�vtnHn5�V-;�w�Bv�5��I9�a��k�򉸐�b��3~%AB�X�z�� �
�c�@��Wx��M��6��)���x�z��B)�ـ"���Hx�EkU�/���^A��C�j&-���X��$h���[aDu���,��M�� �l�����N[�*4�0�+S���O#�o�#;\8����\m˪����{\<�{Y�W�����׹���1�nF�	٘�q��e����`�~-��o��P{�D��U kP��3[�7�g�U�Nz�Y+�,�w6׉N?m؍�^5J��f����Pq�-��J�n��.֬�f�;k)�o�kQ|L�������=.;��E6(�����0�e�]U�	9tA�YQ`ڵ-���1�Y���ҡʶ���b���Ǖp%=Ju{����h/Bd���
�Z��xLΏ�wI���=e�0�DfM�b0m������b�NrmbC�/<��8�<�S�iV��K�9zė�ekqhT���:6�g��h˅�i��9<wi��ײE9%����6{b?T��Y}�+�+�q�ԁ������{W,%f�1�J�yt�bDm!��E�w �,(�==;�?P��!`��_xpCbH6�o���x��&��v:�4�d�~l�]���X�a$���Ih�3��Fd��C̃���vUY�ދ����p�t��^�m������uf��5�s���`ZZ�,̠��l�[�d�n'�	�a��7��� ��֭�mYQ��J���A���o}?*�	��dIdqM���c��(d���1���C|��,b�rT߂��Ҵ7�-)ګE?^��s�p��p2h�3�
����G(��_/��S�1�=cp�]X��s�E,2�~,�QK)�F�ݘ�V��d�Q	D�[, S��<�.Q�Ǿ��X!|��6 ����D�Jj\8\�L�N�JP��z�T���4�_omV��4�%��]�V�.���Z^�I7�{�N	�Oz��u�Lc�0n^�L�le�'T�ɧ����
R�xc��?z�h֟ (�`�҅�Aj�aU8����V���,a3Y /���] �#�uYۤ�l}^�N�Z�d�B��v�z��V0)ȵM�D�awHcv�7��3��B|T��J���R�ĕ\���*4���ۅ��>-��ˀ,[E�(fw�a�o��1J�ըX��'�m"͙i��ʝ�~�����=�P<�̫Vp8��nŦd�� Ʈ&--x#?'���N�9W[{������*㺇&�^�x� �j��w���ݫd�.��g1�c�ƣ�i�2�L7g#��_��|a��=�$GB�ۦ��̫�U�n�F��Ҵ����x�;�c���A�^xh5�*���4/5l*���i�� �����:��4G�h�%�c�N�ະ8V�8A��I�W��,(�끥�I��E�=�l�T�5b[�n8����������עA�4�԰�ic1=���ڜĞ'q� #c�j[��{ot�6�5a��?��	b�M�o�����WPB�֮-��Ę��GP�Q� ���_�x�wy�̓��h[�������캏�"�pq��������)�͍B�`�C_c4ޤ�`�RZX�S8��i7���AÅ�K��Ѯʴ�K򨲫�����	�õPl���1Z�~���5cX�����3�'6U��H^l���s��5`�� ��?C��[��T@�;G [p�BK��-B�@/��HL�C��_���Jp��J7Дo���^ ���͟��^ ЮF�_����Ԡ��V��\tT-� ����֒y���|���~Q�ߌX�Bj��kH��b�
�����_��/*2��L�p��@LA}��\x��2���ᢿ�9e����7>զy�T~^������<ª:�܏&����5:�	#����T��|E x�r�\��A�/�}�	���3��@;�Qb�W�>kX ۙ5T��dd�8;�l��}�x�g]Ʌ�қ��Xms8�^n)K�y|��s��B��ޮ��O���S<�_�N�������/Q"_�x��OC{W%0�y��Л;P�T�8z�Lg:m^���Y��n �3�Z�e� �?�'<����`E��݌�L�
S|cUr��1OM}�ѹy���|(����J솚�Ǒ�@�lܯ��m�ܜ�L=��_��՜�j��!)����,UaU����+Cz��w0��!��r�Ó���!����'��ͽ3��b�~�Q߶�'�Iu�E6h`d�H#��h�;�20+�`@orى`�z�*�:�k�(�X�y��Xtl���nc0Y'T��$O���,b�¹��"uF�7��O?�qO�o)^3o�"�a]��$��{��Q�y�u�HfEo�U/��������ʸ[v�_�{�{OBC�>��{�V�3���5���\�.�D2VQ�ﵼ��W��d�->��8�'Ҁ���mp5C8~���*��R� ����2�T	���kb?}��9B�A�-��/���<�¿��Ǥ~�(��x	�)�Ë�9�2��s~�׸�q��x��MG�!&����w؇�Y�'���:�` �� pĲ�g��h֔�]�`�0ۈ
 ����v�d�Id�C�`/���%%>Q��F�b��O
j��[�����#��}�=^���W�f�:+���d.mua�����������)�=����̗��ȮF�n|�9/��TWv�]�[
�[rKι苷sS�,�d?�"�i�$���G��Ad�ڢ�`�Pg�6އEbr�������!|��K���g��{9W9�)��6-�q�s��S�,G����h)���uG}R�p^�]� �8�������||�%�шi�!EJH�'.�6*A�e�1��Of�C�Py��������ƞ`�"���Zvaّ�?ߛ^�Ei�[>�_�CskAI�RuS&�B�xFB�:��a��x�g�N/��Tj��x��O�0��X�i��Ĝ�J{`�{E�[E8�N"o����,�,\��IT�r�gU`�l���sM"�4���xī��G���]d��}*@�LP�I�ߘ@���X*9|e���s�D<jԿww�Rl�f(nQH��I��wm�O��G���S����A��1�xe�ψ�o�)5��v��=!�3�UD�б� �j��nَD��r��z)k�N��N�6L+m�%�g��D�]/A�|�9-5wV�E�s��1�4��2)�0@���I��V]�}�n��m��)=�8���Ш޸@eL�{ez��5f���u;BZ�X��+�P��Os[���ӽ�"�_s:J*«�˄�'u������My���|u4ď�/���?eg~�╃��'����7�Z?��iƤ�5l��HIU���m�k�p�Q��mes��~u9�w�RA���_/+��r"��y�t�'�l��1�l��	W�����Qym.t��!��d��J�e?��S�GGX9����[hk�����J���L��	���}��$2h�B4{������_�t��ڷ&0�����*1m�@ŵǔ'��:(C��QK<�KQ!"��+3����ԧ��2�r�+����W)7k�ݨDk���D�+!��ϱ��k�N.ES����;���0N �/ʖc���ưǏ2�͢�2�e��Ch,�Hw��6�
T�x�[�װ� �G�����yX����⷇T\�/\e�o��{`M�I6������E~a�O2Sl8�z�X/MzA9����
��s�c�]�;m]7B����+��Z��l�������'�����}�W�c��*bƙj��-໷��g���Ы�����<,�K޺�ZR��)�j���C�Ga׺�`+���#Ȋ��m�Th���;�f�r�g�9�X#.���l �{d�%+|��S�#��*�(����������s;�`�8�au/�1��A��;����|d�`nA����T�������yj_j��|C�Q�T� �՛T<n@\i'�i)��UZ�/Cdex����*����nmh����Y�R2Yp���>�{����94&>!�����ϻ��3�}��&Q=!$FH��z�x��o���RRڴ�.Kn�	���r�K(���Z�iQ��3��^�j-�=��j�~�b�!����=HI��8��8`~l���&�U�Q�RF]�K��\��,��ӇX,i���k�����wH�W���up�yr\ `p����b���������Zp�$�_n]F��˝[Ƅ��_��2�t]�|[+t�b�0~=;�>]��MQ9������T��>�$#4�Ky8���
��x)U�z���mna�X�M���]�дPl��r�P7�T��x���^�/[���>o�: ����c^��Y�Ѣ?�������k�ד�t|� �8����Wz���wDམp�!C>���ol�QR�^r�?e�,P@����I1��8"�a�Fa��q1��R˅��MK��;�
�a�)҃6������zLygF�M�d~�wk����ؽ+I��D}�=��*��=b�u����"$��;8|S�����S��<L�$]đ��6M�Ŏ)+		��*;����~ȣ��"��J���܏v6����J�
I)ދ����o|q��J�T��r?4���1�H6�|bsˉt6;ωA#'wD���Or���9�	T�1pASV��%b�)�j1�����p.X5wF��.{��v]{����f�عuA��<���<0xl�7(��q�=�ڱ9�ɤ����� �.;W^�*��/��������?/�w��Qu�@ޱ+���k�t���B�?\^�Ή6M��ʈ��c�o��߰����Dպ��%jT��k_�@gve�9w�ͽGsT�D���j?�L� ���Oڴ���Aڟv�&��?8�W
�� �)�߯�Gw�z�`{�i�h-r[�)hִt�����+6�	aJ��z�Ȓ�o�c����c���
�����iמ��2i1��H� �[R�四h)(d@!��HyE�/6�7|�|�	�n��RW`P�TU8!$o)��7�b��4]��[ۋ�z!#V1��?�ô��9�̡<w\�k�>_?��[0�@=d��;Ͽ��_��+�����X�R���J�F��}��wє���\���s�N��4#?UK��K�?C�}/x�?fq�[���fC�P50:��\����
9Āi�_,��*�w���l�$4" ��Wa1����C����T��N���h!�%?F�o����nX2��lԑΤ�����~,���d���9`kTÈW'<��t�/�N�/ѻ�X������
��b���D�~�����n]<O��D�l�wEd�<�Z�����y]�Ah�=�	A�8 �G��&M�]*����	Y�;��o�u�?�$��I{}~�F�(�Vc�;}*��&�y��h�'��u��ђ,YNG��r'J���k��M'���_�=��kn���D(&L�mʩ�t6���1�9��[L4�gV�׷�>W���1zՖ�SzpV��wG�p�9��ӑBt�.X�H)��~N���Y�x"��ׅR��� ?�W�W�M To���>�լ��0�����9�s�;���l��G�-�ˆ$���i�J�0�_��`z��Ѧ����E�	��k�����u��q�*�q�W0?\"��`E�G��|�y�$_[�f?��z�^ӏ�y���G,�+I�k�&|U��9y{�d[����p��@�8}� �Ez��WP������/��F-�ح+fd��O^�~�Y$~ǘ=.��Q��|��q�6ۊ���R�w1�;�B~�����(��D�<nY��Ʊ�Oc'��I���t���ݦ@r�u�t�q��;7V�%ݺ�*�x��5N���Ye�^<g�N�X<_��"7�~�b�|��Æ��w{�h&_�ᨪbOc���l��\�`���Ѯ�A)M�*��e�����J�4������j���p0T;��G%\�E��������U�|��N�H�W���9�UK��tuٮ�F�u�)g���>F�>��q�=�)����_�r�Խ�:�]ԭ�Y��f������%�!<�l��{_�bWT�c�T���F˩*��<B�~D�!�E�V��0@���>Y�$|4�]���l����ۄ1 �ۋo:�^�e�/̈�q��Ӂfp�6Dɢ��i���#��j��\�/}:���؈�_�� ��;��Y��]`և���9U�w8�W���
�+���,�h��(!�\y �r�R�m2��y��i����BO��h�6"�_G���YJ��OF�������g A8��x2g�?�۷�BL(��n�>��L��E�0��� �E�cj��h>�j~xh�g�x���n����ܒݤ���
qE�g~�N"x({?�S�>�^��&�/OלXX*b�&�h���,�5���l*�B#36<;�O0�����c�݄�(��+'��'�.��d�f��Z��#Q�WH��Q��Gy'�-k�����SZ9��m5��>k������_FN��I�j�i�/k���F�m-Մ��P)��<&X�^s���տ���9y�������<7i�w����D�1���=tK$P���:����1տ���ŪUNd��
K��Gg*�G������JY��纀��� �l��V]��A�j��;| �`�=��:\V����H=۩7r�Uz��f���� M��Ȁ,ׅ,�d1�����7r������۽xq��1G�u�����L/��z��Z�a�o&G�Me�H��[����D�#es��t���Q}8띟7xa�6¦�Qm�p �z����;�`���P�OA7�W|�n("]>�E逆ׅ�Gi��/�T`J�}Ϧ�
�<G�	KU�,m9���Y�;Wr-;WR��S���D�\ci�@�H�Þ4+�Y�� ��X�A�C�ƕ �w���	�E�1�K���:hE񰤩O3u
3(��䦵�EUQ&M,�0�X>�iKP��@��e������D]cq�.�vvg5Ћ$�Kq���L,&�����{w��hI.��+�Y���C�1"�а��GʕXmS�<�����A �L�F~�P���7�D�g�R�d��_����1�62�E��F�
�Z��"�G�3Ul�#�-[_�FT��Nsbn��\o��2��U:����|����a�\��=���/u4���͵��.���]�x�V���?S���ݤA�B�$y���	J_�i#�0Ⱥp!KN�)�S���/C�~����p�;�q�Ű�ո`�NYx݊�-�w����^��9��s4��t�4��-�࠿l
nyJ�D��N�?�'&-�U	�!<��Q�'�c��x�WR�c�����co�=Ń�ю�~����R�����׍NZK���$��/�RF��?���Ā���-Q�ݽV5�@	TwA�m� �Lم\Kf8�j*v�4�O6�i��v+��1�&c��0��=�l�-�4�0�4�Agh�U��	����-06T/�3U���VI���Z�
G��,eZ�kfj������ѣ��/L��b֐y�T�Z̺�k�-o�"��Jc��� �]��ʊh�Ӟ��z�Z,u��S_����#��U�����k��m�`s��;�'��H�y�{��I�kO(8`G�cR����j�=��olV�DdT�������dVC��POk��0��Ռl�ҟ��=a���e#��3��JL����7�{��>2����e��S�K���������U�S��~��
�:�-O'��LT�1F/B4�e���z.�şo@�#��ee����`�hH(ҙ�g`/�*\] @�"���i�{�G���Xx	;ly|�Blǽ�*?�3���ZL���`q�����u%�G�Q��i�/������`�|l��f�Z��i����\.M-͑�
qE1�8�ND��uo��|S�M 0��\��-��TA)F�W��~�	�_�e1[����˿BxQ
x\�7�
��$��` r,;�A��h���v�j�5��V~F"��^�㈸@�/���b5�y|�f�$R����|�+X%��$ܛ�Ҏp!?�9����Eγ�K�>|�S�\�)p[���li\���׿C��[f́h�)�R�'���-����	�QH��"�zno���K��$������㤟"����"�WW���5vK>+�d�q�pE���v���W��sU�Ċ�B�<�xeM��(�� ķb��+�D@��3bj`�u"����Oz?������]��e[_xh�Ά�y[�x��V��%<���􋅰�z�bfO%��¹�/@�M���1�$�`ÇѦ�"�!Z�c�3ˆ��X�&��;ěB��l[&�\}<g祦��֜��;*nXjB��z�BbfȨ��\ͷ�j�J�Bfz'm�;�/��M�Bf��=F���[��������`��k_9�����/���x���������/�����cQ�T���C��os�B��O �P�=r9S�)~Y\5�b��e�����4�Q�8ҚIᕃ�z)��y{�_4��@��b�_p�U#�ȩf�?wq����n�s��$R�ck)��V��>l�|�^����m�����b �_�����ʢ��7��Pد����S_�"��d�n���b�ui˝�U���*�v+Y�^�l�ZD����hM����/U`Ij�$[U
�15���僶qZB�vO�}�5�eV	 '\S�+&ÿ4"���t��u�����M&�=�?Э�TnF�^sv���K�]�d�9*-X�I)�h��d������p�a�����Z���E1���b��8[F�(�F�r?���,���F�	�fڰ���8�c�/Jqxe"�
�1:}��3���nh�1�����n��	�Cne�"l9ee����c����T��.��e���pz�Sy�
ߐ��fP��V�Ⱦ�6��X!��j2v�2�C��P�+R�ԫ
�׋?=���4���-�x2��u��%7�=@h.�n���8�z��d$��lJ���e�8�!O�B�=�}b��>�V��o�*u�aЕ�I_�V�E�s���ϖvp73�IЂX�l���4���A@����72�`qb�J�(���u��>��{�dM'R��K Z4�Tg:Bk{`Z.�E��f���/w����tC�u�GW�t<�ex� Q��V�9V���j
�+$=�/ٯ��h�,�k*m�9��Υ����{f��2��<����%���AY�ڔ�3�-����St݅��Ֆ��)q�.���e�F�+F���׌vYT��_W�8�Sk��G}(I=`;-(�/�+��v���:U]�����D�T�q1-�����6��"���M�/?Ap#��)!�zu]��
r����Gr����)���'V��l�ؼ�ɭ85Aק��f������r����!H�ez��l���O�ζ�F|+���	,��@k"3�]4�bf�r�ȱ�o��R3�90�~��ɼ1�Tj��O�gR��Q��*���|6��1q�l��a.a�W (!X��f|c��H�ѹt~Nt����U%�*��sH�+�Su�L��D���u��������*���kuA}	+kW��*0�3�v''�A�����&�<P�5a�J�	LI<�ɻ����i�-)�|"�o^=^G�F�Q�{,��0�����`!,Y�����|
87�'o�Pp7[M�8+�F,�F���:(!�X�)�l���BZ�����yK��۩�͸��a�K\��֯��E�lp��s�Б�t������1��;�+�BR<xJ�˒ќ儔� =8��饷o
�iY��BƋ-��T��ˎL�=�o��R)�e�>L���$.��!.Pr��{��&�q�E6V�<�䲷��fg\jz�UoR�f��QA�#&�N|�O�n.(LcH�:f
���� [.�9��V��P3���y�ß��Ӯ�fzL"I��oXVX��7LJj�\�f�΄���jVw�.�IH_в��	!P��>�o��nd�D��r�xS-w*Ы�ϝ���.��n;��3�G:�0<
������������2z)��V����2<T�ӈ�5o��"`�����'xϓn�O
�Yעg���.Ӡ8j T~bR8���b�]ϟ�j��XG��X����C���.V���,)�ӛ�xuV����2��UF/��a��-��7d�VEV��j$����w����DV�L"��-�iqՏ�k����[w�cX��R����*�SoٌV4G� ��s�73I��i�{j���+�<C�/~���O�h8)q���Q6's�rW�[;�zu�է#��D�5��.hX��E�w�1�9�0�银����q���#�'�9~�N��@-�z���Գ �㊝���~^�"V<�e�P#d�b3#F�3��cE�c��C�1�1�ٌ �6�W�(=�܈���i���p� w;�s���>��+$�ɏ��s.-8��I٥�].�Ln��݆@p&K�A���Z@��W
�o�y��}Z�X�nt(��
1jQ�ĘY��9��s�B�@�ƉK[�����<^E��n�T�{��_ZG�l�WC��z�)_�eo��h��)T�tyOo@O�R�g]��)����$���f�0����ex]���G�%r�p�;KcM5���/䆃�`��O�l�Q*I�$��
���&�4�
�~��a�����E�^ ]����$�Bv�M��V'+�_�r��iy�P��ɤ=B�)�ֳ�z�??G�Ꮤ!+:T��ȴ����,�K�=o�L�!�P�Kn�Ǫm��#AueV�^��f�@�T ���_V�EU*`6\���y�kOm�ѽT����%�jH�}�1��W�vϝ`�e.��TJ��ȫy@��N�?��zg0)�Q�Aե�]O���[ ��zܞ�p�
���H݈�ק�FďqR�k�P��@'�.n�幇�e,�V6�V��/�<��u�n'l�Aۯ��شϦW4gn�D��j;�w�55�12bY'�7}224%rНß�ye�1���������mo���kN��c���	�f6; � �4Ic�-�)ؐ�n�2������#g�,I'%;S��蹥� �u׭���񴉀�����+V�|�>Јhc�n� ��i��0��et� �h��{�����G��:�~k;�C[+���u�:>�����HG+���tIL��c�z,ܻ�qF�mJ�j�����g)����6�j��@l�H���.'\t�jcBj²O��q�*.���Wx��<��HZ�����K��Gzp��Fn�&<=�{��#\��H�({�Y����vVkt�e�d��*�L�Rc�\�ʙ6�V�󕾏���.��%�a6��+ۢ�0vqa��uY�$j4k+hI3أ�5ߵvk�4h]qqf3J�z�Xc2�>��4I�Ĺ��4��_�Ҷ��SM��O����G���`g�	��
��z_-�/�4�QL�]�x�^��������r!�t��.�XSN��p���Z�f��pȥ��*lpۛ�+�����)����1@2��������Þ�y!x��p�2i�ɟ�ϼ.�����I�[�n��{I/Na��ڹ
�F�ԉ�M�3����3�aq�Up�iZ��������2�4г^�K�u�|^�9L�4��U<Yf��oE�3��:���)3
�ث��x�F���4|��>��!� .�U��Xg�\����Z�]?��:�����S��J�o�g�����Ӕ�fk���8.�7�0���Vg+|��K���U��GU헛�Z{��a[���7<&ڧ2m͍s4cᒍ�Y2%S	Gn���z��D�G�/V���(��+�:B������Io_n��J���?Lni-<ah�:�
C��8���1W���m$�!�Ș���jGzk�c�`�%��������X��2ٖ������\Sշ\�vE[\��t|`�οi�h�%��6$V(�䮪Q��U����o�FQ_Mj��&��v1�u�>q6~��F^i@�k���{e+ ݭ'���	Osu�8[�c:����z�t��`q�O#Q~��xS�����9Вl�?�@�X7a�/�$�!���ĺq��3��چP�!K���H|}^|��x��w����]�:��
��/�ښ��Ug'��htCc�3�R����9L?��^c@I>�-���0W���ꠈKrn��醹�ϊ�	�)��w�-�hko� r|�nJ���*'�ŧ\�]�rb @��"�i��"�%����Ѯ.�vW��[n(Q5�N"	kt���'��3|N�2�w(ԛZX�d2r;l��������W��Bsqͥ��O��oU4�<�骊n�\ǓG|����Pr�!P=A�V��ղ^�D2�	^������AS��|���G����b�W��}P��(9W���ְ�9a�5!~d���Zt��N'�sU"fM>�L/D�B�Y1iP�����3����K2���������索�b�_�HB]�~�>�!��JLWV'����ɛ�j�!����ʤ�K<1xf���c��Ƙ߄�R^p�e]��vEf8��T�2��K��m��.bg�8����3\}9�5Ft�R�|���^[x0G�p��lp�����:�ν^x��J����~�<�#��<�w���!9�r;a3=��fn��~dk��.����gfl��,
��0���T|?ITH�J�Q��J���0�$tR2�l�b���Qn7T9j�|���8��5��x�2Γym��MG��V�+�.Z�C��b�+"�a�9��R���6��zs~�U}Fy�g���K^�/.S�i�K@f�������,2��}`������L3�tӆ����UoQC�vpߐ;dR�l_F�i�ޔjp �
wCe�@�ls��bE�>=0g=m|�{�����I�T��E]?��?�*z��\�͸��o�����}��-���WFMb���>c�a�����{ڂ��"��y��u��XS}���3���K7��p��{۲�w�w�yi$�U�6�Y�W]���m[Z�󵔝
Ϯ��dI���c�뭖�
AF����{��zb������:G/ 1�^�xރ������j�x%ZtB2�J�h,���J�  jY�v��nEz��q{��e:���GSE0�n�����P>͚{VCo��4�Gs�N�ţJ�^��9K�v��]�2�lC/���6���(7� ��OM̷ϓFm��U��=)mO~�1�;)�&�;�Z`@1]%ܽ1�"�b{����JSlo��0и��-��T�5����;�*��� JN$��gZ�g����"uJ_i���7v�3S`F����o�/a)�;�Յ�X��d��i!-b�U>�8Q�OCñ��
B��{�+��Ƚ�������7.��<3r�j=���)]N�<;Wඤ,+4�K? n;�,6��
�7IV1�QN�]��T������(�<F̖k;���7�ܢ3�1�lt8>J1<Y�ݠ�Eh%1n���!l�[��M���V���y���w���S�i*����s��]E��û�=|(���� ��W⊿�Zɗ�8��H��aF8�sWA�Z��]O�k;��ZZ�x��*\��IB�#�\�C�%��	L�6���'���X���S������p϶��9�9|��t�!F@�x�r1��׿dp�n����/�e����Z9�����0����S���`��l�u��9����b7�.��n�k:����7��4��.�{�Z#��P�]<��1�#�3��'��|
t���������[#���3zoQ�`0�0���^�$!�w���F��Do#D�QAB^�����:�u�]w���������9��Q�}ѐ���4a�l��f�tuf����7Yi�]7����
)4�֛%��4�U�g*��W�Q���Ƅ�#�SW}X����qN�f�ч�o1�v>;�;g�<�f�U�� S^s��{�謄W�B�9H��	�A@��eF��F����G��]i��5/{�V�*��BR��%�b:�Y��|����kޤ�R�Qh�P�K�s3��肒�]N�gт9� �a�\��~|ڮu|��x��"c�����|��)����B��>�ɅW���n4����=hl�&�5��S,����y��/�D��ph�K2&�Ž9ˠ&��Ryz_ݢ��ՆqD<�Z�n:M�և�<�$�|�j�f�/��/ӿ΍�-r��yB�J�
����0�Y�E�;��[�d�L��5����R���D��X	��¿�BI���\��F�Gk����_S� �`Q��AB�q�[W��@'V�#��R;���EI©X? ����c�;<R�Z2#�[�����ay�7X�`wf���0�f����]�uyO+��5��jT�J�X"��������1�Ó谛��cx?0�&V#$n�tݏ�{׎�
R1�_q������1?�w�ɩ�Ŋ6��
�.��ي����OO�~��<v���a��*�Ѧ���7M����'"҅��A�1e?R�rK%�E�.�l��R��!a<�y������팰h}���p�"s�2^����[�BY��������іV��{)h���n&b����R�duӧ[���G�kغ�7N��<�|����=r���O��ۿ���8E㖕�wݞ!���l{k諸�4g^���q�N�ɠ(RR"ԕ%�d6^��;��YkD��a��j=�*:���zv@xכb�ҍc��J����_�T��x�V=פ�7��o����7���E^�{;8�ҀrK����LS����i��/Ѯ���rƟ�Wu�\x$�gZ��C9�q�����~ R0A��4�Z,��B�)�L�rk$�G� {a!HQT)ŦLڐ7΀�p�uM��KC��I�W���Wkk/m�w�
�'`�R�B��.	��l����νTT����}��֏b6WKN�N���muu.W�>���ܦ�a�O.'�=wn�j�bU�+�ef�j0p!?t�s�l�/cU�KpZ,/I�⵱s�}R��`c�J�`��pǟ�>���E��À����)Ϝ�����5P��ci(�8M,R�;ZK�~�������u�a�0�Y�M?y��s����E��Ԛ��2$��醨�?h�9��ؒ�/1>��9d3S���4�F9y��6T'd$O,�"���Q	��"��x�B]���S@���Bz޸��0w�8�R���O��Z��H�&l]�%k�7
a�(�JT�hnu�j��	x�&6�;)p�\�RP���&�um_U�2C�~����;���0�9�ߌr�U�F�ۀ�.jэ��O��l6���ڒ�v�F�ƴ��0��a��FJt���y���o� +#������?j\0�t��о����q���K��G���ջ��~�x��()��p�Q�Њ�̻�\�nu�05�a���i�R��]0ܴ-hx��������ޣ�5�m��{����|��}�&|�3��V��+�QO�e챨��'O<e�����2�"�h�~t,ى��`������:-L�
ў^|~0��������}�:�>�Q�_�;Nִ$`$�h�Gg��1!9o2�#p �����?�;��%G��2]��}KP��b��g�_w���$��*ɼo3A�?P��Խy����l#*�b�1��W�K��4�P�g�"�� ��I��gr�֮_PJ�>�u�e�%����MV�����įT����]0�)&�5�)̀�V4r~6ޤI4�v�����T����5��x�g�Vt|������2r,ͅ�[�&,"r������Ã����A��"i*�>c�M�����91
	�y<ώ1m��~����#�"�Voկ0@cE�9��*�/��qH}*�8+Ӫ��E�.�&�B�r�����r��G��@�(��4�'q���Wof��JLτ-���%M�6}��U��Q���3��$�q4җjM�-���w�_8�rFB{���v��ǒ�9�1��B�ϣx"��)�|������T������X:��w��o�g>Gd5Y�<�_�EՄ=����*~s��ژ�����>B���t����2�K�g�|�ė�"V�5�˺>Z{�S�˦�-��R�n�� ͒m�Bߵ�~�Q�[@IJ�iS`A)>.��9�z,#\[ge�`�dJM6���Q�Nբ\�Ǌ���#�6���=DѨ�>����Z|�ʫ�h�W�͵�y����+��z���#�Y=���4@�?���Ͽ��z�b�Z'����Vg�&eV^�u(g"�-�����"��X�B���SWN��~��fm(�P�3՝N�٦{�u}�ZG��F+�sˍm�}5�Z�������
�7:�R�ܚ�j_^���!����T�U�{ىg�ϳ��
ڤw��ծ�/ �H�w�n���6�k]��7�/j\p��/���ܐ����m��
ɋ�s_/�w>+�o��h�o=.�+8M$Mg�҄M��G#U�!=�͛xqf��
�:v5�PC�Q�<i�Dx��g�lJ6�,-i�4�/������A��\��ڰ�L(;����({ܱ�:Z�ɺѽM_��y=������N�^��C��~�_��r�y�@Cs��&�'�L�{���^pIz3ϋ�x�؇�FW{8��T����/4~��(b�Pr��\�ɳ��K��#��{������|FTꯏ��EI:���[�r�i�+�W��y��v�5V�BX'�$u�R��M��v"i�Mo�j����K^�.��n^���O�xE��u��v�T
���Ja4'��&��� ���մ��¿+ֶ��:���������2S��U��5ub��5�;	�^�	� �R���u��*������G���Xn����ڡ@5����O_9����0�T,ˮ��:0�� �MPe>#�,bD]tR�{���Pqo�~Y�e��e���5�1��J�����,ճ������e�X�l*+���Bm2�/��*�A��z.����,k���q��%h_S������Ed�����?�j��ͨ�ZW$-dzs'�g��TI�~3RgU�n�(П�嵣��%�2��@niٖ����r?��,[�h�F]`}�,�~���5dn�ܓ��^|z=d���H�?��q���w��ԯ@D�JI�MU�yBx+CB�uވ
ᖣ�������4�p�V^b	��������7�}��b�xUKgЏ�2'����u��T�����a�T0C-gQ��!���1@E���0�7�� _@��>/����\aCܝ��[͆\[Fnǔ��X�M��	U�o5�: �'#��q�T!�ܒ��O��_w��܋��%��;��_ň��J8ā��"����ގ��,�XMo��`{��"��Q��,���ʔ��y�ʹ:RԵX�w.�﵁mz���Q���A��\a�ҫ:Q�^v7b���(J�͞���5}�s�D-��+"���Z���7� Q@M*l�f#������*�@Խ6`��i��Zu娡��� ��a3*�.������N޵(���7Dc|�t���Jw���r?�i]�)E�_<��V����S�*��ӷ����"A^���R����f��^F��Q� �MD���Mf熸_�@N�V)E��w�_cL��*���1KKU���+*���M�0�2{a��5GR���O����A���-�P���"�j�U������*g��
��kwa�P�J-f�%|]hOTG��&�b.5�,���B�%��Hm�D��p�Xt"��Lo���^ �
�$؀�5�,,���h? ��E��I5��,��a�BA�?Ⱥ9RS�?���N��f���^r��� �W�ɂ@�x�f�!��?V5_��ԡ��<1Pa����_�Ul �j�;�u�~j�	�	���V3L3�Cf�3�؀����l��8��&)����0��~75=���5���-���-ph"��M�L�~������r�q�|ȡ9�6��]�����ʀ�SWD�ĕY����:qTׄ�����${48�GNj\����l�D6�,��5�;'��F���������9�	���� �	�e��AM���qȍ%7\��	Gbʨl����5��wJ,	���ɫ�;�7s��7�T �=bN]M�~�4��yo'f��)�E�#��P:�Xݚ�xR�i74��)�¾���0c������ W���5()q0��tl8T��g�?$1�
��#�N��;Q��l//@�*kA��;|�3K���z!Z�DĤ/$��-�ڲ,-ͤΥ#��>�Tp�xZ���X&��A�\u�,ݞ	��i��F�:A~GY�v�e��gΔ
�[�U�+&��ŋ�/��3fR4�:�
D��r��9�+�����	�������պ�d�슬P>��*���<�F!V�=tp���O�(������'��SKӦ5;��]� '�%~I���dܥ��Ut��H�/Ϭ%/>�򙾐�3m��P�Ÿ"raoIe��-qUA�S쫊�x�$S<���p�LCu���`�?ȋX�G^�3d�8.wņ>4>~hs��%g��^]f�&���Nx;7^M�!l����C������9��cJ��PG���5�z�cP.K�8�� �>�8s�2M��[���'��ڶÔK󐁾�����c�Ҿ�I�[F�/ -/�8A���B��C�QW*�9��jx,�U]7$ҕf���c��c���3��nu�(|4�?a��rU��i>R>|�h��-�DI�7��SƗ��H��6=;��Q���ɵ��?*_��8�9յx�9��P�Fү����~���&�Ԍ���cQz�W�5�)6\[Qqd*}!ʠ�^��|��-qiN6�s�eP��9C�'����\2�kGزF¼`�ͪK�N��x@t���"�8uc�QT�����q�֐��R������x����>BI/�T��m�E�9GX�\��e�`�Wr����|��d���ZEG�_�*���_�!q��B���Lb=�~�H󋐢�,�Vxӳ�]A��<�sx�DIAo�?W�������rW+3t����x��(H侏q~�V^Z Z�ᰂQG,�V�K�?|�h����m*D"����|��P�ȹ��A<Q��]�� ���|�#��GC��%!IH��XN�2&�����2����x�>g�Zb^UqYp��qV~��(��'����B��$Ř&+EV��"p��:�sv�$Ǚ���ґ�h��I�c�C��J��֌�hT?�r��T� �&�S#ţ�=�Y���F�9,��
ц._{B�<k_�0kh>���������ό�I�݊��68
 
�ԂpO;��R_gB�i�c誓�4<8K]�x&������r���}*�P��.���Ak >d�dX@��q<�?�>��t�1���t����q��H���~�O�$NzU��0��
�ፉP��&6~,�������$��
G�Κ��Nk��c{�PN"h������0�: �¡�i��SYâ��QO���_w���[�1�C��Ր��%;�儸��hE.����Of�d�c`9J�t;MSS�J���Hl�9bF�k�f�8˘�x�`�I�U��gbxfĖ3WPS�j'�"��9��}��p��x��
2�j�pia �1~�����_v�Z�b �F��uD�Jta4�G����	���F�`J͕ʜS����Ad���p�� Lf�Ҥ��F+Y}(����!&�#�Q~B�g/��1��{�V@N��Gђ�)���n����!�Ԕ�#�� L� <+?�RN�1�"�M�����RNmpg�0�c�W��|��O�T��\��-Yr8����ѧ�c��.�j{��د#|�g�r���>b�'�/��E�+��S��!�F\��U�������O;���K���?�~&Ŵ*K��ze䎄m'|Ψ�B��53�e�ƞ%1}�Y��K�ɒ��0��.
t�Q���|��	:V��	���d!��t�J�p�d$گŒ��먪Hu�gd5t6OT�"ԏ�lL���~��,m���Y��C�{|��k�{��^$�?&��	�=���Ж�Z>�����zbY�IS�<Һ���X�	��6�y�4�Oa[�� .�1�~�w���uJ}�3�h�K���gy��!�4�SH巳������V�<��lj��R��P��0������+dp���M?�$�R-^�"��3�m���,�1S��Ei�ם@;&������_�.�9*/1Ѻ� T��h��*n���M�N���J�xvU`�!!���H7��>	7L��� �C���m�հ�+��}�UTi��S؟y~ð6�!^���6��kt4}Qw���N��g�����NJ����#5*�f&緹OR.�z��U�e����q7��J����R��#��<ME�>�^�=��T��D�쩅�|�	{̻��䦿7-�ƛfN+nF�+S�jSV=1��ҒL�TU4DM¹�!�����q�}���sV���qxx�V!�����-#��"&>�{�� �:>��A�+�{QL�3���tI`�xR�L&o � W*~w���!�U��T���t�MHJ:#���/i3�����j�nz���8_�+�|9���o $�K���0@��c�k�B���͙�ݬ��<��B%�������H]{��d �l���*�V�D4��ER��-�(r��v�/�T��t8�a{D���`C!r���!�1�x�]�5u�9}@���d���]�𳿲ubr���åT�~�����P��[O���>�l�7�,��>�p��\�;F;���ڗZ6�W�Nm˺�m���2ތ�v��3X-��%*���t���fvɗ�S�oTBd6�zh�7j_�p_���#��ז	�JOe���-�?���*63[��p�͞V�aݦ|�!��W��~E���ӗ>@\M��B?��Z��W�K�sy�{	��Ȼ6?���(S򄈠���J��y�����%$�ǽ�\j�����@)��GZ����{���C���pt��7�FT�f��V%ȡ}� A�A��@k'7$����1n�����2`�׭��'3b`��9�A��Um�W��\�C^3�h"X��0��CsP*��I���2�/��:��P~���F��:�R"�Ը����Jd�%���"�5�1��LX ��6�$F�&`�� m���Ze��(�Z�2a��`&��~>��ƙNL�Xu�U�̹�b�S(��-D�g�"�4H��/�	 ?YՁ��ܛs�g2Dd��H8���?�kG���Q�j0�5�� fH��ݕJjz'hRn����f�<RX�w� z	'�4�������̕�D�)<o_]%%��~"o8�_M
6t˜c14�E���X���HQ4�{@o�֙�K�x�=x~�+X��c7�x�j�$�I�h=��\�l0�4�� ���;,}�/`'�@�����_� gVOd�kߏ��]p���w����I�3Õ��ϴ�A�Fn@�|>X�W'0ЦM���������ո���P�&:aȲo1z���ᖘ�CO��d�%��/��R|@*yLC*z g4��"t�5<�It_�tE4�/�.l/O2��Σ������n�c�fͽ�+��fQU��ȅ��������7V�|煺�p�F>ǅQ1��yr�>E�M�-�gk��󗇚,Tߵ��NJ���}x��:��c,%�׭�Y���L��~$RIC���P!����$vھ�^�x���L>���!Qw�k)U>L����K�K�Y_�Kڂ�x���xR̗��?��99F4�?4}���9��`X�v�k�� b�L���
,n�>�A�(3r������(A�Ť+:X�]4p`�� ߸�ѽe�����Z�)��j�Pp-��۴oCL��B�}��<q2���MCl�H����`�u��~0wL�Y�3o&�R2�H����8�_�����-�A�/&+v� )%�l?G�)��|�Ko즵�`t���W�!�դ��>�c�6���r�3��p�4�+�g�04׍�켱JH�PG=������@�HQ��h�8���XVH��~�}�U�Ѧ./���Ub�Cv��?�BNb��X�,(�<
 =�Ɵ�l	i�R'�^~��l �Ր��f�/��K/T&5��=��̵������q���8���o��$qP2+���=�*�z�l��8	J�\.��\'^_8�� /��I�E=���e���Bl!� =@�J�#hR9�����h7+��T�}G!���#�FX�M�p�pZ���/�4�٤�ʍ�*?%��?�)Z�����ܔ��h5��:���סi��u���_��<��r�n.O�n�����n�6//+�
�a�W�IO��:���,F#@%-{�Bk��� @C��	
/mR��'�K`U��;�{��d��3�_�2�4�jOz��ݚ���%�������-^M����iC��D@����zm�+xn//��}��'��-�,M��"	1�E[�C�׍��EXa�*^��g9ǼYwO���O�R��A��p��9&��hq��3�P]d��@�`��tW���I�jjb��l��ځ���dv�=��4ڬ��O��̸��E�w��/��W�H� �K�H����G�7�R�Z�C����h�0�a�"�%F�r�l�KX��9�1���K�1��}ϫ�G=�)?۪�lL$�f�ɲ�8���8l��]n^��غ����ň�
��#2��A��x��V�4�w�Q���k�UY�FK��N9{���:}��!�ރ�F���T��{�������$��`f�	�p��������B
 �Ǡ$�0���ʇ�ߒ�q���%(vv�
�0گY[Ռ32���$��2���8�7�}a��9Q�����	i�����T|<��OU�&�'���Pdb��y�E��igw�;��s$zN$t�m�؁���x��m�T��I�\��В*�������B�O�R�d���T����^���'z�Հi]lO�$��p|Ӟ��� 6Lu�m�u�\�r�	I��\,�&�"mGLf�3�S�i*H��fH�/��-j�-�}x�1�^�^8���� 
����
�6��d����;��wah!8a�
59�� '���8������͵�����o�Mje�|n:�H��S��$	C�Q���x1sy��0�89���8����K�`8:>�����U6	���d�A����ݗ�sj%㷾 ���	#.܅nrK:ߛ���EyZ�VJ-�JF��	�}Y�{���N�b,T/��I�����w�<���P>������Z�
�ËB@3���EJ�rXw{���ڋ`��G��L.���ǅ��U�[�cv���ŵM76�9��D�
����>.�l�F�~)�^�z�A�2���<@WiEY�|�qR`�5��1��O�6i��\�w�!Ν =Sű��� s�k�H4M�|Ń� �ˈ$���2��Ԝ�-)3C-�%Y?�y�o�R�*Q�{~x������)><f��^�Lk?�9�M;\�·�z�?S�N���)�'f>��IϿr�>>�=B<"��+'9�$�ih%Ԍ�A��qK��}�L|1M�}ӧ�ү�S�os�����	�B+0��9������^0���/�we�3���xE�\#R����Q��YY����	a���z?z�O����1��'���y��[�x>s�e3���\��w� �	�3�:K�j��.~}6K���"��q*�!6�xf���i��#੷�e#ݨ�"xM�>�}��P0���lP6�����]�c��*W���a�;�Α㼟6�raS^ $���u�pɹ1�06|��v�:N�u�6=�X��6�/We��ٶꂏ�4X;�^�3�������,Ro�o�բ��{w��2ź	>�>�0'hw���g��J�\K4�w�G��8��#.�$��щ��36y$�M�ϝ��"�K�"��E��}pD��W�H�W��Sw?)�}{�]��,Fb���Ir�Z����U��`~���4�N��R��6�i�i��V��<`}`W'ɢ5`��^Jr����F1q����?��GyW���u���0o�wܘ��˅y�Oh��K�����xq�(�k�N%�yb�Q|��k�s��;RΨ�R�h�@��d3���J�N�_�k�"�c�+xo�@]=I���P���]������ ��8�� 2_��=���!�u�$�������3��o�z{�T�ܶ�}z�=��Y�^JW����;�*�+N���EM�,��x�?������1�<1�X�ʨb��/ߨ�<^�-��{�;��.��
�\��<$�0�H��9ow�#���T�+5�@���aO��O�c#�?2T�ͅ�|*$�߆��LvN��mi#Խ�{�������?�a��(/�YO0��h�w���S>˥N�|S ߘ8X.�N9��r�݁���F��e~�9�jSq8'*��,�/F8
Yf�_�Yp?=<WN�"��f?�^� ��b�ba5Wb��Mڴ3���E��j���YT�K�ղ+���;�K.7u��zi����e������O�1ئx ����������1��Lհ�=0 J��{���mX�u2�Fc,�2���Ь��
zn�W�R2U�9a�WQ.}w��&�����斮;��trL�q}�0x4f|o�$�e��Ko���T�X$Я������ӂ�[�s��yͼ`�`y���(�,̈́G��ة�X�^�KLl�8-B�H8sё���x����x{6��QS�M-��RV��Jdfms �����?/ s��V`K�y��}���	��&�D���T��B;P9�)�(�esIn:�N�ح�u��}f���2�'��l�5*�'D׭^o#fYb
xہf.E
�l�T�'}�*��zC*�Οk���"^�S�U+C�%ha���G'���!D:�O(�l�g�[�A�u(��?6];��󩌗󙻮K����<�� B��W���s��T����p���c��"�,U��C6f�y�|%���>΋O����SU���v|����b�[����������;��kJ�T����-��b\�������� ;pi��b��P�?�[��L��u�L�Yz�����ո}��x�	O��9!��u���72�䷚H4 /ip��{RUQQ��[{������d���w�ۨV��"3-kP�`�e�O�N~K����ˤ�~��;X�rS6Nq�pz<#�lWS"��b��ն�l�J?s���'�y���I&N/ܺ�q��u�'��T��+>J��1�	to�lN�c�Cz�����e[g n�>�&�d�kU7��g쭩�����t����::��UUs�
I�Rʊ����e���B:	��0�w���ڕ�'����X��+ڃs��B�L�	O����d�@�[Sd?y_=���13�a�|��Oo�RSK�hYz7�(���ݙ.'$�7�=^��ͷ�7pR��6H@0��5c�����pCyl@���������q��"��ӎ�I��R��H"�+v3,����g���9��_�d(as]��fo��{5��>�\�{�9*����Q��l��X� 99wK|]��c[ΐ��S?��0��P�_�HQju�Ҵ<44��j�i�gՋA�g/j;���������[�EG?�Ӄ�N���( N�������% �|�9q��eV0��^"2<�1�e9ˬT{���+�%�Ϫ$G�1 VK��{\��UjV����u&��7�O�h�E<�1��ٗ�n�h�T3y�e��Kz|�.m�2�����tϣxQ^Da�X��Ko��^���c7���-.����/�𐬒�mg�O
3��U^ӊ{/ߺ^P1!q>����#���SqB�=*b��cN�{~_���c��YQ�o��o+��2�G��1A�Wt��˳[s59`���]w4?<B�ˑ�d���y9�@^�b���z{�M?s���Z�>�_����76��k�/X0!�u@��)<�Lykq��p�&�:��!1h�j�����\��]��5��I�Ca��н��"�"�?}�?�	@�'1��J�o2'��S�����>;�R�H)v��.�TA�����_���{����	����|
5u�Ԏڞ��l'�9�����%�g ��_F�MS��Vmc�G�5Ξ�}Z�:���p.�}9�7~�)�Ƿ�;F�v!�^ч5�I�7o�M�?�\��px�K\N�H;���T�����^�y���1̾i���	�������Eu�x��������ëS�[�f$i��>!�=�{��;'�O�E#�nl����y�ԧ�3}�<����r����s��`tެ��0�6�g���B鹶u.�����r�%uٯ(�VlhI/dU&��h{��uV���m���|q��84��Q�78ǁ�.����^x^p�$Ѱ�.Te�+�NE������.�n�͙�_��t��r�����2�k��!2�$�m���z�k�%����FKw)Ua5�W��AG�&�TKE_ ��Y�-�Z�'˭�Z�m���8z᪏�֜�$����A���	M�(�L��7�����(mK_�q�GDN�Po���a�� 򓆦fu��&��}�txl�ۉ��k���0��|�:�n��1�4�{0N崿x����k��\3@���G��D?r�[�fP�O����~��ȥi��+}��L�����X��|�ZY���(�J�<�*���:ZN~ȝ�3�/�%��TQT�u��m�F���h�M�o�a�=����B~�$g����"\soȲ���G=���k�iY�ױ/x(�?�+����[I+��|�ˊy8��;��m
��J�G9RAWf���]U��ss��-Ƣ�	[������LI�_+G����Y?�ҭ53���Im�/���
�M� qZ�i��=�;Ͳ!�d�l:�#��/��wU�(����@K0�y���V�舆0Ggi	-�0ί���#&v�$w/K���CL���4�zۮk�r�^��_���F����Q!���Y�#$�Px���Wx�M.PA�X+���0��0QI�.����.F�%�.�3����T/E�N���3>���?��I N̲ʕ��,�3P(r�xj�S�[S��ۉM�1�|7�R�f��x(~�|������7:�pn�<������T/�&O\S��������%2(�^�%��W�������_��g����F[<v88:ur+�%� �������}5RAEL�g���׎3�"͹��c7�n�h�T�3�⪟XL�"�>�h~��O�4����K�����"V�'|�!�,WU����g��fLSa� ����`+�g�#��XxϽ���w%'N��>��*
ܽ��8�ץb|���q��QU�U���%�T"i����Rf����ވ�8��+-ы(���+�@?[����L>s6�Υ�R��Q�{̀';�${y���
��ЇIe'�xFh��q�h~���_GW%ѳ���#`#��mBe����/�е�9��1�>�zK/���y�:կ�^:�p{���h���"=�K��;�HVǋ��J���������	�܏�l���}�M��)���O���;=�[��"�0-�:���%d���j�D�,��Ze�/�k�S���k�U����h&��'��BG���{3��<\z�E���[�4��z4��?v�DgB\O��x45��i3���Kc�.�n�o�mO{"��x/I����|�:�s�￟�ƁOXL)9��=���S?�Ц|����C ̧`$�&{O���;�e�������eǰvK����x��j�\܏��U�׃%�����CyB�T�ϪK���"��r�::��M��UZbÜ��,\4����Г�e�e�@�VPx4�q_3��N�kQ$~c��sv^��ȱ��1wǎ:T�Tc�)$\���MC��}��![�H���Q�w�I�N��:�7W�z2��vrѵ���i{ہ�1׌Ȼ��|����a]�q��.h%���G�@��fN�������4X�Q�a�w�`M��F�N����y`?�,�2��z;O��_�YQ��<Wp+s������-;�{k�+��⺸�����k�����&I�,7��a��͝��RN��FR��侼i���|��#�D��i�2=�T3�K�/�#���:`�M9�陸�vT��tӰf����nf'��G��:�:����&f��P���_$�It�Fܛe���sOR?�d\NN��{�RXTyc`Zw���dtGX�#7��NE�J<1�F"\��~��1
!UgF;��`�F��i��7-j%S����~��3�^%7��M�a������d�+��0�/��ߙL��O�t~��H>�kn;(G��H<��s���s��b�"�6������}Y0.���:wK߲�R�h�� g��dM���bn`�7��>>XsC�מ�T7�!ʝ_B����4����0*6CLl���r��~�,f?=��h2�t�W�'�,H�w�S?�}��l��tI�4��˄jn�>�,na3���	%7I6�Fvz��_y7�����v��#'{�+¶�R�bW�k&��p>�P��K9�t[U���N1Z����->9�ۊ�ġ�*�Yǡ���e�׹l{�[,멟�n��:5�+Mmk���剠�i(M��$��L��I���%᧸g%�C�oL���i�G��#:��&�p�:��9�%��134�D�g���'$d/i�ѥ�ܢ�����շg�mx!�=���4<o�5���\Y�P�l�~JD0��� A�(�c0��9�&�`��0k��aYU\V�&t�()�_��NgqHF����B�/
�f^��ޅdɱ_Q����f�ȑ�av��k{�?�PFq���G���ĺ�S%�?�#�
��(sA:y��xJ��qIw,�U�ľ�#w#mx>}����_�&XH�duS�\s�=C�T��6��*qAƽ�(v�����Ȟ��8|���؀��8�'�>"���5�r>�RaP($��K���e�9͏,����i��ls�R�J^�Az^-��]0hX������Q�6k�x��+ O��{]�/<��9��}l �g��XGĚ�%oR��oA*]Q�:[R_�+Y��s����v�3��t��>���T ;���qE��Gc#s��h!���0#y<7����5�h�d���Y'�
�4ͳ��q���g���H࢈_~�O#_4M��U�a>M���&��ɋ?�jg=&4635ф3�X1�f�f������X��7F8,|@�~L�a��\o5X��ҳ�z���l�X%у����3��s�|p��J6�k/��y���ҍH(��*1@�x���A��*�\���;��3��06���~{'���:L)F�Ǫ�+��NQw�Qɝ��L9�FHO9x:d�9:�kf�?Я��I�S�ԼjWT.H����E?\���^_'��*���;"h�`Z�ȚU�d崦S���������%׼տx�C /���T�'���6+�z��tJч��&����q�<���8�I�aЕ���!O��>�9�kR0�o�b4�����TR�	�6��ba�b�id��Đ��b�K�F"��'��#1��q��{u^E	2ߟIbTp�'��M�o��%�u�4a��UIX���S/$F�J�xu-���Y��nҋl�[d��H�5���i�>&P8h8
Ny�R4�Yh�ӧ=��t�%�fU5G��i��K?���&e��G�KR�b����\��(�,��@��(KC�<q�f�5M��/N��8�7���O�C�C�ѻژ��{��!3x��Ȳ�ǹd�֧[[GU��i���@��֚ꟳ^����i��֡���9�S3@!.�{�Sm䊌�
�����DKF�Y�
��N�d�rk��D�Sv����EVT���k3:�3��%Aʪ��.�a��b�9*��h�XY���UF�?�pD�ԑ/�,�"xG�e�wu��g�k��9+YI�����k-�<K�"����� �t�c�6N�[o��Q�D%�ec4R3��\ʬaM�<fh�4lŞ�2��f&l\��?��?����pι���f�k�>���-Ig~c��r����K�k�A�HZ�j�#~Ͽ�y}ߟ���KO03*��!��)+Ϊ����=�s/��7�X�$:hOM}7Q��|7b.ܾeL���øK�)�Z�'9�l��������E��7��Jv���_�z��u\/�6��n�qp^�P�f��'��`����͇ة�_�F������_D�ə����c�����Ӧ���,5A��	��i�K�UF�T)���*o��a9�a� j�`�zխ��o/024za����a:ۃx����P/�ȿ��i���ܣ��/*"�� ����te*�{0o��o�6E��"vS8�z��{|�+vgJ��>
h�>��M��.vά�m8䕲E|�y�/(�#dK�;��>�߸$��*OGy��x�S)0E?�a9���wu�G��o� ������}/�m����$l����BlU�f0P��,f1U4^�v��L�ͯ��bG�[�'�)�sv�ļ�zv��"�	��9�Z@{'�ƍqx��P�5�j���<Fހ5J��ۜ��"���+����\�G5"��C�ޥ�<���BTs�᯲(bn�X,2�43)�y��ѧ7M/��'�u�m�"wo79�E�&��T?��������@�{�з�B|��~ �[�p���\��t�t��Ñ���S����S�����! ���|Nf<�⒒�@4��#�j��t�������VX|Iv vJ|~�JCY'Z�tG����];�A@)Mtr�P������#��B��B�i�y�
���[ܿ�t�m�z���SKӱ�t�.A6u:m���8}�NOi�ni2����/Pm_-��w[���<���讉�Z]>h�DÌZ�3��@W�J�>s�3`[LAQ��p�7�Y\,\�H�&Z�4_4�=��i�����3��F�]F��wO
�l(�?s� e	��os�H��s=cJ����[}`�ݕ6���u��Dy;�tז�����b|'"�oF6"��$7$4M���8�%����5I�����^F�h�p��}2�#�������G/�O�
�I%�����"+G�G���������.��˾U��Ҩ�sS�&�i���9�q�etg�c6�v6�a����Y���ʶR=��4�'(�F��$��k�ߐ Z�^j��������-U�os����Eb5G���8�����8ʄ���d���Qu�_�=�6ېm>�/_`hT���:1b3]�Nh��EB|4R�+vY|�101�Ň�B�S�;���o@K���&��H���S�1�=�f}���ʽ�������>��od�`hc�����-�q�`��l$lft�o�,Koa��*��|���@���(9"�e���eZ�>8r�$}~+�2��w{�B=��Z29-��Y~]u��N�xLH��K
;+�\��1�%�(F�!��w�N�@U�{|��������u�U�dfB����g�K��ћ����,��m
z~��;��WI޾�x��ˮ�`f����3e�D*� ��{[��50��A����ⷍ�ޥ��1]��v@?�&r�o�AK���[|c#����i����$M�,��a}@�;S������!�ߦ`��m�~B�~�䪵/E�_7�J{����C�l��xB��NI�=-��T(�l�wUl������6:QG����6�O��"�3J���Ǎ��C�u毾$��w)L�����[	���L�x�\1܏_��<���e�B�o�����ߡ��߀+��Zv�Ֆ��
�������?�dW�N;���j�|p��3�-�my�`G��59h҄a��K��+A�4�x���Z1}ρv��
��N�%��w��] �O�lg�gC.�y�GٯE_s���A��GV�O�.��������T�F�5�n�# ���~��q��V��#!p���8V�F��|`
f�첊��hn�WfGM>��Ia�)�%��k��W<�%k�@羏ZeijL?�ua���y4,^E
�}<z\k�2@`9-�G����j��E>��)^d�)e��2��7��Q
�s/�Cf���|�+�e�;��D��/�,E������q���Lӗ[��~��Aj'��� ��'z��G���݇b���3���c��>U���R�b�O	i��Dn*T3����\��[%b�I�n��Բ�\��@^h0'Q�ܫG!L�kS����[���(��ih���~}AG�X��u�+����*����k.�׮@����^���
��?,�t5יijQ���
.:K���j���1�ܕ}�g���*�(��9I}�i�iz(���Y�jJ��(�C�KE
��IZ^�PS�\o'���v,�K�Q қ��ʼ�{;{g^�揜eQ�o�$���s&y<��F��M��~�s�##fu�+��2C����N��*,�}�½��e��z���3�����ْ�h�sY[E�B?���`�'� bWBMw뎹�C�Fi�#�KGO��2�"��H���0da㐿H�yu���UK׽���=�2ET4� �ھ���Ӛ�+a�{��.	R��b��>5���Z榏vʠ���󥥧}�:~ǾT^?�+����V�P��+7����Wn�,��jܒ+J�|�(�U5I����Ts���H��s�\K����Jm�{�Uu\\3Ƒ�x㢀��?$��9(ݟހ�����,���Wl���@��m����J��X�i��ڇ$�SA�N�ⶇR���hV����^��b3��>�[�G]E�qB׷����#��_�F}z�)���oU�o �ś��q���s��vo����� ���V��Ѩ����oFV"��h��F�e���}O���)�x~v��!�7� �q�����$c��nngi�FG���ZB�na8E�5�ι�O�$���wH��7���1MO ��|G�ZM4FoYz���_-#[N�Ht�{���[��0���S�\A(hW�t�$i"I��G�����[�҉����Ė��$�Z�BS'�� ���ަ�K��h���6��Ggb?tՋŰ�*���.�mN����?��P��uEގ"L{����B��N�y�&y7�2Ƴ]���}�k���ɐ)%��B�N<�T���LRfГ��
�Ads��mO��@�i(����}f^����?�x��Yo�
x�{�e����\k��q��\P�?�B�"& Hh]J,��[N�2Q%_�-O��[2M�:�|t��7]�:W1����2��Ღh|֞-�%P=����{c��L�o�D���B��jUMqi�V@�Ϳ��Z	� ;D߅�F�M����G-P�����3� �����_~�����F����;���J�����pn�C�cΗ.��7�;Ǜ�S�][�_�\��Ú���Rdp5ޔ>ӁT�_�����&���ЦtpMp6�_��[�iZכh�_p�5q�Tn��+��1���K�T/m����M��0>ɶ%�I�)0'�5Su������a������|[gv�|;�����?-C��������K����"A��ve�9j�%�1�ۼ�"R,,O&f��^��G�|t=�.M&���JQg{���
�8S.m�w��j��-��+_�əCK������慑xI�B!a�t�9[���؅tV�����K�U}�f�)0RFC�NS��t���\񏘮�abq���9Al�|�|8_�OC��9*9���4\�ʷ�Ж�L�Xϭ��l�W�&c�ҿy��]�S-q����_Ǯ��GfJ�<�LC%Τ�|7�:��)�^Ü?�d��f곲Ar�F�h�@Q�5m���#��A�$�\��P7�PU!z!�
4�˴�x�*�Y����pZ�v$��w�F�-���7�����RFu�7��	"�m�0��g<������a�j�ك�f���DiR�<f<aaIwy�9��𹮺P������b��V�&0��0]'�c�.��園�Zx�ܒ�(h����p�eԛ�|]I���n�����[��5�J���I|2��8V��[�" �@,3�]�>324pR,rWSa��L�؆c���K�B
74��ڇ���鼴����:拯����Y���W����G��Q��"���Nr~�*l��e�#a1���������S���ڌ���]n{g�.᰼��gM�ß)���1�6��~���VQ��A��R���;��H��*���*�|�a�w(�cj�rXto�S�7�K�±�<�z2v���z��0�$3������U��U��Lu�n�#�YK�����=�:̉��㷸�I>r�u�~���٭A��:�E�Sb]W�sL���soܜʅ̕�&-����b��U*^�a5��.���rԎL�ܼ��}��B��y_/5.DΣ��jۮ�n�	N���'�>���N�:ˁ@�ѧ%?o���F%YL�*f����Gl�h���l�J�<�Q��=o�*���8�f
e�7��뱀�t�s�zu�У��Mm_�E_��3��g��U4���Z&�#���L������`W�1����9OB�\��篡�����x1��W�60Y&F���,��7�2����l�}`,��^V� օ9<�^-�����/��M�A�z���Bp*�Ā߲�7a�z��)���S�V!|]���>�pE. �-�[� v��|ʸ}Q�K񛋹f/�c4���~�Q���6;����a���/�������Үļ�!{��X���w��vS,�=I���g�6��
�}\��<Rb�l�I��G	�5����� �	��%�G�,c��Ț)���'G6�������.����<"�&>[��.��_> �4%�[Z;"�6=1�ݥ~�oN��x[�̊+��dA	��a\h:L�m�a�RY/��x�+�f/�_GW�QU���3^��d\�v���i:��i{C���=lXӼ�D��W�H8c�̜Y|o	�2�7Ji�߇8�hΤ�7N�Oc�g��T+�����r�5#�. ##����:��S�m*�ka%��=LE�����}~Rc�]�3�*�L�������&�΋�i)�)��:9"v���R���)��m�o1V����H;ͺ��])҈��m�m��ܿ�;XSA�j�h�<��Q�Ü2>i6�+#*��WTM8�1�.^�$�ћ��p%���?'��&�+ɘ..��ì�,��p?ܞ쏖�Y+�zO�`��d��a2nE{8%�*^o����G�[�rkyk	)� ��aG��˄�N��,��Qa��m������h�ޥ7���$D��6��DO�DT�	��a'TU��rDԟ��?{u�[�	 �by�QQ�0w�\V}j�$��c,��2�X$����U�������JR32�셮%��
Ի�Գcxc6�:k�2_��ǔ@��~���Y�ѩ.� /���/jB���^(�(��l�W��\|�ta���(^�_ۗd~��dS�UO7ޔ��"�8G*�;�������Qߕ�,����X0]�^N��f&d���Hho;PU�WU�!��+ae��E��i
Q#/�?�t�v�B�I�a���|guFE��e�%rC�Yx�XT�\ka��4/P�U���O�1σ<�>˿�����@���a�v�����A���k�-�zޤc<]��2j�H���C���R�ǔb�a��C�W<��8=?�K����Ve:�gD�b"{+Γ��|t:���yRI�ș�ރ��o8��q·���<�xo��i�=G)�!����D��PŪ2�Aari�(�ܦ�t�	^��:�bLN.��N:����TҸ�l[��O+�+�2����SU�������s[{�'H����m�ay�����ۿ*�!gS@��:y%b��P�Z��$�پ;�L�y펹I��X�8
E�/q�L7XG�VfH\��-�%ghV��N�Ȓ�0@�NH����w�S�6G[����ͼ�m�S����}�Ύ��ر�~w��7)��yi�0����-v��0��<�E�F��d���n*N����G�����ٲ����|q@�m~���c�/�U�4�{��7���=6�6�<{RJ��t]�π�
]w_P����!��6�����T	
ױ��t/���G)���Ƅ�ғf�Ȩ�� s!��W�6��t�i�w��9��,�A�ߪ�o9��l�W|m�q*I�M�Z�߳��ܤ�t�k�9�[���ʘps��71|t��g�6q~�̄$�Kj^��ᖱ������`�n�%��Gr�訞ha�M���H��޸»h:�S�LD�B�rp��e�Aõ-r��lϧ�1=����ŃU9O&z�_��	.X��bi��h_*⾴-��sZ�s$�rH����gu�fv���8��)#�M�bA.�N��y ;`�E� V�R�sccy�[���}�������/��O�cJb-�����QA��2����6��`$L@�k��c�$V�ΰ�{���_��j!]��~2��Y�*�����x���f} YH6���U��}_�##�&B7g���'��]�0��EI� /��z2e������fV��n��_L�ȹ�q�~�,���sJv�j~řY�,<�I?���`+Y�����;�����o����ҭ���s�U���5�0��2�8�A>l��[<��\�(�@4��E���e�Do�[�P��ʙ=`ò,��1�iptBڟ�~l�`���Wt9q��=��_+���,p0�V���[�ӧ��.5E
�����B�/Y��T�����i���*�F�?e��|�9w 	��ū���],��&�捕ӼĢ��!\vK�v��h�p���7RKj�W�υˇ�TqM4��n	�3+'(���f�-ۭB���d��˖Ø�i�Ou���>̮���uSr��JSvM��P���X��4��������O2�k軐��щ�W��q�Ɯ�����q�0O�3�����]þO�0>�&�d�9�����G�L�]��(�L��:���{s���X�1��ß���` 0�y��H��.���Ro���{��R�yW�#�/T�hW�����C�_�ͣb{k���3�I
�f��pR}��|� �F.� ��h7���rc�Q�n,������J�����l,%%����S(X��sU�=? dR���,�`�G�ٰ^g5JB�.oថ�$��-�l��5�Z|�5�2GFd��.Gmm��={5��"���>";����}�|��-�O�/�C�d�e6�g�n�,-�����Κ��
>����D��6�FOM�`�vm���������a/���M��K|�4�����R0^K�������Z�,J�0yw�5߾Hn)�<���zNB���\5�C�4W�;��������/���8�M`~����`�!�$��{��o)��t�k36p �� <�&�K� Fw�8��l��΢� /��Z��)ɊDː2"g?+�M�;�Uٲ(]G��g��^e���]�m	@���Z��h��@��?ޟ�Þw��M g�q�˂{�s��es�) N*���E^�bYYOc�lC	w�M���yں��jT��r&-���o�[}���s~l�l�"��N"�J
TM�+N����:
j����a��_�m"hb�"�'�<�g���=#/�"���z7�5���d���9�x�g��[zA5�����7��Wi�]������}Y]l�/�o���BW�>����	�ob'nB8��+m߅�n���W=�5hu�_U��̝�6��ϸ�5l/]�xt�y;��/�]!)2^�+Th���������o&>��}����iI�)*Yێ�g��	���_]���d�L?�i�R�B�)U������ު9�"s���jb�|�̑X�-����F;��W�{������0�q!�y�� DRTS��2`��*;暑�D'گ[�ˈ�E�Ҥ�\z9O坬DIG�v�����1M7�'.(�*籈��������0��ܭy�~�A�ؕ0O�%��o�߰Aa��u;���1m�#C�2���禈5��@�(�c��>xB�Ŕ�靽�V����M�@��-Mv��`�����#����ڕ�B��,��H�a&����� m�����p��k3�nL�Hq9����'|NQF@��	����5��rһ ~F�ӓ�5�/퉺?:�D��Ǫ��G���B��l�3>z�M��^R%�ć@�3���[q@���s��>>��-���F43�u-j�<��@[���E���-�OeF�Yu_q�g.&X�ˬZ�s�D�F�ȸ'�!3^A�71o�����[1�Q���.�oq�Vm�U�)������|��1����R��\�����d�S5���x�m��5omcq��]6B:ם	�ү<�"d���0Q<�yA݇�43ﶸd��^�N�U���o<�]��\��P��N���V`��r�"�4E
y��)�B����^tmq7RW�[C�?��wqB��X���w+��ԷG:�SX@�OK�MH�Д�ބ�҄b��_,���w�(tz`:��IW�x7^wy��|�p����c>�<H��ƽ��mF3�n��@�cI�>ȅ�=Be�&J�P`�m$Q��u �d-=�S��1�5)[���:=��������x1��i#w�1�H&�Ƕ%$�穞_2�b7a����p�	$A'M��{�k��c�&��\a�u*0 �T��oW��>�$�$���amT��>�Л��/U@�Z�]F�p> 8�E�*i��P�O�r}5	�~M ~�y��EzoxU�`�a�Wd�G�aoRD�3�}��JSh�?�����'�Ƅ���R���J4�C�`e����K�鷴t8~GK��1�g�l�zc�M|�ZV�E:u-ʵwY+�
m�6�n��n7��Kh�*�u��t��C
�(Q�u ����m��'��\�cZ�Oߟ�}�R���*ϱ��\<��$��p��j�M�I�c�^�&lzA���Me������ݓ��HN��>8
����/d��J�MV�3.w+2>� a�RE^��]V�h�P_5[�Ԕ�6�
-O�ć�&�g����}��ȰQ�3/-��+���JRfe	3�_��e�`��q�'���h����P�������͙��?�BN��M�1Ќ��/:%�N˷� wOc��ʛt�烡��k��j�f�zދ�宰��*~Bcw6�!�$�o�j��M��G���,J�0�Rv��ڨ�3M�_�'��
	���@�m��2�]�i�Cb�0�j^n�z>���A��Iho� �����4f�(P�.�|��!oX��v�b�٥z��i�]��A�ʋ��\�Y����2��0�Y�X+�Кs��w�4�L1�V����/Q��ޒ5<���yj�!�q$���T�Lfv���@��uH�ݟ�H�HQi9�AN�avU�:d�x5�_�A�f%�����Q�v�I����Ƙ�CR�і�����=����ÿ�p�7͋'�ݾhy?N��E<`l!H��!m/������s�y�9޷e-A��m��7 c4�0u:C�^��w���Wd���Kپ���L��p���fQ�k�u��,�so����n��k�D�1�S;5�g�k)��ܗԙ����?���Y'��#A�)�ۛ����iB6�q&�B�z���Q�B�����k�`ܼ%����|��B���ϲ��Z>�H��.�ˠ���8;��<p���
%h����ތS���_�0kdJ���|]�yi��!d�nd6�;�-4p�U�V�i_��'��a��og^������`>}�9)���Wl�5n@O��X��3���q#%��D�߻�o�gj��'ߵ��[Zh 4�}B=BK�_��k�9ryj�=�o�����_�yj�i4��}�*pA���~Cz�}����0Y��.}zqG���*���!އ��&��Vh-��e���?��} �TGZ���!*g��H�r�D��_"�[���W��4�ǷK{f�>�~Va��0�G����9�C�cO^����S��c^�	6�m��8�3�lx�<a��M�(|L*)��W����~j�n)�.��s2lrhz�'B��I���osQ�t�Ey6T�?�69�H�?�-�\up��� 4旉��ܗ�;�oS��ʯ8��g�16~w;��,!�x�4v_MP���'�}?l��4���iʫ��:}���'�	�$����5ֲ+b_:��6�}�D���\���Y���<�eVŃRj�2�M���D1������,�R��R�t�"��3-/�����LO��+Mh�8�B�1���^r�fg��1��"?p��{K~1kT݆�fTYE*��V�3�Crw\�VH�H�?Ŵ���]7���ɭ�V+v������T�[��99>G6`0�߈�����ZcVc��b�b�>�3��?0)�YD_��up����㏱�o:��@w�߇�a�?�R'�I�?���*>
k���w&6P�i'�q}��a���JT��Ԛ|�K_'���@ >��z���rpT��ѹ��Cק0�Z����u��ǷUj�-��J2�Ǵ6ҤA����%����=��v����,O��#Vܬ.�Ro)X��]xA��ufv`�}J+��f��ez,�@<�O�����	7�#��)PxGaI&t��cyB�-��~p̵z����ۗ&��pW��/6?ݱטs&%�3T���u����kn����3?�U��o�#��bsR_,�#�2�2�uF����g�'zi�V-���>��I�jL�֒u)*����Bi�>f^9 t<��@C���q����T�夠���f�C�d��)�CKo��c.�I=[���b��T�ߦY�U��h�޼�&v���|W��w2_����}�A�v�AN���Is4HcP���k���݆e0g[d�ɪ��X�b.I�`��$$T�i�*ݟZ�'w18���ڝ����Mؼtj�J�{uBy_B�M�v��K�&hj*���t�>7��iw����¨ѺW��`��,��0�K�{�;���>�F����u�1�ۨ}N�+o<,�S��у����_,B�,z�YJh�ATun�6=��cVL��`�X/��	��{�j�-�������}�c��Ȭ5��Td�J�3D��`�^���L1c��ƞ:3��Wׯ��R�}hMJ���1�O��9�S(�����o����Fd�ݵ#p�����`(����GO��(�Ʌ
�-��=@�a� J�%E*VL��S,�,Ŏ0`<`�$t6Q;S�ij7/N#�A�8�q�->T�Ћ*Y܌3^�ޟx������f��V�n��D�I���C��i�\ρɌ�X�a��J'���Tq;L��@T�A�x�ѥ�� �L�՚p<#�qi�=��B���]A������D�{���]-�3֝�@��#wõ9yDBԮV����`���-��-):f���
��@f�>���b6�Ή�RI�N�΁���<4?�B)�߫8�Yj{�d]�ǫ��*��HmF�ry*��ġה0w����/�kH+�+YÕ��F�n��ŷn5���4��5iݗw��o�eZ�BNu/�{������߫zVͼ,��ĵ�yj��.��<&�2u��{+�PI���a�M�}�3l=�gN�N|d-�)�?5�(�y�99�'�����i��]����1��2�^D���&ɜZ�`�ՓoB��V���y ?]%?LC�ƣ[
o%��V�!�Vo�6��eF��҇.:��^��Z��j^r��?�=�\�)U�++	��>�b�l&L!� �������Vl������*�ǣl_'?��s�/�Ɏ�-����� ��-d��U=�v��.��\�!�F]i�XS�*Z��\2�)����j[�X��ÿP�dC�2\�xx�iy�V��`S�=^F�������=e���ZM��	{�����Lm�W��	��X'��;VƁ[ȏ\�7*�A/�۱pM�+���`��������������z:eQ)6>�n涞��L�7_'\��Z���zFϲ�_͐c.0r.԰�<�B���˱� �l ���x6)3�5 xԽw�ԇ� dR��b噃��YV�����2(�*���M���>��Bi��A�OJ�'����Ow�@��st|���1��j���s�	�;�z��vu���'��ao����]���_��)��� �D�:��6{:�GQ��\�S��k��)�ݗ�t�����{8Ϊ���U>�h���b�8Oؙ����5���BP���JWu�f�p~�S�} �U�l���x{o0��NOݮ]�𢺹��j��;�e;D�þ|��Q�H��J�);w̕Qo���K#�DF�����a)b52��������qiaJ�iR}�����'�Ͳ��7}�{���X��N�YG�;F&!�[��T^�:D����B;�u��ja$�E�'3����t�(~G; ا�NH��+��
�P`^��~�\�*�Whỏd�YL�Y��3*Z�#�6)�K�ū�(�s6M�+��ED�
n�Ev�j�]Q�~�VI6���AL���<��'�I��[&��5\:������P���ȷ��c�E(�Â��8��U�
BƎ���r�i~�:!ī��iy��@7�7U[�G�:�2$�)PTJ�u����^0
�B/���&���}m���>�H�1��{C�n�v���w�� {7�ؗ�~=�A�An����[���Jd�l�c��|��@���B��&}�$$���6��>�w>��zqa�l���C$��ac�;��mR����(��h	���o)iS�~x�����)���OS��W�:��6�r4d���G�n�MJ;iH_��.%�K�v���!/�F^x�v�"���Ʒ�Q�_��{�/�������:vf"$�4&>BtKأ�T˪)������j�G�,��)d�yͯh]����{�Rmf���_^�Y����C�X�}�c�! ���LJ�4%��=5��R�ܗn�4�8>U��ML��^d���=�l6Q~ ��<%6�v@��{̼ұ;�{�-�6P�	���w�����~��y]��`�h�m�����ub�.��	ch!�쮔�xcó�\"��?���j(��f��|c�J9�m�]"m��fdWB�ia9P��$\u�+֞+���y�"]Ȯ�Q�ݸ>ժ����P����P�(؁�ګ7-yS6G�9�Y1Q3Ch{�t-���I"��'c
T�^>Q �o��hz��@ӉӇ���+44�A�=��_w�dd�b]���mH����§*�9�1�%#2�u|���ٖ�����E��ձ�B�i"T�ӂ�B�\��#�'�٨� ��v�Oɸ�f��-�`��翂�xL�Q���O}�K�A��"��-K���=M���hs�E.z\{V;�ƻ��7�m
�(S�6�@+Ab�?�������#>����v�-��1jˮ�g���o�Y]&�h�?�3{T�Q�9�Zh^�;1Vo�m����A���m�X�'����T�xm~Y��c��X�5ף�W�v��aFg%�,y�n9I����b�>o�p�����)��$��M�K,G�h�)�^��C8ɿ��b��G/���eމoӏ N�?���XO]�$L�C="C����Ǯb }���Ww
x1�yZ����3��-sy�^K���,6�9��������.��*� |�sg���'�R���ށ^]���"%���Ą��fF��[�/U�r�1O5��:;�CIiH(ͳ��}k8*�ybc�^%ށ�B)E�ߗ0�2��� y+^oq��L�gjo2aK�t�v48����[��»��]>��r�~�� <��߂����8��y'���sqU31�$5cX\ǐ��X��:p�8t�XW%<��f��k�7�2xe70Ub��w�[L4(γ���ߍ3��U�������e%�\��or�p'�=���ؐ�JGU�[� ��ٶī�ǀZ�E��=X���j��=���wuL�#a@�U!ʩju����!�6��D9��bJ?ʶ��5�TW�x7�w�����&9�E�����ͣ<Ǵ+��e&�;b��7̀��/ݽ`��^����36���$�ښ5w~�2��gx�vB V�žw���J���� �I6���n-ґ˂qn��li�'���>?5��@A�(m~�g��H�#�]��+�hϑ2n2:�®�#��D�T��#����<O�t�#�ѣG�XAf#k�:�ϒ̢��8����4�w��.��Y������;���wqeAS���.�%�F��NdET��m���mo��� �W�\����m6�I���9��Sq;͘� 7����4a���uS �\�m ���%7#��{!DѫN�_M�.��\�x'^���R���#x,I���gdz�	�����V��_!#87o�T����s�&�L	ܢ�!M��t�����#��ejF�
�C�T��6�=ɗi��dp��$
n����*ߘ��,u��!�q�X8X�YA� ��S�"k3�:��첤��g��Hc=T�����!�.k��R�Y��nJ�J2�v�Pn_��|�M^�Ǐ�t"FE,_ZE�:���B�bca������,�'�0�&�۳�d.�k�k0�}�~��y�hǓ�_p�oe�]�*�M0���=���~h;���o��y��D�G�t��?�ME�Βu�`<)v($-b��U;Y�o�ҝ��#�ژ�O���:�}���ɛ��'����/��'=g�ԟs���3d�O�a�Ȉ�k���x�fb&�!�rg7��܅��HS���G��y��-��7�Ѳ,\
���X���/��qFs�M��=?���D���f�{~d��x�*	��R�2S9��X�6�)�5;��mV{���?:��ٮ�����ԝ|����l(�1��j!�!D�F�ql.|��,���� 4�>�$�^��F�tB]��_�>��8F�a�!���s��5I)
MNi�^T�Z�o����L�ͯ�{H
/�Ul�!1��;���x�iD�Ye-Co\s���N�}V�����=���0������Z������\��^̿g��, �o�9CI�w��8bw�"�#����Ahi��Q��C7�§<�-)���<۔}�J�d���'{�/�2�/�@�[��۬@ͳ�i��g
���M�!�L]!�d��F�Y�N;MD-M��L�j�)�^ ���p��٩�1Wp=��b�bVAj �Ȑ?�ns����=��o=�1���b�G�>����mk��@L���ߓ#m�c��m�;��$%UbXH��^9k� v�	����	^IUj��i���Üo"bA������T��:Vum������;7)[>6�}�
x߆�l)�@��ۯ���r4\8������Gx ��@g�D�%8Ԛ����i��`t�F^���t�_ռ��0��/�v�d3�q����]Z��}���z��X㲇�����Xp����h���ϴ��B�ei�$sv١������*sE���lY'�5}��\��C.%���8,˱{pi��}է&w"*�s�E�Z��(��"�K�:溔f�*[�-�d<2��Q��Ә��Yu�΄�]�F�]����F�/�Xw���H�:~'�܎1���.�XǱv[h>$�
s!ǅ�;M��E/������w�P��EXOF��t�;ľ�&ԥ�F��y�c�AU�Z]�H��έ�{H���[W�`.L���PU������ݿ/�J+����=>y��l��d"r.ߊ��	�<'�Oz�+���I
}��AA�\_yFB/
%R[	�+M|�"}ʝ\�Ftܔl�^D�ո�X��3�I�����1�����G#������5K��2�t��9�Mp%��"��n���^���M���-u�7tF���:�5'��tf��I������A�R�3�J[J��2t���kC'^�˜s�c���&��gT�_D�/�T��U~5c�i_x�� �v��>4��+��[&'�qqF�MkC��]��N�'��<��+�{����(}�s�o�l�\�����(�^�$�������V+�9�;:�� Z��3���^
T�\��W:��*Sx�e��-P3�tJ�z:�!5O6{x�V�"��Y�Q!��\,��m���;c���OVvy�w�h>�4�׈_�.WV�Ln�c�����_��\N�#�;T������8@ǿ%C",��Z�˹A��#��Z�%z�f�W�2Ca����!Cb����k�������{<������8�5���2x�9��N���'�H��֦,����A����W�:�Nq�[	�Ń$�x�dH������/(�7��M`o(��p%O���xp{�"L�����$Y!�!��}gĕA�e�֡$�Tde��p?�?s�۟e���?��K��5 �Ő��2T+� �N���_��Bk!q��dC+�(��Ǻ��6
kT��r $!11!;Bk�&.�-	&������<&<SC��n����'�w�9�U��r9��oڵ%��R#O��X��ܡ��C1dh��j����B��j���2��H���y��]-���@�F�ЈfI�k7]���,4*����dC�����W[#���=bCkXю>����~���a�?�JL�A��ס"&Y���T�`��ץ��,	L%`�گd1��c:�dh,�C����4|�A��ǈ�Q�
�E�$��W�a!�d�xh�9��BCD��ċ�R�������:;蓄>O�Z/��~�U	,ӱ��"�DO�U0�����$e	C!�X�]$%���<(�Sdg�1c�Y��s� �~�B6�0�W����xk�m����W�Q�)��G�#Sg0�
�� j�	!���-`f��#(�$S��h�� � �*`��������̅��L)7ȥ��Sǚ� �������@�L����fX���l�D�����C���@x���i�l�� چ]L0�"D��&6&&Mb�'�B?�J�0���x��<'���xN��!	�5~��� -    !1AQaq���� @`p��P���0���  ?� ��o�1q��A �V��)���d��?���j��j��2o)ex�gME?$Ҩ�S
���3�N4���B�f�=�{ܾ���e�e<�z,����7$������ �!��0+W��� �Ɋ��S�6J����䖲�7��@F��b�k���!�� ���zE�w�%�ܭà�E�Q �ھ��@�V�R�%����.� �2�lA�i�����YB��5�p�5��Pr��� ����5<lG���4#���f�3! �������� ���GC)����f(IM���n���!��&� �.1(#9w�n/����opԋ�1o%/�l�>��鋚-��Ն��PE,���f�~����UX��� ,�ŀ�K��� ��;''��������@ø�� A;�ܺ�*�$1�E�t��_�@Ny�+{q?�K�|���<���k�J��&��Q�Xs�5#���g1.� #V�s� �j,�WK��#������lY�w�H;��	פ�R�q�	_�G͉�J7+1,�uU������\O�	fc$��$������(�-�]��P��U�f���*d$HG�T4�����^�����>_�U��#�<G�=�%���T�?I
���ڳ� ��~B�m�}��N�,�B��i|��x�S��,����_�|��bEDl�B�t�4k�(�B(QY�������<��� ��v��H.��5�,�E��xb��iI�\7�=3�8�Fφ� ��Z���țe�w��)��NI�Ka�*�Q�ЂR%��Ք�����T���0�%���W�|AW��Q:��0� ����Xb]C:�+)"X����L��nx�d��O�ŀv��=f��^}�kוp�fe�f�.i5�R�Z��M��غN�t<E.I�A��������V��2�}�IE��ޘ9�2Ӗ���ʪh.�I���	ճqMR����r��E�ł����H`pTH'Ut�pJ�vq/ѝ�Ac�m��["�Tۡ�`nZ���'���Y��\N(��� 0r0��uޜn�89!�@���/!�mD>��5Y���(-.�F,���Fd�}�'8�HC0�k�?7�� �X7� ⦣���C�� L���̱'�Y�� c�"pe�_��!_��	��dˑ��$g���-�u�87-�'|��<1���szㇲ�d���K��0��!�9��B�.�y�l5 +J-��������&��ҦG&9����Éx�S�o�D��Ua�{�fmy�ddQ�]�I �aO��C� �E`��V5�D:�W�QQp:��
jX��"���gP``1��ܻ�+=�c1$L
j�`�p���PU��1��,ب�C�
���a�՞/�P��uC��
��#��$xP]'/�CbB�7�~�Z|o���g��c?:�+KG�`��o¥�-\>Kf̤ )�d�8�>=�Y�����_�
t��a�Ť�E���Ld��p�I�� �������9�	I�4˶�A�B���ۤE�A� �;��(R�Z4Ƃ�0.͡�?0-�h7,�t�h��0���BU7S�j���i
լ�.��S�jQ*�Ѷ�7 2!a�{�����\�{�A����f�6��l(u�d�wI(���{!ױR��:��~F�-0��q�;�(T�q�d��ӛ�)}ʄ ��T��0�� 0���ZԽ�Ɖ�� *��0"TA�a� ��"hf�~+�1��G�U�]���/�k����ϩ�U�R���A69X������Ja��"\1���x��P`�E�ƅ�(�³j�~D�`�)`�D�n���WPx��X.�Қ.U�`�X��:�T-F4�0���� ��4e���Zi����b�Vq)@�l�2E	���ʴ��(9�fG�w
�5�M/p
VR���ϒ=�la����s
Xp��e�*�!����],3�
؊t��\�	�[�� ��2=��S��-Z�5�F/Yf�P��%�K9G� �[��>娜L�/qU�v�o�e*��ӧ�+i�EX�	���P��-�шL���aAz�Diz�R�R4e�����P��q޻d��u����R����V���I�#Wmobȴ�`��C��wEs5i�����1�X���0�/∁���-|hi�Ԭ��d��1ťY�r��
�e��Aj65Cp�@�9l*r��tġ�w�#N%��7$�ܸ�� ��"��2��SR���J�6�/oAk���ӨV�Ȫ�����V��ܠ���F��vze�����%���U�+�^��),ӑ60ivO�X�s��\:y�����Ynt�������&V+�2�;���My'(��Z�넳r�?�(c�IdD6/4���
�7���-��7�(w|�*�&yM��<���b�uw��"QV!y�5<Y���5�R`��Uq�t�8
��\0n�q��P)�Ef"-����f~����k��=N<g�j�|�W�%�H����D� `"!� ǡ�U"�]za"�7� ���X]��K/�
L;pľ��;>Vy���JK���+V�!�,V�`���H��� �q0;_�e�,3�R���"�����,�t#һ�����-]�S0`K]&h��	������t�TZ��Ö=7�	w
J�����(��b�XvA���rO�+�10I�eK)�b��3K�x���ӊ�i���*���b��fgcG}E ��~�Ԍ[����R���$���9g�>..Y[l:e��1썂��(2�d�lt�R*�#�82�dۂռ�Ih<DF���t�n,,ɑ+Z�*X@rD�1� ��T��p̰�|/"�F|K=q$f�r�70�S��R���� R?"(X��C�|�� fp�tv2�8GB���P�4���~Ħ)0�z`e�	�y&��W>fE�E,�
�C{Y %��
t���-�o�{�4� ���'�kᦓ��Y��y��_:f����ch�|e��6�`��&�41T�MG���]�f_m�F�b�(2���%ea����m0��
;��2Y�$dĳ�3�\�1.Mʠ���b+�B���L"e1I260X��
fb��߿ �ҿI�*D^%nV����T��F��+@\A3�x��J���$�ae�M5l��r�r���GmZ¥�.-�%dP��W�H�%�T!b�F�c�Գxy8��P.���;!cG%?R�� /N ֌�E0�2�(\CMVk�Q�TC��zуo�4ˤ��}Rb�\+�9AmY�0�IJ
�G��!��ޥߠ�t�M/u*ًœ3J*��P���(�dFp�ԪYJfRi_c�Azj�� rԨ_v@0�M˔8g����p�"ĉMU<��_�>wY�����G� �ٚ�
6�\�1=n������Ĺ�w�0^l���R¢\�9��u��ܑ.<�0̛��X��6Q��>H8�FQmc5�����]P�k,��D�`�䀃K�B�VĴ[��@J��W$(V*�V�DH� �^h��C��� d�jb�j� ?h�Ed������:��H_�~5�l�� " x́���EP��ܪ!��'�"σbi���̶Cr��㵆�0Ԑ�t��������	r�,[��lL�[�����L�wԯ1�`x� ���������)��Է-�[a+�,�p�D9��*��M�U �	`Y��$尾r�2Bi��*�Ր5���h]W�����IJ���
�Z�p,1�WV�ꅻ��"T+<����+�1u.WwI��8�|KD�n�^��,Gt,;t��3�+�{��6C6*���(_��5f6�f&,����!wRˉL^e,<L�XM�1[R�lJ�p�Q�b5(H2�lL�̣	2���Z�Ȋ=�D3X�CL��q���G�2�;�/��hB��&Z±/�b*��m�ol��+��#����2ȩd��^.��t�e�Lsj�'p�ds���n�
���L&Xo�9�+����';�.�� f�M�U*� ku5��q���\�Vƥ��k��TW�Xʬ���m�q�.f"��c���3�QODv��sP𣋁m��\�Z��z�x(�y��!��(�	E>����yb�6ĈCc��0&VνB�5��>\)V�NȘZ�����Mt��5M����Xl�q,����x�݌�a�e�$q�w3J��F6�[�u@��J�i���1,��µ��ы�,�]"��� �!M�O�h��M�G���T�a`	(���/G�{ +�n�Ĭ��-�k����Ao$s����^Ȋ���W�$�ؽLj�c����}�z蜅hz�Je��ZWl�C��Q>��$�ω�Z<`���B\�`�% �L&s٩Z�&!��7�T�Q�4��3r�gO1�M�]�Rn>T��� x��-�7�,e�9�䎵��2D�R�]�8G
�^_p�O�����p�_���;%�����i�R��An��*-�����E�f�Eo�ų�|����P���G�`[���� ����rD6��Sq�7����r�����n��:��1�p���v��E�����19� ����� �#��߄�`�6��e姇��єd�tֺ_�R� y.�Fm�g>6~��$[0�U���&قR����p14wq�[a���r���2�_�VTT��;B5÷�3*�nP�${��F�Ċ��X���[ݰ�*L6���PeŸ��)1F�9j��ԡ�6�q\������R���ߊ����;R�ls�y��jX�g��T	l2X���Պ��P=L�X�$��]��6�8R�w15*"�bj������-ǴC/��ăU�ܡ1�S� /C��]+�u��b�
!��V��,��ṷ�(��n��P���S�lN.�	yeM�2J��Z��d�*bP�5ܷ�����-'a�2��#�[˘.�槥�CY�Q��]�W��e�<�਄4_�9�]�45V�K�8�����k�$&�2�o>�:�2J�Z������h��UKcM�_`����� �Z =R�ҭ�H�@,�������*�	��*F@�</��ݭs*�ȧ�ZM(6gr!KYc��Q]�w��V|��(n�Жd�kR��G#�'$uť�
�Q5��ާ�	���'�mp���
0��,u�j]��L���:� ������I��Po�!��lS<!7���l��B��nr'�����&X�Hb
�X�(�T�B��2Q�^#m�3%��]����e���)�Z���?��&��t�Y��X�4����D�5�?e�&�X��{��m�v��(�ᅋj�D��(<Y��KH�����z@O�	,��F�m��
j�%�9o�d�e����"7����-�a�_/:�6�� !"�i�8R�%D�%�c�7�.#�j��a���k��cx�t�bX"*���s6:~�byJ#��J�Wc��o{Լ�����B��c��5��DFF��J�~��;k�,�b�EM���0f�se�̟	R���+$lhVA��9 Jd�-�ih��L�P�Θ:�D���%����%E���%g��W�ĽW,�LV��@��B��dR�Y�q��2�6�#�A���7R���_)c���� �VLn:GZJ�m�$��AYq��Zh�Y��P�EJ�%+^eӐpʎ��^����[�.�b��.���������*��(��c\�թ�������S|�2�14�����X[1�����0������cl
#2٤��FI�P`�-����*��x�`n���b�K�\G�i�$�S=��2�=�Ԣj ^N�S0��`�	M7�*�v��}Ψ�]�;
aD��I�5',��}Fg������a�{c�C+��#q�K�ŬD��)D�2�H(K&��S������]8�s��є�߉�k�[��(M; ��[�S����L�L�*S����6P��[#��iF���4�CD�&�[���(s����]\叟D��\�F��~����}�0�w��j?�Q��a�	Q�\��=�<�qீb�L�t��%�TBFژ2���?e�K#>�;��q �C,"=b��q)&bo�(j|�����7e��}E�'h`�U��҅������a�� ����Ú�s�X��7�-Dؕ�F�.���0��(<�����5,t�ʡ�9��U�zwǆP��-�����c�	t�-5꓿1��k�қ d��S��\$09��^�kE��®TYy(�^�LA��R�Ӂ�"K���ʪ�QP����=FZ���5u/ 7Lo�r&֬c�+;��kS����J4X��ဓY9!R�M0�`�T���K��ܿ;"$�y�p��tL�a"�oFFgv&��+Gb扺�0A��*&0T1k��|I���a�$��B��W"� oi�FF(Ii�`�y����eR��;#�/��#���9��6h��Û���Z�YM������`�U�Y���nS��@�u)dY��7�8X�W¢�,��jLw�x�-���#q��� 0���Ǹ���b�߈]�]A�Co�ԗU@�35̛����݁^c�.Hu�b�Fl��0+ +Fz�r��|�A����3b+�]}M�l��,PS��"�oqf/[�r���T�UT�B�3g;i�0|.�Ք��z]�y�0�޺ch P�!>�P��d���X�Y�a(d�u9���ϙŨ���&��o�p�F�a#�_�L�ae���ad�(����A\q1��.9���JS��_�r�� �lzp�Q��EЧ;~��>kp������,��n�14`u��DZ��&m�%7p))Q� �P�˃� v;�%>ɱ5�E/�aݓ}��B���>�T���������,��P�Y�x_v�=.#֖T�&�����Y�V#Q�-#�=�Qqr��˥�KԨ�D7 B垅$�Q!���ʷ���u%�:.���<|]��1�Q��j(��u*R� ��AI^e��&�a�LT��q������ZE}̋��ĸd�8��]V�5V��1ZÙQE�2ο��4ȺؽKp���rC{x�)��R�;崶����4M��m��� ��382m�C���X6l]��/�t�eJ�5�j�$�@��G\M��Ġ���e���P86�!�R� ��j�$V���X�P&}���Zߑ�f���B��,�������WH�H-rr�
^u����r�|n!� ��Y��Sv�8WT^���n ��p���ZV<�hBŀXwn	 Z�+w �_d f ��@�r�Ȼj�7�}��	��eJ��1�D v�	Jy���T��O�2)�����bF˃�B`�(�g�R��O2�˔C���sdg�3��>"��-]Ե�Ss���˙p�\!,�Ľ*�ٙ����
�fn|mc�ŋ`Q��E"S��-UAجC�e�eX��Wn�z�#���9r�wi�@�j:jb))TG���Pf�wU�F�RPJ,�l=qP�;M����2`ÑkOѸ~�'|��?lE2�u��d@4\�y����)B��:��HV+k{��Oa��r5�!��U��+P�!9��CWC���J��"�[y%쌩��M��ĂE��%���^�/J���7xc�f �hD���W1�9O�Q�
{�����⎼��Ś�1���}�O�+8h؜�3�\�t�bn)�|>!�C��ELJ��+����@����p4P�� [�Pi>	�dqi�p̶�c^��J��㤌����/��$4����Y<%W���+yA���U�]�
�k6�K�XQ�*]؉��}�0�:l��"͘���bf��7񚥜j=�_1�k�ۛñ�1��ԛ��Ch�FU�H�{�aU�"��%fVF	p��X4s��P�-�\#���J�ߘ.��M��Q�]$�e�������u`5
�Sȏ���aE�k�}���<���k��/�~)F���H��2��"��B��%Sv���Zd��LV�8e[����%̅^w�!�<8S�*ʣ`i�	�swq�2���� Qy�����_3��6kQ)ji>����<$�{�.$psz�U�V�ikT��]���'���\3Z�Ea�`��B��p�KܬWX�&v'/{�.qu�H��s$���0��Z5�0A]2�e@�#��:��R�v̋����P��������2����< �Xv��b=��Q5)*W�Q=���&~�c_��T�J?���Z����@�
��e;f#��X9&+8�L��˖%�pm�R�}1�_T�Զ9ś�5S
�����\�$� ɇ2C6�$��E�	�kg���H�˥�%a-DU���:�Y��B6G����jnVD��=��էQ�(9� �����zʫ�`��#'��b-�Hg��d:U���{f��-KLc-2䄬6��sLi�+�L���R��s̮jc����L�Y�.at���P������'���8��\�vC7۪��2���`�g��ۗ*~���ִ���Pؖ����_��K���J��稝p��RPP�!�i�u��&�K�Al5}�uò6`U�^�NN\�DPk�:�_3d�؆P�1���v�1��̰�� �ӈ3�ԣ�Bz�ݗo$-B��I)��]�W��҂d����� ��n��7(/�&v����"a"{%��j�
``���UR,㇃��!�5M���^mM�Ō+=�A�dQ4E�%3D�������T��Q���5�iAA�0� ��B��؎l���;�.�ۘ��7�;t4��hĹ
�I���3)r��y5� �c�(ڍ|]���?"U(��F�r��\�,��u�@�Z,���)r�\2�%��/�I�i��pA(�Y�b�-�i�)Ӌ�*��q* (�D�X� �r�����pOYk�z����	�A��g��~m#� a/�U�nm?SB�\�!�T�o?�@���"���_oT�����g���h,ǆHx&9fyAi�w=SH=�/��8�e���h�0փ"�Ġ[��5���mW��Hf�>Iq:j��d��0$�D��YQ�ܹ�ޑ��x��)%����æ駞ez�	�Sc�Ps0�c$��b�c�1D���m��X�̃[a�1.(W+B�eSw� �*I��o�c*w����I�72�犽l�9[m����!eo�5��&,Crk҉i*M�T2�CR*&y|MR���@Ɍ}��|,a�1UƸ�,w.3�/pLXe ��Zm0���k�S-�������`�Ly����FiQ[����1�U��!n�#p�a�L�<�du�,ak�e�]���=�y��L��yb
��v�l����iK�qe`�[������+���ʀ$����U��~�����*��c"�r2���	���� �b�y� �f�f�� ?q��]�Ed�����?a\[l�@��HZ����7�)��OR�2^��y_���w:06����+XO0# M.��I��f��{9��10�D�X�3gO���rTfL�/}$�̤��y!L�g�2ƀ��%e4���n�S�e-]KljV�3pd�p��Q�����؋�,.f�T�@�\��%>Ƞ������~ٓzAR�D�0b+�oܓ蔇��^�}�d���e�)R��.;	�T�5JBT[81XYi榯�ܲ��L�a*\c��M�\~s
G\E��Ix����+)���x쉡�w
-�;�Hwp+i��8����^8��OR��*�����n���\1��X�hp��N�'0�l�w�D�����T`�a���0�35/��k�5�e�2L���0`e-�7,�� +:1�����2�oȟ䜅|b���g�Y��ASQx� ��%ԭ�1�X��S2��ϙQogCw��_Ss.�ǫ���-f���K(�u1�}����ߣ-����P4��_�!���uφ]��'Zx��M�ɀd.Υ_L0�9�r~�-o�E
�����Wu/��,75�=a�e"�D�Auq�.ސt�|A������P�c	r���"��_3
Lt�ԅ�c��_�Zu�4n��p��v����~3B<c%�1J)�!��Cq+WBP�7b��1e8E|5y��$%��f,i@�陎J���8R�3F㖛ĳcr��DV/�m�ʉ�ŵ�&�\��,hEB4�i�M�V�*�#�)169���?h�pM��ޣ�G� &�6BR1�I5��Ye̈JC7$Z\@@�'
#�a�? j�g�Z���D�
�E�l`�轜E����]V�%C%YS(��)��&�T����\�Op����Qit����z�Imb*������S.*gmx��,� �ncA�[WJ7uz�E�w.��A`�M9��q��6l���5̬�p<r&����jp�c= ��P(��ʂ�.zEI�3��ɼ��eWy{u	xzE�$�Gtj�� �^���&����LO�[�c+����t�PIʼ71U&�\����k
�oL��*��*3%�1ˊ]ҵdB/]M�i�-4���,��J��b_:�A8�ĺ�dF�|�4@�I�6c%L���y���b ��X,�1gQq3��ܹ�)����*HMD�,e��4�;G��A}'.� �,e;M���e�DS"Z_[�)�b-�}2͟K��!�o��Q��#�*p���U~O�f�2�`7�w7vu�9��G�r�����_i�ʺ�	�#�d�4j-�����M"y�N�H�Z�T�����~���o�
���܃p�$M����So���T�P�� �DAj!d ���!7���E��B_�#l��5*Z�+/ ����֎�EW3i�h�E���3�y<u�e����C,��*GQ�5M�&?��˲��ej,&~M��6��Vؘ1\��.��+̓~e�i�w<p�� �#-�ZKf�#��-F���9m�����7Q��e��[���FH���� T �(m�g̻��.�PE���im2�vٯPU��[�
D1�J��ؗgR�pPwC����D��ۨ�_�[K��sH����%��dh���%j\Ӳ/7�g���7�2tS�������?���<�c���x�����倃V��'ZN��faR֚�̳z�#��a�XKPQ.[VBہ�[ u��C'M1�^����C�#o�Y�~V��6�-��!�<;T� 9a;4���.e�
�0�5
j ���M�,>0�/� ��m���̽Hm������_�̖a얒h�3��C��Te�iq��j��:��4�3D���:��h��*��b#|.��,�0��;��4�Y/$�h9�:ّ�L��
X�.n\�*Bf*��:��b�Ɣ�ѹV�nx�H.�ZPښ.�P�-�2_�Z�Ij��.��v��4L��a�a�Y)� 
e��+9�@j<�U*�J�b��h�u���[ ���e�.։��KEuQ[A�yn��fV�:K���q�Vۿ�'�P��9�a������W��鋸�����%� �0��[���n�v��:Òa�٣=ͱ�U�b���m9�'���"�G��03Ua���;��1U�W�x���sS-�`8�L�H���(��s씪^78���E�xG����|.7�Z��O�>�PM+2o�u-�ng�,�׼���KB?��������L���c�b>�z���NQ�/Qe$�*���=#�ݗ6D�t���isw�����8ŋ2�zŨ��r�U�$|g��Y�c,��0R��w�Y�5.�s��m^bj�?Re&*j���x���6�.ȻFhrw0A\�����|*�%t�*`91*�Q'0K9����Rɪ�v��Yq�x����D;F�i�.K��Qp�z�����@�%�<JU��
��X���N��	B��"9ܼ�g���JnP�����zn?{���K�W� �;��ޘB�YA.27���[Z�TƕvZ���\ZK�<<$bѪ�����6���E&�w,�)��DY�k4�gKi,6�Ą�j2A�ɒ8/�b�
�� "���z�Q�9�i�%���%M�/� �$@Yk<��1��
|M�9���E����Lڦ����M��-���1�Ƅ�y������J���b�}q7��`��in�@73�����@P�D!r�D�r��50G)g��1!R��`�  
 q�~�k�t�%�\��� ���R6B�]MT�.+�fpT.�%L�3"੍�`QIK�72
��<����ł�2Xĕv��<���1z�l��)��K}gI����#��	� ��fYdҖ��!o~��wL�\4�q���!��>�
��p����N8��8�=�]��.c����t��dN��beJM�����Ț
��ʣ:��b.��O�V�O��)��⿀Ӿ"�����y",b"@-턒`=ý��� <��߅WU*ۛ��0�ڈ���qޤy��,L��b���X����c��ؿ�l�z�nq�6f��w�XO��E������7��l1<1X�8T��S�c6���B�_'#.?!,ʵ��K9�XVB��/����3�4�F8�P����b]jm�Qm���-!�a�QUƏ��.z�~�H���#��R���**/�y���� �� �zb4�,���o���6p���9��GG(@� #�F��/�&'4�܏��^	ei������.��.�@���FiI��mLupn)}��V�:솕����K7Va�)�R�B���B�_��)��D"PX������ sB�{�阮,��"#���YY���Q�l�ݱ��s�l<�Zu�S�x/���8�z��&0�2�3�f�BGk�T��0��a�ɩ����:�c7�s���0��5:9R�2�RF��
99��T
�����`L����(�8#�q���km 7x,6]@�+����KL��Y��-�i�/m�y@�A�����f�)��PP	O�4��R��Ƀm�$U���˩T�Hb��X�A��"�T���9*������=<J��3C\���fR�f
*�������CkHB�8)�]�)B+-�	T�k�*2cl
�짃�$��\��Ӳ����E���� �
�T��n�����.O7?����K��9�� �0X|D$ˏ��it�����ȧ���ćވ&��o�~�}�+�Qa�%���#���lǗ��£b1�s��-�{+tģ}�{ T��(���it�A��Z���*�?]F��1Y�K].U�1TѰ���h4v�q�*�Az;"�s	��(\�2�5-�-HLE-����%�ZE���f�D�0�U8��n B�|B¶98�n��$��E$|E��������y'���<E)�Y`�q�$���\��T�5�R�$-�1����+�\-��#�%��ag=^�����k9G�X���{�ǂG��C����� .�3��F�#j��)���+,Q��D@�Ě�z��3w���?%^�:Ng<��9�M��
�����*͛�WJUї��;A�"<� <��Z�%�=��>g0��it?'��c	�x|�o����#���:HI�Q���˓%]<K���B����a�)��r���}V��"Mʗw]��'r�Y������U��^�pƐC��3�t�;hg��4����g��[i ����6H�d�7�[+�ƍ\i��Lc
=D��KX��b���5.����45	L�Ŏ��`E�N�p�*���xfA����rK8���� ���Y��wH��T9��*��8`�6ʏP*���+���b��_Dr�M�ᆡ�S.�	�j�Jb�":��`�˿�7�f�c�qU��`��Pf����9�!1o$�B����%e��,U%*GNm�. آ3��ei�x,�?'�1���q{��U��8�?$i�;Dg�� �M�&�b\5bCX���՜� �.��e�q�P
eҥ��X�-*U��ߣSD'�T<CU���`�+C, qr�i��@�	��D�j-bg��� �J�5PQ1�6�����~��Sr�8�C��L
nǈ�Ai�#X��ۂ�[�]�Aq*^l��O�Iuz�8��awAD&�^6�+��9�7�e�;Y<7�1ʋ��X�1��{3��ò>��"j��KJpq��(츂�Ξﱆ�K������=�k�$T�1�]�{�c�a�=(w��hrK��k��vK����DI -r�`�t8�9��@�����U�,�Υ>�X �q�0�|M�q�����J�0����Z7Ip�Aa��!L���a���е)韸�S�I��-Ss"�3d֪-�*b-TF����On�JW~y�H�`jJKS[���"ʢ`^%�p]���%Ԭ1%�H��fY��웸�K%ܰ�ň��Z-T��� i�/I�[���U?$ �?&e5��1)����S����O�� �bi�]���0���;�+��#�r��*8s�zn
�P=�& F�,�� TviPF ����aу����!�á�ɿq#e��B	L�h��p��v~&���W"��׶.r�,PCm��՗��>�1��<�)
wh�=b�|E�����C�'1��ᘈ+� ����E��0��9���V���'�2�� �sM�R�t���E.7*���a?�19,Q�y�ܣ��y�ӶT� }bc
��H�<^U�TҦJI��	l���s�Qi�C�5��$��.q*''�dZ�>���q��f�DTp��dob�X�òjY�]a�2�)�c�Mi�'(���P�+Lݮ�8��i4�nN!j���:{)�Ȕ�\d�t�C���9&��Ay�&7�������JS����q+��ط��U�W1fn�;������3^�ӔP���e�A�sAE㋁U��K֬O!�La���/�E�H0�=qܨ�<G_�7��wr��e�'�Ļy��������W7�E�uJ�p���2�6H���Q���|YH�qi��_���(B�8y%ڭ���8ߟ�XJh�� �R��aJ�5q'��Y���i_�Q�6T	��'�+� S{1�*�i�p@��1NIyC q`���DЕQ"t�7�+).��p�+�k�7�{�VF�o�D������~�@�Mfa��ƙ��T�&�%.����I�Ň{�&%��/��S�7@��>{��nxܦ,j��i����0ik�p��KwCX�@�)f"��@��-� puJ�7����������fU;l�
o��Q�n�w��-}�~����.`��1��q��m��20�"1��#�;��_��Da;���GkXCDK�wI�EY�	Zī�SCI���e��h�9#���:��s�o�jnK+����7����NV%��F�9���|s +ej�;�>�HY� @�@��P�.�����'ɨyw�vWF�B���h,Òr�r@�eY�Wu��z��upB�DiIvC�lTW�@
�lX�/Gq(E��b����J�b-�
�#R�m*ߖ�m�3UA.�Je�X�N�FV����v?�j�xp���ĥ	�&y��C3 �i�^��V�c�z�rxe��G�cmyܥ��u���q��l��P��0�XBoL�����d���[�R��,yFt��+.
���Y2���,@x���G�������#��y���ل"�ܬ-�R=��.Q�I��|�b#�a��̂����9!�?�xA�[E���&  "��8�ȍ�Q.����ƥ��� Zվ���s?V'�]�F����+�A�1�ӾH/X��p��s���Eܤo��d� f�|,�\!)l�L���R��2#�W2 ��V��
QD ��c�0]$�EoR�b�.�Z�G0�fxܮ��YD�-J���,[$)Y\K&�����.��	~�K�b�.L��;��j2���7��i`�3��ҙb�B��"��:Sqz�0C�����r��Ux�390:�QЖS�v1R�߫���{P.�q�`4�W*����˫o�˹wȅ>b���0�͟�%/����2�ExMЏ]�q�'� �z�o3?q/���?*�M�.c��ͦ�����n|=�d�L���c�k�I���'��;�VnY��'|/��-)D��c��6s(]�>�т�A��6��u,�f!C�"�j��-�@6��Y�ĭE�anD 9� MfAbp��`��q䚉|�6��s�q�-!���bc2�&�A�iL�1Q�^�b�n�JD��z���]�EY��d5C�6�CEp��x��Ln����Hu�m9|�,)\��"/�`e��C'g+:���5 �(��Th�h�q��`K�rx�⑒�ˋk��pʰ�0�R�[|���Lw�\��c-�.�y|
��s�E�^�Y��C�Y|uu$�5����д��� ����l��p˿�A*_&��E��s�����L�;���&-m�����Żfy B�|�l�JQ�(Y���Ř�����j
K�u���D��[�2�t���r�kx�&[��L��]�khiQ/�����>�RS�a�f���Sl��Q�C�q��d+�YI���Oe�֠�c:>���Ҙ��q1.\#FXm�nv>�qU�$m�Z�l`�n��S�mb����ukO=��9ŐT�s`r��i���/T�R��u������.`k�]��`�p�L��O�4 ��T�31Պ�ȋ��f��E�0|	<����%͕�@|Hli�M��EL,� �~:���o�b=�TE^�Ife���ƙ_�b �p�VaĆ�J���0@(̞W��LX�0��K�+ɤ�h����P�Φ���$�t�7gb}ˤ��[Q۷���,ʃ��TF��NZ��f�*�Q���r�q��Yq�CNI�\U������ڦ9qV�5dY��ˈm��j5U�4���y" �D�Gܱ�İ#����l�d�{�j�q��C�n��O0O2�*����I�1R��Q�d>��֬ �PL���(Ӹb8��� �dx����>`�Y(���5ʓ���W� �أfG��ȤVj��n�==�%�Gq2�aFo]]\!o��`���	\��DT�F���(h>��1M��W��'�ṲlJ	(�'�)���~'��
��?8��evawp�|�PP�fl0=�+� ��\O��H.��Y��8��h�[�xvL�!�٥� �F�Y��:��28J�,�[(nQ�����Aw*T�*�F(�5c�8�bP�̰�$���P�^Q"7�D,Ʋ0̡��Ta�q4֢]
jo�n�(��ߊa����.�����X�c�D^n&��y%��P���J�3�K��������	�#���c_��H㉎�� ��QЙ�Il���Hj]��H/�~H �%�P9�3Z�#�zeb�ʿ��ǩbէ�&1��"l9�]�tV��5��e�d���3��nA�����+K����y��]�
0���t�%�.?1�.?$���?G�`�QK��1������X7�3vf�T�(��2�k�UeO�iC�.A����w� ��dL"x��r��4�t��_�:�dsn����]���ȏ��uQ=�l\$W^��#ln>�%��t���+Q�eBÿ�[1��]ʰCr�H��ZY���5���ab�
��RU`@���7L[�kW �_6�V�\��vDQ#�h����*��(�M�Gi-C!ܬs��E���d�Y"�^�R[-+|p�dƨW�FG��Ú�S�]��T�چy|p̽���d *^k�M*!3Cw�m��b_k����iO�o.\q��C��PB�FV��!E��(ή[�|l��͡��.YE|^؛Ώ�9#�r�+>,��T��K��%�$4��� 	Y��%���3*�r��PL�O�Qc,!�%>IECj���1�J��hT$2�Xܭ�L�9��]>��J�M��
c	DRة��)�5cEښ�e���,��"�њ�h�\XEh� p�)H�����Ȼq@�k�ٍ&5PT�4S5Z�����J���pT�Z��� ����K:�����ʊ?Q̔Y�,z�؊��MF�&|�h�#�����XC�V��9\[,��HK�-Q}Djj^�q-#T#< ��;5�12L-�m�Z���|g�v=�l�v;��C[��j`ҜeC�"P�G��5 Ӆ���r�ְ~�՚_��c�;#J5s���.����jhf҅��, ��.Iue'��(�<����z�7K��e|G��O�T�_������.����d�0X���1��)x�e�L�%z3��-��AgJV	�jUo�á��!�9��:�^2������:�ŏ2���Aun�JS�d3�~��!Ĺ
cdT86vd����dPH��1"8ȕG'TB�Q���0C�f��}O�>��	ܲ8U���]���N2[�V1r/d
�/d���Cx\�.-�i\>��.c��{��rSA�Z�+V�m����?�(+�1�v�.�x�)�p�UE�ơ.��*���p�)r�M��b��NU�#ko&b��:FQ�8sn]@j�D%g�ZF�@��kP#��5����p�~�j߂,��RL[��b�,E�Vɽ-@��9��.ԉSB1#`31��rGb^�f�'�D��I�Ĳ�|f�FR|z�,�ե��A��u7a+������X�F���
�)3,�(�j	����l`��$�fk �K*
CC�����F��+	�D�B����b�o���Ҙ�kXܡ�c"b.H6K�0�MwU�sYr��#�*��B�0��ZB��]�	z�9/���G�&�G�d�o�& �C�&V�k��*+�����d���."�|1�"h��u�*h�M����:��	�wR�)�L�������;�T�į��ٯ{ZV�Bv#�����M�j!��n�UQ,e��ʁ*['h�J�>)l�p�cX0*�12b2��t��6��C��������L�wQ2&(/Q������0�-F+��q���f�9#�_��&��F��
�|��j�	[�Q�q貒����?V4�����&=,�ǘ���0�T���P�8���P��",�H���1��ɥiS/�p��)Y�T�XDV�ܫ�2��P�d�ĆF����k����D��\Њ�'r��REC�fm%��,I���>4n�%z��{�*��R�?UJ���1?�a�8Zg$�\ g���
�����oK��%8e���2�E�o�V�h���L��R�$n�*4,�c�$�F�P������y����&��es�2�/� ��&d ��(�2�:`�1�C�:����K,!WQ����[g��%w`��I��!�")4��� �P��̻_�ٸ��3�y�Y��+̶�$9������  �	R��3'd���pDoT�C�c�'���Y�2�X�$��G���ԣdR�!�G�+:�<��]�$�6�i���.7E�/M��4�m��e	E̤��� LR�`��}��!+�eQ/����2�qaNe/�*>0�!���d7���[*W�k��� |��R��5і��#R8�.;AAܱ�TT���v,$��a���T��D��:� &x`�h楰�� 2�\���7��+��cݍ
���Mcf� �B�㜥�Nb) :��}�����ipf��vT"1��
틐��ށ(�X�{􊅯%B6��&
� 5�KZ�H	��	/Q(�fh���k��i�c�~�ej��C�
U��H$+�YA\P�Q"�G\��PT0i���� ��)�H٨�.6X�J(e�Å����k���ѫ�)�7(���
}JF���h2#8�F�<s(�h7��Ԣ�}�f��`������ĵ�.�rJFͻͶK8��j�J~�~���������,l��-'���:����G��&�j2��7�H��je*w�?D���2e�@PKS)QK3ľY�����E.8K�L�B�lb@�+l̲���V�?�*Ш�� �b���&C�Q�YB��bT��chD����d�<*�6-�g}����q���A��q�����,��F�M�	n6�LXdM��\^��^�r��B�\W���9|'�K�EAR�O��d����`�,+]��Ka���4�+MU7�
$�14@4"/�< Pk���eԺ��[���g�qi�EG�J����ҟ����E[�1�JT1���J�
�(a!�8�b6�"%V%�")�\�LQi�vL��M9���*�1QD�憥�men�jQXhn� =�4�� 6�Q�V�t����f�p|/d�g	�h\���
ǥ��F-�a5aȸ��%�K���s!!��4ޥw2�xR�fj�?p<Ū���,��"�(L�PR$!���KLzKa��z&">���F�5]ǰ�v/����DJ�j6��������R�uQaV�£`�TU�-CV.R��W�3s�hib>��*���� ���$
u\�,p��Ԗ�@��H۩^P�lī(4-�8�ee�`��*黀�6)��Wsb�d���Y�ޡ8��c�P�uKLP�^%����F5;v�&j�
��FG����pf�Yuj�W����ҥ��P�$�M��:	z��N*�av^6#i�9��2�"&2�"��[�t,E~S̢z�X�+�Z�E\�P�LB,n� ���H�od���I
�sČ�%r���.��^`�Ho4���@i6���aE㹂UXt�Qe�[�Ua9����Qr��u2�0?E1eؗ	��M���ţ�؛""���ŶK��I���	v*.gH?��L��R���_K
����Dg�8�,�X�(�JA*D�	D��΄�`a˦5�|d���:�؄� 夣���#��a�K��cQ,HYp��/`��6/��X�f�:�*��@��+�"#d�u�j�@~xj�i9�6��e�a��}Kk15c5.����1��C� F�2x��� #<T�ݘjV�e��=!���ו-�5w��2�cTJT�:̆.7Z#�WWÀ�Pu2 � X��pCO��62$���JF�Pc���2l]*Le	��˨6m&�KbV<��@�-*'T�h��H��DB)�I��pz6�x��	�`?pܓ
�"� P^)��ժ���gԨb�����m�K���(5��N�,e9�s�#���FI���=0�%��HF�OQ��b�M���@�*�sBt�jpN 9�����-`���P�U�a���.y%�p[��(����P�-�lo��*P��i{�-0��`I�����$�#��b13\�r��H*�e���o2�jG"����y A� %Z�d��� *o!,j�a�\	A:
Dծb��
>�T��!����C ��)Ķ�@������R�oS�½� \���7��3��G��R��3
b!`j����n\Յ��@�S\X��PkdW	F�a��
����!acB���P0Rm��f��0}5>�m%�:�8k.�	� �W�Q]�LA
�����@1��(��g��Qz�'���Z=J����	��ٿK�\��+���H��g����"�=��^��C/��޲]F��$�9��]���p7n��
���T$).K�oO�"��`��!Y��	so2ѬV���8� ��,Gbi�.<��0�B�n�LE����I�}�-PBwCD�Tϲ��Hj�&��L�]�F3Bb5������F�� T61%q� *͑�ȏz��IR�(��s	R c&B5VF�0��e�JX]A�&�E�B?�(��o*�ɰ'��[�0S� �������s5���-4�Z�Q.�֥�=& ����`���0!��{���Bq������K]�������x�*�2ùma���Z*��Q��Bw�m��^��׉�E��� �U���������u�ɮ�������|%�Q�{c)m�1AA�L���C�'��50*�5� `xuò���H�z~���c2P�s�\��⭗bs����dg�Y�Q'5��E6
��,*/�,uOH��U0h�OVK*��K�D��"�6q)t�Ħ�Mg��вg=� �*�`�-�
*���+4�:���w%(�q�2	ȸ�N�q�C�@މ���}�29�o�%�6��Nx����fk���5*����л�us�Ќ�ib�i����R&g	)|;M��6�_ C�7 ��0���f��4����a�ܽM7��R����d/�ej�,�.���*0M;�9�9�6%��3����?��f �%Չޏ��5���k�U7�ET�A�f��.��f����X
F/��t�d�Y��o�qǲ���Z�*�'qQhi�� �����*"Q|�]JU:�՗��,����Eͺ�1�'˅������e��D�8���Ȩ��*�F"2Y�>��UF��q$ k�H��BgB��Pt+�7P�qU.�sL�	+jS���?���9B���(��*����$VR
�(n�J$0�<���8C�I�i�)��通ں5�G�ކ�kI�t�̵t���)%t�c�x\[f+P�w��Y��6凅�N0����n��|%�5��@���8�!l&�� B�ܤ//0���2��̶.���3�� ø|)���V���.Yqʢ���0|D��a���p�@2� s�d�U/��W�ˈu�8}�\r-�/	e>�V�;2����T%��c<�)�!���1gEE�^��"j�	f]C�C�s	.���ϖ�6n"�}DR��uB)[\��fs�0�㚌2��q(�6J�j��u���h&�lqH�P;�����Ӯ�z^M�CZ8�x�/&�圄C��Lat�0��\���F�tW3�.b����@"pM� y��Z��,��?R�}7`,�W��
Y�� �Y� ��`Mā�r��7�p[�k�GU�O5T=ff����Y�ڣ�~���a�p�Pm/��Q8�<�(p�ў��!H��R�.�ʩb*�T!h��E8�~�Tr�i��{^�$6c02w �C��n�ѳ��H��O�m2ԳDj4;�h�bȏ�Br���ijè7\�l*Z�zZYWKl'����!�(�qًʜ��Ɩ�r���ե�̎3���j5����S��MC`��� iX9�(�7�c�"͝u�!$TU�Od+E��5%����מl��lf��YHN[�H��j0��Ղ�
�ch?$`�-Î�p�$v��W����5>�9��A� �(�.���K��ߺ$�:� �l|mIb��M�	[��!^c���!�m>u	�D�n��qC�CҲ`�Z�P����ܮAd�-Ժ������5e�Q>t��}�8=3JٟaXCfb?���0�`.0�Ķ�%�5e�X��U�OB\@^��]z��o��L� \�WGj-�'YV��ȅ����4U�`�P�S�C�jۄوtqI���1	�5�-������jO��r�48�4�o�Q4X���A��?�P��� ԡ��W��)�Za��ղ=A�Қ�qx�/wA��mv��RE���M���<�eQ�K�Vd���&`��1꫙�Z�l~���O�Qtk���-�
�B����̧!+�?�T�h
��b�y"����s�B{���h­�%���$J�^�Y�UIl��1pWr�PN����� M�s�j�Ƞ�1��Ps[!t�aQnX��+Eĥ`��wu(��aN��v2ᅷ�[I��Ljc�m�o����"2KW�p�k�V5�岭�K�����F�X�f�$xB���8pI@�%Z�&�s�	l1ޣMH�] �X��Y��+G�QЮ��T򿺆�4�&�^����0fѰ,c+����*0UT�p�`vJc�B�t�����`m��\L�c�P����"l�?%�h�Ĳ�S5*W3(�'{�%��A����5���� #5���Up i3�rTC�+��*��tY��4��^�~`צ�!��،��"U��):T�ʸ#6�&21.>0Ù�ғK����_��G �.eOq���EV���e^�9�spR�1M�5`�V%NF4�Q�s����AN�Op=���=j[�rf�Jm6ZZ�f�Km�}_�m2ܐ���H1iK�/�*��������-��4!����c* ^Ւ�ȣݧ��NGC�!�!Щc�.-���H�)���<��=�A�е� [Һ��.]�x%��3u�XO���Տ�D��p[�AG�QI� �*����3d��%�"KF���qPÆXXq鈋��@.XM`3w��'@-d�h5[��܈��؝F&1�$ٯ=U���3�ͽ� ��G��pZ4M�ˮ����+u��vQ�&x�!�6,������Rz�ʌ�t0����
�$�!��4���@&b�aܘ*�F�3�8�CT����n��MF�WM����X�� N��-�:��4ӓv��n��)�b�M;2V�`д�����T��7l-�����b�ց����ف�J�/v3���yUrW�v�)�;�hAKpΈ�*A`��!Ս�*İ�hBc���R�]A�EڪwD��˂h�l�B�C8B�r������ ����C/R�)�}q�Q���!��h�����j�o��6�!�g��/;%%sh��G�/��$}dQ �v�삭���\��˞��-�b5�n	��Y�ah��.1�\p��D��H���mN��nً�\�Z� 0�o��[8�\<@���`�/$+�X��U2�| R7�|�ıi�����c�az0�Lj��'g�;>���j�����9�L�H�}T��e�#L��tp}���8KA����N!g�R��$>{,rJ��e#���0B��l�k���e�H�.S��q�s*��R6�ְ�>�[��.R�~����7��Õ��J�mh��*�od��*V5ME�ަP1�1�>��f��%��1^U����)u�Z]S��f��u\����.TP��(��V�ª�Cd�^� �[�D�ØK
�eM�eY����Vf�"/��x[�׈�Q)��E��b�3d��Ӥ�?�{����!W��ޘ�p�]ˢ���3����!*�2��6OڝX����]�[��	�:8��� �C ��L��ei@]���֠]��^����%���h^yu\uSI�ɞ�*@�Lt��Ae<�rY-�˥S�f\��.@ǀ%�b4�ܣ��Y�o���X�p�j�!�^Q�� �s���� �xĠ���2;� v��!� �c@��� _�������b����J��[i�hjĿ�:�H(�u�õ�u2!W�`�x[d��U���d�:�l��Lkf`.a���0 f�P*Z>����t\ �o�
J�L
#�bg���֥̅攻�����P�܈ڕ�0����bf�m ��d��9ص��F�vCV��T2�Q���ђ(���$��eVg(�k��RZ��B�Do��~Y���+�p>�EF�λ�x�nd1���:�m�r�P�O�2��K���#QȈEk�k��pv}��XS���(�-~����!�@j;���_�s��0Bi�lO�J�0P#Ún�bk ny�w���Cz?QB��s��+1R�a�4�`eZ��0@��T��w1i�����{������.:��u�צ�K#a]jSqe2��:(���<��B�p�sV�X�"�s~%4��i����<>��5����!Σi�Z�6q	n�X�',�����1�rJذ���X'\�u-~'�pAn�QYRWc�J��Pi���@�a��2��~�.>#	|N�0Q�.��=Dz�A����X��2�X����UeO"2��!�ƚ���H��ۡ�@�*Yiay��l�a�� ���$�F��0�ܮ�Vo� (��*p�$f
e�[`�˺M�ǫ��~�n'�A�qt.�ku*�K, �,�]K�_�\������ �5(q)Y��ъ�$��02��K�I����&���(4������y"J���/�R�E\FC��`���,s�2�F�Lz�ce�f��;�9�l-M2�ne�U�L��)n���S$]�B�$:/w0$Z��G!O2ܘ��~����E
�*-ya(@�y��s傇�v���3^�B�
~�)�Q�	�-Z��`)wbW`?�T��uU%�%̣��F«3q8B��� �bS퍱T�F�	�+M@k�Ʋ�]���s��T�s�=_C�}����5�5}��u�jb�$N]�DE�9����){����`�����U;l*�J��0����{]��䪸�/�M�\3R���̈́G"Rq,��K1".���@ln+�dbX�Xd���Q7)�ٔ@j9v���^l�q�)��1G,� b�ݏ�f>��XQ[�����o,X�6�e6X��X�GQ#���"�<����A<��1�HȊ�1[��m��Y�yo2��pm��+/���$�z�e���]�2�Uĳ��ᖤ���ťnv9`ED������*���������S"U�U�߈����H�I����o�:JW-��Q��hu�d��9��{���\�J8� b�9@aI�s�.�hS�peV$A�0
~����L�Abu�Ļ/SNBXe�!��Yk �SMT�he]�Ti�Z4H�}�َw0�:�*�ZL�a��=Z��6�f'0�Gl�1��X��檠�>K�l�G$%m�T:q��ʏ��`��Ρ�H���V�f��#gqqHQ��7԰yF��d�pu�<�%����E[ K�������6D���솳�p��e�8�*F��Dφ,������:�%�'q����38e�7���#diE�����~�րg��n0v���?�*�kr��(6N��Mī�60ט��F`D-1OPDs�.e�6B%�2�'���<Xr0XR�%�X|K"Ά���e)���F��z/������!WBs}sm�J#��H*���:G�m�PߢR��j8*��f*���T�VBZ���>�#��[b�'�ҟ=ͯ��Hqpi苁�Bk�i�Z��-dbA.���ʓMh��l���`z ���F��H������&��J��-.�n)�%��u����0>Ь8������g"�g��Cqc#��o�-��{%�2��4��O|�_��TQ4k����R#K
���#�N�/�*�r�^��ux��ӈ�Cr����ᖪ�B���s%�E��F�p��PU�F������B�	��QM�	Yxu�-�\�a�d#-�+��z�����Ah�����=.�9�G��065�˱]��J�͑T)2�B��p��-�4�:�@}�Pبled�K"��g\�7�)TT�3�}�3�s	.�K��t��G�LW�H�Ӊ�5L�Uk-l���F[;�5�pw8!�[[H���QS<-�.�	�"J�G���h�����Z%����]ʥ�ԡ�e@���D���%�0�ōJfo�5D�v��G�+���(����z��  4��s1(��w�Q%eD�<�_�v���a#A�E`�2�ٖ�h�!^����_��Q���Yk�ԬP��]$���.�F��J<uFe�LZmy�ә�
z����)8k�
Է�Ⱦ`�=��L���U�B) ø�^Ip�����빑\\�2��e��������p ��Fl9Xtm���g~m�e[���'G�[&-�{�R�G�}�b�]�<��59
�9���H>��p�X1|9�e��7�L�0\I �0�&��V�������(���0�n����Ɩ� ���� Ip�po����Fp�`j{�}�Q�9ewlN�Nn�W^�����U�OĨ�[�"V��3]��EVD4>�#�4���O�(,]�d��r�t���1-a
B�w�e�ʟy�DX�ͷk��\/�r�e(��jK�Q����kY��t�w����n�V�B�b��W���I�v�QZ��[Mĥ��Tt%j�2����&�=����F"�gWZP���O��m&��v�I����q�x�h4��Ǚ�I�	� 7p�5o�x��B�G�"�K��p��e�w����M�<�f�Z�s�������` W�t>���1E�R��Ԭ������`��f#gqk��3b��jf-u�JH���WىI-:�
����vb�����4۫�j!�!��eeV��]Y�o�>Ad�pnU�j�栀4S�K�1�3p�b�A����xal=�(�Cu+�]E7�K	`�p����J�Go��̹R%�X�W�W��j�Zaf�G<�L��̿�*���GH�K{�5(7y�;uC,�1C�cM�A20{Q
�|�ݗ�������*W=�C(���\�=����R����^p�>��̹\�ʩK"��e���<�V��݈��ΡU�Mtʋa`P�q.�ר���o����Gt�E5�L�#�P�F~���z7���UR�g��X���L�چi�l5�,�ja�-�+3���۬[o�M�*��;a�U���b,�b�+�ٕj+��q�X���F'�L�j$�UlȇtV2�3Z"��tk�<��B�Щ�R�*���0��cpl��M�����!�"YJ<����Yv���P�d*�W*���>��� ���.���6s,qY`��'%�J����d�\K�4��6�I��*,��]CU�#'¯�AE�}��ק�C!�QA��R�b�A0�VV	�����SL�%T�퐃�.Y��%ڊJF��}w��5�\}�J�A��kz�tQ,�q$��e���p^��Y���]2~Ё�.�N݉��R�)J��a���`E�j
#=�`��Vp���x ��-ִ5�<�Q���#歌t¦�;��Or�x"]@*F��cn~#�m0^ �f�×<�f���A�L��%JQY+n�#�۞�K]g��տ 0ʨ��P!�"�D��T�'��7���,+I�]��� /\��_-DB���� (UD�,� ��K�˟�0���^J���,������ZL�L��j7�l[|D�b���gn���A�W$
u
m�E*WpQ��R���h�H;�R����\��P��ވG�ƥ�%J�]b!Ǫl�Me���$�zb"��
0�����?��J�#|{{�r7��/Aw�w���4{��m�a&F(�Ī�2�s~�U�����$E]�s�J@�vA��a(�Z�%6����r%-�:�!����}T{��4��U�N$NP)�d��e�0T)� \C"�c��O[��Ѻ�h��`���Q��Z.��b
�@4�̲܈C�+������2F+S�1U<0,���OP@m�"r�J��.k�z�Y���@�_����L��9x��X���^DuC_�]<�"0莴�byV s|��6�^Is�상۾���(b:�3nH77����\ae�V�C�uĥ'2�b��P!k.rkw)W
��U�`���J��S
�	�e`}�V�1�����5��c8��}͊����bU��p���"���P���L���%kHט����J|��0JҬN"%�2��63��̒�
E���yJ-��j1é�$)ɴ?�-�Ԩ�R��x�g��-�⢅]�^!��El��Z�H��Z)bP�W�������Y��ҚT,�Ol�xY�f4_��<i4�ś��R�i��1����f�̩Dt[����E��0�>�F Ļ� 5��0�����ңSQ���d+�Bv�K���zf%�3@䌒Ѷ+���,Ŋ {�=Ъ��W�͠F�}� ��	�o2 W����8����\����DM�Ii1�߈��1N�
#��,�T{�%�d���ň�2,�@A�-x��P�e �u*�O$ۇ!1�ljHi%B�ʖ�>�r<��L�uo��F k��k�Md.����<���;m�l��WP�Q�̸�$@g�B̼�
�C�X��FZ���j���U,�����_��O�4o�^� R��� N�~ܪ� T��C- �3���.of24r&I�m֤ZLu��#���u�T((���Q�.pUĂ�1�(a�r^F�[�:�PG1`P�3��Qt���bY#\�d��� ,p�J̗�����bg
1i\c�ܭeY�@Gg1m�i���d�"%�B��tzOf�^ t�{�h���`!�\a���0�)x�V<R��6b�L��&TX���~7��!�����'�F0�|�K8�Eڛ�2�$���Gj����2K�S���n�����*�*KR�R��F�����FՆ$��V���tP,�J���P��3T��_���&�<奚e.��Ӓ+	Lٖ�9������5�~�E�s/�\c���du,��.*R�����Ddp�
=ܳ���?R$�_}��s��p���,�������G1G��ۉ%y���L�-�F,��p�f�u�]}���Q��-��?�+I^Ǆi�̜��2���o�)��r��x��!��T��x��G=�o��zOJ"!w�]A7���9���Q�*9�����Vs�=��?S*��!���z�����Y�u�DAa(YG�����W|\(����_�_����:� �����f�s��\Į�%���*�Y�*�K4Aa���1-VZ�q�p��
ۿ�/����p�6��`B�j]�ս2Y��Xq,�d�0��{��� y�$[����11MT`;�y��k���o�&�I�Ga�G���
�@� *Nf`$�o�]�M-�g�q�L�҈�6Gp�E�Rc{�~�zB���Ӏ�I`���G����se�Ħo2�B��ȥ2��cqI|�,������1�,u	ΘA��!�� ���F�����1U���b�d�� �i �nx1@Q��E�Tݢ.f��V����7��v�q�!���&�(Q��1K5�^w��K��:�ĩE,���̫��tQ�I���C�o�0�L�$~�����
� ?ф~�?��G�c
Gh�j�f�����p�QW�2]@	l�s(W3��Je���Yq�����,N w�P6�Z�4;��D��KX#C�"�L ���3o�d����J9e��b�p�����Tq��U���	_#��5��px�N�K��aK�o����0�|��fl�#�6��Q�dw~�#0���`#4�pS[%�2�H�����e�q)b�־���k�{� ��/̻WQWX�������)����_�:[���.+_Q�+�c�K9�F���V{ac"����1Y��N���ovwJ��@��=��h���(�$n�U�d�y�\n)t�GW��	k��h�Ix_��0H�.�)vp��� ��T<JBEp�5�\��R�Y�bЎ��%R���F�3)Z.���z1_r�dy�	E�Vֹ�w�S��&Ǒ�ܕ�"q�#�d%���c2@��L�C8t�W�`�WQ=�_r�)��y�f\�	C�]�,n]�`� �
�,R���b���#5n{�mT����Z���ه�����&T���l�+l��� �� &�Ks�ܧ��PŊ��{$�x��!C�.Wp銸R��H�u���b��q)4�W@� C�%5��Rz�:�]E0�B���}�˃B;�J�h��4�~�ġ	@���e��	��J7t���(��1�!��/$�vj���.�9+!٤|�!mUw�x�LE��à�XѮMY5��xJh��b�Îffk�xܵ#�0�S�\"�:�*2�)�J��u+������Ť�fk�n:�������}��8����YXe���a�����������̌n����A՘X��,<�C=����Y?PR��uf�W�}&<Hk�J�bz� ��n�0,A�7,�%-	æ
l�$h.��K0� ���m�^�e4FQ�el��R�J�\0���C��	����u#4�l$��B�F���
m���+���p��6V���C
�b+:�`�ӯ̶/:�B:$
�R�1`U��E��VҊL4��.����Hi�/1[���ʢr��_�Fk�fmn�ࠧ×�Q��E��^KRu}0E���0�X�ӄQ����Ih�0��|5��o��ZX��$:�ń�����	U@hJ_��`���E��жD���bBa����TpĪ�1���0D>�N�.�U��\K��Cz:��O-ڷ�)HD%���6��K|��[Gp�9/S�
�p��Ї8M4��J�i�3�p�),R�Ϧ%�mW*<��g�<���+8p���dk��pla���S����<��c�%�.���z![{�� c�u�Fd50�%}���Aچΐ����ݔCҬx��Ȁ\A������;��?{7"QӅ�ƌSHW4AN�����e�A�`�O�T,�n��9c��E�ck>��*�~�d�j?h��X�-�����Vw,��
�s���\Z�W�(m�
a]y�-[�ӄ�>��A�1P�E�c0�w.dce��q`���o�%�� $���7ŝ���nt�M!��#���Y2���&��­��R��{�% �`�RYy�\�LǙQ?2����ȊIg�6B��Pf�v��}͇;#�`.	w\����@.-B��5nQ�ǝ�Cԭ+,ja7�
�N�Tt1�>��>e މێ�v5�C�k��{Gop��/�i�Z*��^�g9�J�uqY�=08Ԡf83xh�4�y����-6`�٘�32f^�����Rɞ�Ul�-T��2G����ط����A�����=�҇��[A�Z*�t�A]��.��1��%����fR�� n5Z�W��M��&��\u���f8�������{�����+�ؚ�^�����:b��cl��6+C.�`}�˙���8��C�zJ�)WT�����v0�Og��IʔO̗��O�<� ��h�n̒��s��hp<12\ L��-%$�o���%��<�Y�V;�>��+����s	Ʒ�����G�1�[q��{9��P�4�N��*�P��LQ���W�	R��y�E�l��W��lg�a�
�P| �B=�����2],t�Vĳy�c+��)P��*�`���q�K�$V4�x���# ����V��1-f+%��`�g����3X��*�,  �2D��_L2ݒ��
��K�$�.LJ��w��yGQ:e-����Έ�g�AT�\)�d?�0�ۉU}��S҂a#@���s���V/��R-aC�0dLP��Oy؆ݙ�x��A�F��s��8�ֈ
�`;j))𿀇I���/�$�=�G�ïB(��S0��M����d�O	i�R�<DU��z��l��Ä�� �t�+C����b2�R�F�2�@	bh�'�}QKF��(������q+L+�ew.�?� r�\]4�"������RmTP}�r� ��>��Ee��2�@�����|ˁPI_�d2X��������-���b�r���$;�iXj�#����*U~�6������I��"m?R+�}wJ&Y�=�
6����+�E���Z�*�����N��"����[�:A�h7���1Q��u�V�R�ɐE	��]l�,R���J�.4���J#�Ւ�y���e����by�g��+�w*Cx�P2�\b��i� 6g���M.Q�4�����Ɂ�� >%�:DHj����]^�@�.�Nv�ba�l��b������ŋ��Zj�}�`
 �
��K�!N2"A����4�~�pB�����%[B�es���8!�?��a@e0H���k3Z�Z��A���'e2���fv�s1"dl��-䀩�hs��1s5P�B[n\�u�x��s��\��n������ K���{��dg݈��҇�6���:���t��D��)�;L���c?5����V\���	��%�4a�A��C�%$�_�H��Ku\	�
�*)D{�h:S����&��� V���P�Q�������3Jv�,���(ԩ/�����j9�]@sƺ=�exe+��L�VVW�18Z-��+6@��Gd��n��f��[K�+��Kj�v�Y���YC+�$����`���2�eyr|@7DI�s����y�#�P���7���t��o�!U�U�j
T���K���^ز��')8xa ��|�����P�\1� kQ7�b�)2�d�s�r*��h�f����%��<}�k,����Y&,Ɔ���	�be�Q^����� ���2ڈT0�2�rkl%�0nX�ع�����:Ӌ	`�je��R�]#�Ɵy#��#���f��	+���e��w��O$JDe�kWH��3R�f�2T&ܿ�����X�E��S���5��2�U�L��M<L_�g�����Y(�R��;��"s�����v�\s�6Q�:�DIU�98I�'ì�!2M�� k.��X���lM��ŧ����wh�c���K�����2�c��2��ȕF5 F`���w�pN ���ƆW��y���`�~����o��Ӿ��n@�ƴ�1F�n��%i�Vk�a����3�$v�����l4��f�u���&f=7��]ZJ�,�l�]HSGc���l�P�`� IYK�XTC`+�[����v2�*Joadɞ"T\P�-VQ����;D��g�_����#F�Ს��+*AQì������z��Y`K�W(�?��l��9>+Hd��¦1�(r��/����S�jP��e���!�����&lj)��H#�G�R0J(3�(��Ŧ.c�/�m�`��0c���p?S:���L�hոA(Z �B������+���ڑp9�j]M��c�pL���^���Y����Y9C	RUq �1z��A>��)\\B;����_��#䆄��1%�p3wTc�fj�+q]��s�xIU6,�=ď�Ua(���̦��aI{%��EKQ�`q�u2Gq�?�)p���Gi��������3�S��b��`�F�Ⲣ�L�x�ՙ~p���\��pKL|IP�r��@K�Mҥn����$���?
��U�1�2����|d��i���8&��JVʔ�n0��y�!�2�ߙYvj�K�+e�*�9TO��0��Ҫg���3�D�ԙP���P�\���(I�m�\���]�ں�6����F�R�D��j�i�Q��(5)��a���(:-�HD�8��@�a��{�:�X"uP=�j��WX3����%�p���O�Z��X0��U]"�{���0n�,�,�\SP����,�.��R�o�|*���ă(�/1f6s(D���ڡ�U�PY�3���6�K�X�e�X�g_ڬS��3.n\�R��ibK�G2��8i�0Ws{��S��5H�eGL�#�G!���f����\�9?�,���e�Oɸ��>&2�6��{#(1�)+�f������Q���.*�HᛌsD6�!��#t�0��Aqc�SA%������b���.��> ;� 	a%ŏm��?ڑ,�K�ľ%FK�C���cԴ4B0{a��=l�{�1����*�F��H/B�
Cd�L�e�چc�#
�c�$����`��f�� \�MlE�քw0��yh�me��|:��q.吰�K#�1	q�u2���ԙ\��.fr�?b�1��t���a�L�a䖭���`�8�t��<_�j=Q�/�|CQ�Fb��vy�!��12�/�;_�&��H~��֠@�WS�!�b��П��             1` !Aq�pr��� 	? �5�DlP�� �{��vG���[��f1q�:+:������ ,        !1`2@"A03Qq� pP����� 	? � �X�~y99�SN*(�S''✍S���(q�����F�C����:���:X��Bp�*�*8�	�c�%C�<+���Z�Ouc'������u�@�\A�u�76��l��p;	^��{S�7}�?oמ��pB��\��wV��57��l�_'{+��kv���+H�I���ku�|��j;K�£���YCTq���O(fhP�Uu6�O�(�<Dc5j�T&�a@G����|Iɡ�2�:����Up�F��'�]� z_�+}l(U��V3�y���=8�i���~7��}����:q����PK   [��X��@��  ֈ  /   images/e8a1ea1d-d840-4bb4-a734-95947de726d9.png̺W\SO�5TD� �H��A� �7�E:��((Ho�BCoI�U��N�H3��	Ύ��]��s�[6��33�Y�Z3��kM%*rFrD���R��	]yq�:pGWwwx��l����,~D}n2x+y뺿���������9�9{�X{��{�g�I3�@�A*/���g�,xd��NG'���z�Q�H>��?�`NT��(H���`(�w>v���Eꝭ!���h���3O��(N��k�Wcclq/2� ,)Q�̪��t��'���M���k���x�_�Ҍ��9�#ūW �G͔���b񟼁D���w���W�/V׼���FM|��o������俿��˓_;����wcD�����i����F�x����mR�-C�T[�,G���Fn�7Ū����=1Wð��pm�~����Yj*�-���ҩw�X������{F8h.ӹ�}o���)�q>m�YG��G���5�J���W~�uP�|�_�_~Pf�)���?=M����"P�ی���C&�ѩ�ӽ�M}M׀f+~�ߞF�y>(�<^&V��==����fΈ\��Rd=8�h�2������W�/H��X��g�{;!��h��=��X�H\��QZC�Pӿ��o��i�:]�3	X�|��x��q�	h����#�.��nl��ںY��ۤ�Og)hF$��� �/TJ�v��Gf�����rq�vJ�R�y�I`���3�*�z=5�+Yͯ7�I��L�sD1z�Ё�������� ��k��Co�����M�����ޫņ���8Ϭ�����ps$�_w<&j��4[�J���f�j^�5��]\�`�:jȚ��j�7�}�t��2���JC�ܖuڏ�vEOO����O\�`le#D�5��s:iͩ*֮9+�q�37�d6A�U��cMG50��Ȣ��r+�9r�~?횓i��U�H�G'ŦW:J�~�ˌ3�2� Ο��}j���	~Y���?\͘��V,B-,��u��FI�k;��ޞ?/���hz��F̃�ŉ��!��w%5(�FI��� ����`8�  �j霡)/�Nsi3O
}�!��k�̉d�b�
a1��t7����*"(@��	3����	��6e��}�X���t)��V1cq�e;��I�	�A�<#����\����Ĵ�V5y/r�)�l�/7��+D����cPf�e�g��f�YO��]�5 ��ΠjO��U��7�y[ň�
h\�T&s�]���-��Z,�WR��$w�HA�O)����"���Јԍ�+��"��`��z����U�9;#f3�Ĉ#�&X7��|�%H)�77�#����<NA��\�7���O/��6Ź�L�2�CFBT���;�G�;����4�O����������;[B��N��ݵP.�wJ�r0�z�ݸq������|����3w��@���a�-(>�]������������2/��h�����_���]B��Z/2g����@����ۤ�-����A�	<n��}b
�2���i�؟3)��]3�>�>:�b��Ky���($~�-,�dv�%�ğf���l����GT���@�����;L��@���b��x�mp�[<5Ե�US���H�3�ִҮ#�ڗ�,3����w+�kT,Ѷ�x�Ia�h�=�l���7�Q-nTZr��_ߝ���)�i+Q+���E�v}$�g��\6��1����[d@���c�'�w�3���4��3�K��<Q��C�iD��&kel�;Wh&X���8x��Yi��k*K�����껅�5��\��!���ٔM���y"f�&俩���Q�5b�e3��b����X��/�~?l�	�~Q����{�+���5��'%��E�)�|����Fb$K��>"���}��~�3j��i8����속i?��"�k?���Z#dވ�)�]�`odևX�خO�����L�r��d��1���?��m��q� ��0]����W3�[�����7M��Q�����\�\�w;'4%Wƙ�h�O`=e���Z6/C��ݨ��H����g!���W��� ?���}|���ܼ��BpS�z�4ҸEmF�ٯ{V����7���I�4k,4T*����B;��z�B��Ɩ��D|9j�:�q�������������ҳ�D�&�/6��^��I��m�B�,K�͋igd`x{6-'sj?��u���5�*]�o�YH��,���6Z��Lz<�Ŧ�x���WJ2<nB�,i<���^+�WJK<n<�L)<mǳ2��An�,���q!��o�Б�u�Wk�Ğ�r
����>�01���w�x�?}�E^��A�+�V�m�臹b��LRP�I��<��+�'sؗ�љ/z�0N}�&�4�P�e�(��x΅���Er�Y&Hڡ�6w#��n���a�����zv�K'��˕v����̩�����sE'ה�?>
�9��&�!�O��vL�-#�M�R��+�������zm�\qBH���)o��v]jv-Q�!+V{TΖ�J�z9A.�����E���Edܨ�-\��*��q�M�O�W�F�0���C�Q]̚-���B$��������L`�!.}Y�4M>5�
Zb�Ub������V�>�s.�)Lx	W@��h����Vϰ�&P��z�������Rʷ���U��q�Z��kf��k���F��{�T55W��OL��9m�������H5�η�-]J�.�t�D�@���ݪ�9q�c1G��X�n��t�BO�79 �a0DW�e��+V�#���s|���c[5q/�@n=�ŇؽP���p�P���E�b$�%�1Č�lo�QHN/h'��8t���D<��a�]�dP)H���넆�}���������h��, ��0jaη؜�����ԡ#�҇-R��c����ojFBs�9����R�ֶ��NڤubA�rw~�Py��l�N�	��v�a�{>9���X\՗A�[�@�����}#U\_�+�4�,����7[�"#�Rv
Ȧ����⋭q�.��p�ϑ�Jz��c�Ve?������R&ΰ���I��\��cc�?]�ș+CW�`系W�����������Kf�_i��S�I�K!*\��"y��U�篂(:I��d~�V|��?�>s���'�V�g��<��w�ش��CH����߂I���`���-�Xe���,�'U�F��8�鶵��*`1�d�z�����rg,ǁ��\���d6N��A���Y��<��WA;��-��4�������C��rLӌ~k,0]���{��U BÚ����z��m]#䐐�I1K�$�����k��m�
}�sgɳ��ug�Sn�R�/e�?EQ_=W�.�+NC��_�)���q�lf�F]���Ms���(d�2|B�q�A[��6��(X�����'~RL�Z%��D�h|pg�� Ձ�>�z�x�+��n^BB��0Zᐂ�)�����؜CΫ���X�rK�dA_�R�aa�c~nT#c��dD��P��w5��m�!�T�!;��	iN��
W���陘���4M�W�N�sq�{���f	̊�d� U����Y�_�������~ST3V�]�?�ŔE	i`d�]���և���'ǜ�:�f���;�nqԬ�f�O�r�V��L��A8>*:�0fV9�v�B��8�P�w��wXc�4��N�ڵ��>���ֳ�n��_�������ɨ���i���� ��.:��꒖g�$����(h��~&隕���w�am���^�j�9I(�8�>N��L[�6W����΅2|(����ܦ��Wo��K��LH
6��q�I\�x�X�DM҉�<�'�mk�wmC��-U{�|�.�:���z�E��L����~߿μ+��u�����]�7��xQ���DF�r	�4ҞV�j��!.�P�8������Ӡ/�?���w�PҮ ��ݳ\zC�}C�ܵnË�iMY'�8F5=��OU��� ~�v�FN�3pl�<�����,6%��!�X?���+�D��P�VC֚[�w!�<�L���hTg*v�X�k>��m�2�:ɏ��a��K���ƮT�{C��h�:1QY�=3m�i�o��e�m���'�v�Bb>� )Ҧ��`%�z�N��3���hXO챟1�f���R\��Ԇ���,�g��3��W���j)Z�В��ԑ2hʆEYc�et��VE�j�!k���oIsO�lU��W�j��~��^�t�D}����@GĬ�����������,�}j>�4�w
��>jvNyY8ug20��ڳ*'�=�VC�ưۍL*�Z�F@�<~��3���N)�pRص��G��m1�
�a�M'ud����[{�M���"c�V6MB�ɓ�l�P�L?����?�Gϰ�<!����e$K�	\D"c�h�8?�q~:H�qq��0��I��Tʊ���|�@�+ 獸����@�`u]���:o��"��ݚI��;l����V��	5R0�}�i�}�(M�4��wΖgN��l�An��Jq�6�7�V�^N���j�&�����\�A|p�~i-~RV�Z�m��uMriiQ�u�Xd�d�����ː�$��A�$�����ee��V�W̌;�A{Y1�D�8~y�{�N����c��1����M02S��6LquW�6vbΪ�5e��`7[ �إ��?�*�t�$�j�D������'�Ӆ%Gxc5tz���kN������Ͷ:�xxX�9�Ji�O����c�d��g�UM�ٰ{�ro!,0��n��iB/y$Bj��v�hx�v�wz�(��?ג\^������qf��u��j��l�׎ ���"A�l`��aߐ�󥯠��w7`��%-�V0/�����o롦%-��΄$���#�B ��Ŷ����r������q�S�T;yJ��ͯ������>,��*M�op�T�צ%��CM�&׌+Hw��n2�.��9��~��$�I�Z�ʋi(��Ғ-.[�mj���6n���T��Kb�V���m!���}T��CM%؇�9�||[�������Im�2C��r�H'?�9Ƨ�'՚z���۸%a�rK,�4�_`&���d��~ߏ8^�
�_�"D��������3L|+Na�SL�K
ł��b�U��|�l��A�'G�Jq/j"�0�L��i�	��B-Jo0�Z)�x��έ��S���������Vם�,���ON�>����h��X�.��4&�Lg�a�f	T�0������I��Y�E�t�v��8��v$!����-�ᅲФ���0zyj^eZ�M�"��ss�&�����l�M�٨����y�ޠ�,N�Qi�[�����l�k����e�Ί]�>�]h��J]l���c���ЩZC�����9c��=2aj��}:�4�:�>�z�abی1�"Q
,��<�hbY�E���hq�yI���g�Fr��Q��D�'�Y����IХ��L�k#�~�f��q��#�"g��lAH����c���p��yչ)��Yer��6ηA����Kd�Z��փ�{�[Op�"C�NĐ=�*�>q�����R��DI���頿�M5N�.4_���J��0x_TCx��'b9�P�br^I��s�$Dx�U0���q�}�f�|�P'#4t����v���/g��n�s5 1O�Enz��V���#)���)Ά)r�����`p�}�uҠh��T�����4���+	<����&��!<�t�o<�ĵh��;_V��h+�` ���ΌR�M݉�Z��"��V>�l/,%TW$��:sb����_,�q���֍�?��h�s���H6�;�Z���J/b�3��2Hs`��]��c^~����rI%*��]c�b|`%�
��x`ó��AG�"m�~�KÛ��ŜJ"B2|��U߉V�J��N�9�ݦjxV.�-w�Loڪ��t�]�dֽ�=	h ��+��$��Ճo�"����=,��%��h�s��&j�&��0�%�:T��,]k���R][���}3oW�2��I��&�T�"ؘ1zFd;�yQ �ג�E|�0.�p�ԄN��4�W���*[�a��$ ��9����*�Qݱ=%W�Xz*Ef|8�uIq2�zDU}�����3����p9Z����or��p���=�˯;`�a����<��Ţ*H6�)�Q7S~|[�#)��C�O/�+�g�p.f	�k*[Z�|c.?�&M=m�:
��G���@V��f|)iie߿++**r��"[��f�}�[���m��߆��^aY�J��V������/ �sc_��Q5c��ޮ������k�ױ����A.#��e���0���?�;ay�5m���V0%%eINTF���M{|���-�R"	�C2U�� 9q��_�Z�HV���v�Ԥ�7݁��Ӈ�\�	�Q-ᦨ ���Et56z�F����OM��742�!H��~�:���0�ʛ���gh����X�/�V:K�]vD�w?|�0iY���1�ws�B�L���c	�1v��b�%!�'��T9gN�!tֺeH�HL���uSr�[�L��	؃���݈<�=N�J ���"Evvvch^u�k)����
���ɂL1����ؠӭ�QWRGC��or랄Ӓl+�p��x
݊�\�m�ٵ_/�toz7R<�Hx!o�Ԃ���-,�7���ᩓ� �=(�d�|ǟ�oaQKM{�n! Snk�3�,.fu�����ew�(Z�����Q�)�pX��Fc���t
����T��kنC�R�#�����wد�;3�-Ԥ�3J��8F���'��)!�.����9�y���Z�d�X�<ǒd��黽�7JFZF�'�~]�}��?x���;�@O��O��bYJ�P��m�����������Q��š��������jj�::Ӝ���++5EDD0[[��x���&���R2j3-Ɇ#ߘds��v����?�}�.7��Sm(�������I�C,V�d��릕�K*�t�;Q����ip��9���ϕF*P5D���u������S��@&�W��ny��UFVV�1���3}�⮮h��6vp�s@X����3d����������$#����&�dpppjn�a=�/�;/"�����&f�����xxL
�ֿv�Kρe���SOP�7��<Q�Ȍ_�k�*���P�Ʃ*
{X|��I�vS�d�!i�ycde�n	>��wt�zd)��Y�)�ZU�����䊗�BxTt�nS�S�ɹ�oׯ_�B"ˌ���=���X;���f bpt�ңrhc��Է��:B��hN��+��L��FD߭���������^��RȾFi�@ޠ��6 ���i\i��,�}���""���<��{&y@&�B{u�2b���}�f��\�$Xt&�#/u��0��Y���Jy;�M��5==��
>yt¿��?s�~������mS�K¨�+_r��ή����֤���^R��\ԫ`§�3��uu�pQ��NR�k��Yd��������U"b���c�?Z`nl����m$��ȇΩ��cR�^�W�>zu ش`��a	��{�;sy����!歁�II��U9ii%}l�f��馊g˃@� #7�-5Ӿ�l��b���n)}u5� }��=�̀@F��ΆA\L�ϳ /ٖXgj�B4��w�H�A�5��zw�����S��֖c�ߕH"LkcR�[PB�		�>u[�sU͖�����;��W�"��~7��ݖ[���H�{a����Ey��xS���1�F�Z195�n���~+�	��[T�Q3��J��cSx�ޭ�>�7svr�ɖJ[b܅TV���n����s����w��j��;�g�1�!2�ul :{�[;gX�-�����)g9%�n<�y��*qR$�xg�#�����"�aճX�j��N2��=�651Q������+� >�m�_9�]��jDD���ܳ��:��[$������%&�GU}���	<5Z<<�$���b� �_׿~���K�nF0�*��#0�2�)�舣�=�lIU�H���ӡ������Jss����S�)��6L���?X뛞�o���X�iB���WjO=����|?O��t���S�����\y`\fc���@����/?�{�𹩩�{�7���6���=##� (�[���������h\��[t�
�b�8i���(腁Jk������s����E^r%��B��O�7
�gn���������LDm��QO&ho\;^O��c�����[-�Y�����YFՌ����D5UU�kǍ�ShV����\`���"Z�%�i|��o� �@���fD�)��\�Y$�Bm�/̵ָ����PYb�Rwɹ��]�j��޴���9oprrJe�A��cW�]���g8'2QF������4 ��2����x�3j�`���3��E���� 4�.�9fd��k[[�Dm߼.Hi�<��Fa:�.�u���h]7�''v?+zP��"��7���JfX��%����;�lnV���|��o��ӱ�l�EH3S�LEt�	�\V���n%�Kz��3�O�FJ����^Td�y0>�PoQ}G���]zZZGo�㋚�8S)�Z���Q3����R=cc��ꛀV�8������T'Ұ�1��W�R�#�R�!��VM���4]����$��S{�G�kS�W��ͤ��N���:%�"�
�������a�t߼�����,n�9�N^�g�ԛ_�H@s3pW$]vI�ޢ�7�'��Y�nv�O��/��k=����.�ږ����ڨA3��)��ת=�s�v܆�V��0�
�=d6/�����395���-�� a��p�� ��9t����|q�Ν��
�8������|��Q���r-�_�uw��Ǧu�w�kؙ\��̨V�Fn%{E�4O��&���p6����9��M��J!�`�;��L�Դy���X��n�ͽ_�W�4�p/2<[�3-
yv����|7H�"p�������Y'#�|Sçk�9Ms����>���[ZT��{��� ������x�(�qi�k�/Oҳ��J]�Ѭ�:NP���|�c�d�oW͐v�"c���WT��}:��������6S#_%y2�����Lz�̌�	 ��s23'���^����~��Ξ�r����9@�ۦO���ő������U�V���|p;�je}�H�>C'�Q�N$��m1Wk�p	�򬾈�t	�̕;Z)�����ǓDT�ػ��bOb+Z����/7Y�|��TZU��P\hm�ņ�M:;��$��2����ͺ����ֹ��'nS�`Pz�Y�s�o�l�^.���J��d0��Ч���ٻ�3w���ڦ��PWw�����V,�6o�xN�o�Ҷ������>��77�jco�U|kuV��c����K�~5Ӑ���i[p���m�xZ,�5��D���?�{��vo#�z�5�=��rOLL���A�.�;:�~���+���M�$�QCs��������#�ۏ<����l��jlm9ﺕ�Zxс���zC�N�)��֙$v H�	��5O_������v�R�9��T搖��q�Ѡ)����&@a�$�G|X�Ŧ&,(�ld��S�����e6hr��MM�C"���gs�� T�����!��Q�@�'�����p�}0�y
���)�T��n�B����� ���pM f�H+NN�BBB�P���v�'����V�����G�("���h!kr�8�]���\hFэ$���������=t��S��>a�з�ml��0Sػ=[�/w�,NF2���K_$�t麅�݁OZ�(��{�"���sNx����SS�@���|��n%޿D
|������q�� �.�^��WA��|ek�*���-w��h�oqE�a|���Dwgg� ,�VPb�SA[[{�h����n�+]I��96b�̞�ܣ�e�M"g�F�3))�g��Q,����[G�o�W�w��%����m]7g����/����S�PH=�
�k�r�L����̅�e�	��IP�����!�	<ʾ�#Yxm�yG�� �p�=D�1t��HM��>ۑJ�YSo�o����I+{� ��f��̻����Yʪ��P�[{Ҹ���3�����nN������ଦ"�_��S�
�a$`��)[� ��d��h�A@&L��K����H��0���� 6Sa�h`ut��Gf1\VH���Ѝ�(��I��N26@n�/��P6T	�h �-�k�L4�n��y1ӌO<h�����P��w�yuuu�V_\\L��& �k��6�����#��4��~ ]�ЙK�*��A��o9�~����Ф�M;Rj����͜��T!�+�[���g��� g���&1o,f�����^D�̌�������J����o��-T��2���>FF���S����RDp?�5"��C���;�d��:Scqo���
d���KT�X�@!���L	���w�/�Pg�^[t�7ng>���Ą΅qЊ�2F�o�wI@a�5�4u�f�ַ~��������	�Ɖ����f�0���X��^J*M���]���^��~���a}z
��)�K�o��?�x�yب~*S������n,C�qa����B]��&6F*EX�|#� �K�LYB^�%jB���}�����3@�24�-.f�M�������:�/��R����`�3B`�%6|��V���}���`@X6�/]?^��3>r���V��o {����:~w���]e��W�5Ǟd�����S���R\�7���{34��͙<�U���Z3n�Gگ�Y��YC����3��	њO,�����[	|���
�ݻO����O����w�*"2���Y�4+�@�H�I�� ��JCU�t�cgM?��64'���d$��t�*;��q[�.��H4���,1��&�Ў�k�Ɖ���p�Z�`d#�K�V��m�X|@5*��2Y��("����y���3�7l�2wW�1������405�Ϭeq���Oލ��5�V�`d����	��nV�Ջ��F��\��ųn�u����uo�}6�ǷWK��r�� ��)
���rX����u[�T�74,Y4�f���1W��e���`�����g��)�6�����fԕ�,n1�_�?��y��\o?��S#"��^���{��B^���N��xI �fe���s۾~�h1'[�]����Pw����Г#�-�(a3?�aD<��X=hP�̚���Ȣ��颍-:W<�~(�/���|V|	�Y X�"�e��9������F��^?�th�Y����f��߾��x���ԡƃ@���[an���a/��e����wl	��c���ɒ�j�.gr|"~g�Nr�y��I�^A�"���(�OR��=�["h=�_Z�}��\eX
�2�� �H��V�,v� n��(D� >كy��
6n� ���+���6�2F,'GG���hkp>�yv�훶Z�o�{��^F��x|z�r��R��1��W�����+�Y	*|~bő��g�?u��zO��.��I�T�&{�@2x�MZ�%�T����j���~GP���j�>>>\�ԣR��O.�SMv�AѨ�����B�pJ{2���C	���v�1��|���Vnyxv�����	V-Ҿ�`Ƃ�.̠���25;z�{h���zu�®�� ĥ�o�Q3�vt��LDD�(=��Ӌ=k��o��Y;8k=8�8
l5���;<:J3W�c��47C�[ZVU�"L�F�5��C�; �K�U|xkHᜤ�4'D��8����+M��69�
��{�c��vp���s��b�^�]X9L��2��D�L�ō��B�;��]�)�a��x���:@�i�<x�̘��)$]brNNN���F�'
�� }�V�γ!��w
 �P���5����۠0Z�n�a�B����-��CC�]�ݧ2�*��8M'wꩌ�>L�]��4�V_ŕ�=/$?�U��9�}��w���Q�/�%`wJ4�M���%;$�[�0"N�G�;�<:"Q
 #W2�.�����7^��jm���2�zگ�L���bN�X�>���ëCv�]���$b��pI�Ü�W}=~e�q.ퟌn[#�=�ˉ��,���/y��-��?
=kG�{y u���d�EW�`�0I����d�v(N58[��]�M�on�3�*��D��3��zk@��|�o$I�N�~ky�s�v~�i�!�S���F=N���Z��	���Sup�N��N���q"]Ȟ�<kyb"��Q�(�~ww�.������^*�,,� �rʬkiM�|f1z���R�v���E�>�w�߄��V��քߴ"6:��K0�{ZZ���x��'ѹ!F���&���v*ï������?�,k�Ov�w�n���a����=�ezPϒ��t��2��f�lS��Ohkk��׷pj+^�u����s��g˗H�`�B��d�P���ڻ{�+����	=��*�l��x���xأI�{�B/ٌ��^������%�w��}��rثg�Y���ۛ���^*�����"����F�,bf�@V�|~�$ku8Egd���R�S��\�[i>���-���F�U�?��)B"� ���g�-^+���������訨u�2K q_`�H��3��z��|�{H���c�%����å�%������ξP�8��~���a�C^�s��E��.�j� �7l��Z��"i�*�s.�C>7��h�m������5�)���ه����p�В�$��� \�39�>�m������t�Y?���b�!ٕCp�j�ʧ߿�%$*���pTQ�؞��P�����ga�G�b�
)))��=q���σCC���@�(�c�h���-,*c�T�SZ�	�����)�e��Y⻿L�؍6��k�}�Y�W ���>,�񨚼�&�qnշYW=�[��g�)��4ۿ֚���j�����}��e��Y�i5��`�[�M����g�WG���>�ճ�]���
椄�'�����
�_��~Vh).^�:}���#��֯�������oa�L����Ɩ�ؼ��u�
�?�g��l�<::��lLOM���;�qjf�nedbB�A���b�,U�
�/|���ʑ��f#>3�xJ�m󽠜]�#�QB�%�
��J-����z���Й�f:Aʻ l��NhZ-ط/��Ϝ.��{(q�z0����S�[h�U�H�5W�ǎ+��T��h����%>;�G��?��/�&+K�����~n���(\�m�� M�^�%&����7/ ݎ���wu�-5�:88��e�=T{~D<��b���9�j�ʵ�8��� ��ڣ�%05�gŖ�m�{�v��gg�LI�1]����������G������싴��<��Ћ������'��?^��m�R=L�))���w?�Gv5��&/D%�	�?��;��둞��2~i���J� td�^��N �/�:'��X�uתu{oB<q�BU�G!)��e���d`0`��x暐pp���q�@iu](�`0�pMӯ��>�)�4�M��������p� ̚}~�u4��
��od`K��1�L��۝�������ǈ���+aw�R��z��΁�վ>[>�����{�z̖!}���9��ᴍR{G6N���E�e�A�\N�-D�p�Ѓ�z���M��[�r���:F66�w�6�� � �h���WHN�d�!���d�0�F;{/
j���_�
�������Ҭ��u�,�`ȴ����;RQ�1�&����N�����v�O��E:��5Pޯ)3��!@"2�������LNYM��)���ޯٴ��j���S)����X k+�7�[��9(I�8��H�6���QA}p�R��eG
�Z�i�%�G�81��:���c��[�n�P8��pi_J8#��h�>J��Y�k
w�dy������e���p`"'�׊����!�du`H[�%l��.�qq�G���Ӯ�:��e~��Šs�D�7ٖd�fB��ˌ�.���}��;��-w$A�̌�lsm̶_�$��{�r�]���@(~���?�gX��.!�7�\�)�>�Z6n���;�?�v�*�E�������#���_��x��U�ܒ~�3vxx�g`PE�o`���ɾ	,�X��$|r+�k�-�.��`�'�i�yW�˭�%M]-a�r1+�u�K��S�cD�.g���5C��Sح?�t٦�b���g˽&gp��]|P�y��������K����N6�^F��ܹF]�0숰�RK����NC�OJ���Ԃ���V͖ML����Z�:p�Hc���"�h�բ
H*��R
����G��vڿYSC�Yˢ(HYk���>���� I��B��j�ڑ�{%�ɫ5_	��C��%��k!�q�̤N�If2�)�G���s��Y�Z�+�q��F�:nZK��z��+�4ǝ���a"��U���ů���xX�<�������]f���P�	�
ُ,�0]�oG��Z�&
��7l.b���n��
?���UC��7^B�	R���?q�]���m�(��Z�@��<���짽�F�f�,hu��C�ķ�E���Vt���?��g��.#�`������J]Ϗ�����jèm�&�M�� �w�3_`���j)I)**����l��W�tu����0?��z8 1;��E4t����m� q&�.@��\X���9:���;dD�J�5�c#�VdT�bƒ���[��F���ݩ+U=�Q�Y�D���{,II�g`�~܂A-T���|���]�y�Ƶ��3��P[�:�CVB�@��<,��+J ��E�U���M�d�g8JzL`�њ�e����K����E�f[�sBa�+Y.���=X��hU]0�|���i�>�S?�i���U��:5�B�y��Ex��0U��C����Oxt��CTD��n��͟t�k�s������}I����Q��<^S���
ޢȟM�X'�O��"�M�Jra���{�l���Z�J^�v��$���*��V�y��鎞�>WNv���~Q4R	��q����|��2tTc����3O�{b~�T0T�6�6�b��d�*:��d��@��`|3��N�����h���xlj�[R��][E�Y'�A�~U�c'1���֤�ƫ�r�{��SO�#ˣ���>ǘ���ͱ�Q��u4����L�vQd;�=���:;&��������3��Ĳ�Х�4�����4���@&o~�PW�8�u��!�D�BKZ��n���N�23�5{�$�u��D�$zڋSV[���k)���	��#��B :�/Y���֐��6�WJJ>��1qq��MM�����n~N4���ˡ�����E� ��q�'w�	3�8xL@	���ܟ=��e(P���#5t�aK�����?J��γ�$���*Ô�G��t&g�	8Ε�;_�B��jl[�a�����Ҭ�P�������dzZZ������,��(D�n��Ĥ��1�1-&(�O�^�X�hj��@ܼ�N�w�;@[eA���o�)�(Ұ�%I	-�0�W���%0)�0	j}Ǐ��u����������w��=�L�C���:9��ܣ�&WWףX,Ƿ�?*<),".�����v����(@	�ȭy��m����ծ�@���
�	*�Oe:|7?Mh3�����-���D�k�e���0��� 	}L� �҆0�1��-UW~+PYAI��3�� r�Ц&� 7_�g6 �ه_���l �HlSss���?YDMKOo�D�H�d���f�ʯ{� ����f$R$J���>�=��mA��f��,��]0L�閞�B���x�O�wSS�G�w�L{\�H0S����&�����-	��C4���	����w�{�,�������3���w �E~��O�i+..~� �<�R�6��Ի��g!#I)�U=�§�8��d��(~���M�l���(���΁��٦t)��d���<��J++g �Й�.	kd��{�컫���08���#+�LGG��6��2���a0}�18���Ζ�ُr�ա���m�c'�Κ�Қ�E�j�I��6��j}��ݏ���:���!W�v�_!r+�b�d�VYm�aBw{�@���_W�;l�T���|v�(���.��{ tW�/%Ԏ�"r[[�u$�ȼk���-SJ�Kw��$f(�ٽL�� �֠�|���7ܮ�羊i��ѻ�=wfCV�8D�PN
�q���ŷ��~��^\\ж�4�lo���&122ޥ�ξD��
�,��S�0a�u��# =YZV�V�G<2�=���٩ר
�uxQ�ydU�D�+,~w����!�/F���z���0�UøQJuu'<9�/Bq{R��gmG����j���/Ku{|�+����e������\
�eq6��q̻�~����2TC;Tkk<����������+W?Ͽ�_<;�H�չ����*��>2.!��~��-�'�p�\\:fI���><m!��'qj@�<Z�p�&>�EJA'.{���-Y�[�	ml��d���&� �4rh��������)�m�WtVa#����P	�;�KO�·5�����
�)W�ɩ��#a��s�P�kY]�nEEfs3ޮ�)��yV	I�}�~8;g٦&��/_.�0�J�Ql��	'�+�0t����$����c�śE���:����
;|ph��6�[��FJII������A�ǎ"�(33�$���5�MVB�I�=�5�w���H.��H�ݣs#|��6W���T�$�k(p%�Q(^#�}B���p+��]!xo�{��1$<E���e��R������ �2�uo�}�7��w�"m�9O6�X����kp���M��#�14��ea�S;>f����p�?�ݳ>3{{siB=.�F����i�ꚸQ��"ȣ�HW��{U���{HGP�(R�!�B%@@�މ�Ф%@B�Kx����Ϸn��]������3�g�7{f��W�m�N�G�^�>��0�2C����,		�A������~t�^�
�I%'��a�E���e�>ڿ��� Ej�������̀f��y��d��-�<;����Xe��R��z�M�LyE���YAB`����'$$�#�חu�o6y�V�txL��뛲^�߲��W$�<������կ ��h�-?��x��4_x� ��*��wN�d{��Իǀ[fyhV��eu{��8L����l����z�Y�����I����l�g��cSOU��*Ʋ0�-G�Yd"�ϒnm�Y�j� R���Ҷ��3�b�s �Zƍ�-Ve
�?£M���۷I~rE���j(�#w�3�2cA L������#C	?��t���w�ja���snj2�K�K���F��ӛ-Ɖ�%z�>�뜊^�|$'����$�hy�hc�p����+��C��oFQ���t�)��u�}�ǉm��OY��}O���"�* ��z�eI��|����ȳȚs��A�-�?�e��G��X9:�ʨh�!��Z�V�tbς�F�#��
�}�ft�׽�l��㢝�R���D���g����V����b/Ox �i@Z,R���
�8�^$��e0��VG��۫�Τ�5�ȡq�?Ϸ���� �&����5��u��E��	�'R3���'C�b9v��ēn�+Ǭ8͈/K��,��Sr�و�A�Y��6ķ�Ɔ���e�OJ�
_�J�S��S(���[Vx�꽞�G�!�p�;�v����Qtmm��Oٕt�+������!X ��þ�k)���/��5�?I�&�7�U���	0�3W��w�>��^��d0>�'�t=�3����m�����R�n���=n	�Z�׮�_	�7cq��H�4�5^��A��V�7w%�->���E	<|Ϟ@���|�|	����sm���[����{��&p�]x�sk�L���Ɨ�#�s,�I#k�D��m�����ֳ�_���l"E��討���u.*��? Z���I!����U�0��2Y�y��`�>@�3Ic�*��AO'J�d���}J\+��BE �Ҿ��E)��j8t��;��ƈ;6Wq�,�<>��J��|f|[1�����'ol3��׵�g���D���[��CD<�ޟEſ=a�UDY���Ŀ��݁h����ٸ���vZ�ś&}m�=����e�0W�6r��R�����[�|��B6�9����ƛ��K�[��G�5��_����)e9�g10�D��[�D�P����Z���j�Ъ�j�5���+�)��\|:�P0�}��lH�� U��bk��%&��'��)qޣ:�G����Y�HO�'��O퍌�I6`�S���i����'�ݬe��������`2P?��A�<�>1���%��Lw�r���qD�\�a��bA�y�y�'�������o�r��I��qjU � ī>��#�(Eo1��d�C���*_|��6;�z�<���`�ˮg��U(M��{Ǻ@I���S�}����Բ"놨���݉	C�{7x��i�O�AC�3����|1	�H5'�y��Lf����>�ax�ue��D���p�h���)��o�߰��5�ZZ��9)����(b���4�� ��_�j��'C/y���{j4��o[���+F��G��U�A�&�h�ݠ~k�g9͝��~!/kr�o��#�It��\㟺���D��Ԣ��"���d�R�(�w�&�0��C7vǙ� T���'��]0\�}b����Z4MA�G�k@���[��(��ыQ���*L��$�$c�f�9�d�}jt�ć#T[w�ؕ�rDc�K�e,Bx��f�A�P���mJ��G!�����-~�l�\���'�}[#������[�!Iov�@ēl���Uq�g���^$!h3o��7'Nh��;�1e��	�jC�6����n�h;��T�0�%�h7�/ ������/"a���♏[�T��
|W^��Y�j0I�]�T�9�0���(<'Rc&���5�<?t�Ab/̆<Pô�֯K0e_��V�������k����A���q��>nƤc�\����T�:֕#%�Ԙm�s�����G���]2I��� �R�t)�Q0���bk@�0��;s<��/�E� I�,�*��'%۫]�'�hhn)(ĕ��w��^��������L'�#g��fF����^������ظ���o,do1�����(h���M��3�s��oB��M���zƽ�w�T]���K��ܫ�SwF
���E
�ŊQ�FR�K�6K�Mzr+_8R�{[�$X>��%�]�c���<6
��۠��|�l�HbL��d��Jۖ	.b�IH^l��kj��q�G4��3%���)���"kV�,�gIr�.����>XF�愹�({���c�Х�W�[]�5�C��Z����I���_~_XWx�R���:W��2p)��������x����^�k��Z�1*\����I5d(g}������:N~�<�/4��Q�3�+'�P'��	(�/�.����G;=g;3�FԎE�i���a!qUaR���
Y3|�͜X��^�>I���8jq��BCᆔ�ZX��	��(k�k�a�g�<���fW��%ÏTR�77?�+v�	4O���GЃAY�y�����w�Z����O����[��#��Fj�sB�w'����]dTh,��4�x���������#�	9hn��7�?�����	� ���"ړ>#W�l�}15��ͯ����6�mQ]����&�:Ȉf�N�Io� P�[��Fa�ѡ�;�.�)u�@��U���=��6хt� X�Y}��Ȥ�HE]D�Q��"�¤'o�#h�&���V~�������[Wƥ��t�8&�&��U-���u52{V�Y0�7L�Wt~%���^C~#�?��Ʉ��DIp���W4zm��=���4��:�	�(�E�~R�ৣ��B��p4��i{8�%�*R3欳�=���>�Fl|�t�*Y,U���Q���4�)�>嵏�D������	KD��f�r� �]��_�Y��SsRS�1j����8<Ύ���z�7Kה<��:�����'\{�w�j�X]����பb�$����z�3L�@	����6w<��o"`u�TyM��1q�!g>?�f�[�;��������X�Q��m@6ih\.D��E���� �_j�`���3�x�����x-���^�;���������)�������O'y�Nt�Bܱ)vk�8X[�Deo�����{QxW$��Q6S���t\���`���+~ת��ᄬ&�����p�^�I��Ǚ�k��o\Db�8
.T1C�܂�t�N���rF��($^�a˵'i��b��=2�cc(R���;�Ɩ��>�?U��z�G�&�+OJ�ZT�M��Ϥ�Ѫ�G���W�oU���G�N(�{�vHy�b
 ��ڜ����Ь{M�;�W��'bV�[����U�Hb�$Fd��h����6�Y����;��ibF��E�p��B��Kv��)ׁ<���$���B��ŧQ..C����O���w���z�V��d�+J]	�Ǘ�b��(�\಻��4Wq��WUHGǸK!���g~zLژ��K��ݘ��`f~bD�jĶo}�x�S�~��}���z���#�'�����hF���믭Ѝ"�E<�#� /���<x�4�A?�u��m�6*eQ�k)��쓌�6n�f��"W�Cé�Z�`��sI���jHd�DFB%w�����'���5�ޏ�h�r�W���hjϱ�N*@�&k4G�L\��aL-��||��BE4.�,�#�$�;�����a*��X�kT K��2O3y,Vc��z�`�L�`l�[��8?H^�
�ܩ<�h(���"{B&H5S�ϡ��ڳ>��=o4[N/��s���L�3�� �D_^�]='�\
q҃�О8�kuN��Vx�eL�jE��&n�D�;�����ٶ�=X4z1��>��m���G��=��뗑�=�,Qa������������:���<&F��%B�Z/Z�(����/�\0��ss_�=î`�z�����fIJ��+�&�'��e�X�i.*�'ܐ���+�8�>�}"Lv���ޕQ������M��������?�ݩ`k��]_r��*~�����HIB���==�v�\�U�Ӛ�/���C/�+�������م!���yN��Q��3�ȿ��a����/o�ȺnI��A�]<�
�b���,�oT{��f�o������d����4�w�?
�5��H&��"(A?��=�`
������|{�jc�=��-5����s�7%)I*���Υ�d���ڻ�N�ͨ-�'� J�(M��W)��E���|�!|�#�k�%�_�=֐v��mn����S�׹x���(����w˜�i �rS�L���Ј|�N��Mq
�[��~�.�@V�j�#�Z�Uzm���)����o���������I�s3������W�����M�&�2<2�Y[���{�-^G��E�*%W������A/|�Q�|/B���F���,M�C��DH��Wn����'O�l0�-����cm����� "�%��}����h����ml���t�9��:C���a�f;�|K�������峳r��O�L�|�ud�i�&]�'V���c���Q��ƾ�ic��ʼw̛o �&L��)�Xt�,����4�B���ӶY��k����%/ VѤ�M��h�Izv�-�1�9���D`��)��)�L��I,J�4 ���η��X-i �>��T���昌4�N�`��� N��#-e�Ŭ�}�p?�Ap�f��W}��A�O�"�Y9K�>��5��>=�����c/�Q}?;�~k�z�9�nf7(�,�8�tv�C�P��`�5%1�RD�?uؗ�O��g��G��z�r�D���5T�)��6�#�b]�V	�m�4�fgk��?�~@lF�c&�i)U�A�#u �js74'V�����-���j}Z�$8��Rkd868�jI��a�zh��&�_*'l�B	�����a��c��l��8��Hu�|ս�S��?Gި�v��fJ��x�=��\�a٠UMy��0����8J�m�4�u�����az���dKhHž5!�d���V�e����t�����H�Ђ�Rw�wc�`a��A��(\oc���"���{���Y��X����F��n�2��!M��Y��K�Ǎ�N�5�0O2"��
ߖ)�������׊a���X@�pviBy+|a��%�o	�|����g�R%�mn�����)�x�U�V�'���A'0�|#V�;hN�-t��	&
5����-7xM� ���\�`�`0�A��%���u�sP^JBW�*��w����&�`0.���vz�$%Mz�o~�}З.�'wc����y%ó�4(�
����6h�9C�>�Q�0�����d�s�����y��!K�
�c�D��y�a!����kZ����O*Xᘟ'!�P��]����vPsнqeO����_B�Du�)���a~&iÑ�o�p궕���=�r���K�5,,p�g.l���w�[|��Ò���HF<!�т��?6ϰ��T��i��~�w,������Ɯ;�_�a�'��B(�ƺ䐦볖��m�\n8��o#eu�I�@�ι��ҵ�T ��v_(%���)�:��ٚu��G#8���y�}�D%��ƚ���ޚ���5=cY��&�of���'Ak�g\�u|xk��KM�ŋ�7�ۯ�C�������x�Q&�lA����n)�UQʷ�F�ˬ=2m��Y���e��1�E��S����u*�f��n�=�a�cK�V�N"6F���g#&�Y.��/�K�=�m�۾|F���Y,I�6�Gy����,�1��,bZ��A�d�dOV�m�RawΊe��_s�t�gL��V��>�A\_G��^abd��נ3��mG��ޯ�73�웥�(}�Jڝ�t8��.���!#���nG��W��esf��߻r@��*���E����s�j�����h����^�[L����P��,7g�D�4%=�w�{�����&b�{"X+ ���(K!GCP<���eRۅlM�"ϒ��l,�>��T�[,��?^H�r����\�/�����E)�o�z���x�ν�*��:@�湦�˽~��׿ 
2E�36�n�,0ȂӞ�sc���B&[�gI��SN����P`�GVc��]��S��i���>��Vbh�����z� ���@��M/�6��y'�8޾{/��fk�A͍��g&�V����=�n�Ȏ�q������7~�����ҹq��N������G�
�a�f&�Ĺ)�d�da??l�u-.u���� �����3-2��F�}�Cm� A��.��P\��3�Z/s�8?m��o�ZHgwq��l_<���-������/���SA6�;����+��sl댏��4|�=5`�5�|b�����*S�_��KH�"\%�bX>��F7z�0Uf��?aCl�mIeN�d�����!����3�e����O��ۧ��+���VΕ�ۄ/���8D��6� xK��i�T���H��,53ʈD�<�n�&���Y{��)�|��s%H��!�rdyEr����`�ξ��h�~J�H7N�7�x�K�Drd�aR<2	��a�����u����bw=?`�V�e���k�-}����JӋ��f�����[�9���L�<�΁�������+��v�U�b@��� ���`�ca���=�2/�0!U9��hn�q��+8�0��Z�Ø��k�d(���p��V��M���u-�͵��2~�g�>q�l����_g���y�Дұ%6�W}+����5��i����_܄�gc8նd��\.�@��y�3'�1O����ONa4g�哦���t-�X�I�n��+��!	���-�#�晋�$޴��P�����`��L�����XG�'�DEz8��śE��j���!뵀A]o]Q�?�s����<���+ϖ�i���PFm������eb.e��Fn�A���sm\ޥ���x�9pw�a�G�kG�LVp��2�����I栉���R!M]J��_+n�Au�� )RG�L󓂑K�*�n��9�l�'KUg#���GXH��ft%���U(G������ڗ��w�ql��D�udx��׻�e-+]p�2�R���Z,�7�j]}7�]�i|D��+�A��ZH��)X�R �e�R2����إ���G�u��ӑt���T'���Aa}n���	5�4�UZ�Q⬎u��m��RO�{wc?����ب(x���f��l+��/-��z8�02��I]�]��{+Ti�8�W�	6�<5�У����R���"T�Ү����L��a�P�^z����(�Ѫ���|�{W�;�i�S �\��_���F� �&e�aڟ��fA,0�焎$��r�5���$��"d����U&TG}��������l&��HG[�_W�7�I�|�"�6�&oc�������͏Ń(ƥ�ä}�_�n�����yF3%w?A�q���+y�>�m_г�D���UW?��V�V�V�����j^]��w$O����IO��7Ä�Ǐ�3�ZZ#o�r#�tZ�@�e M�M6:��!�Q��J
�K^���݄���J ve|�3]�
�_=R������1���$Q��c;���~mLԑ�s1��chx�>ieӵ��>�W^P��G����:����xpTq�a�[~�����>z��sc":�*�8~���fQ,�Q��ه�D�?��/�U�u�DiJ(^.�+�ikY
�j��Үr�_�ǲ�\e����f=�D��ѯ)�Mb��Í�쫀�k��K�+[-cw�u�J2��#<÷.�7L��'�8,_������z��I���s4L�	ڈ_�YQ����}��2R�iM�J�[����c�I��=q�v�r<^9P��5jsѩX�������AݚK�!(�)��i����A�g�;|�����4__��|�]C��v>O��'�>V�S�wS����,��&���N��?(§�>F*�&��lD���Վ�ܕ��7�G���lO�K
I��w.���$�PO
��y¾�G�r.6�9�9���W��%�*�}�.1�
��ݴ��#�8�P�4�:�,�(�r����̓�t�LU�2H�?t+�mNN�0Q��
�BP�R��M����'_P�l}��4��e֙��O�4W]����"�ErǾ/���n �Jx�U�:=!O%��˂.~GD��۰m�D�{�&G�J%�:LSQ|խ���H�o��r��ݳ7=YgT����=�o�SV�Y�U+��A_��I�@XĢ2��J@�����r	�2�Epײɟ�(����g�m��S�%#�Ǫ�Z����
<�vO�y��;�&�(a����c�{S�h��,/%\�w�T�Y�r%�i�_l6����D���#�4(8��h�t��I3�mzd�D+�$~���әW�W�4`��_�T.Q"�T��b�� ��N�x�\i>�Y�-�P�{\�U�닉ŧ�����_��=6�>��n,z3'���W::)T��U&N���zCoҭ,>��+;����ėx[��fd�c�O$�C�DarSy3��g���t�+-�}9V!8�y�h�i�'x�8�&	#�{�hD�����P��xsoh\��/��#�]��=�%��W]���"���I�3=�Ap��i��>�_<�_�"M�J���S[���P���985���b�r���/ȷ{~__�<|�����i���͙L��'<��A���,O=8�Y�����#WA��	֡��
q �+�}�W�]8F�����`�`���pJ�:$�!4��Y�F��#��'�F)��<Q u�����^�M �M��ր�(�s�t#����z����*L�����о��h�#���"k)�77d}=d���P�T�8�0����b��P��oO���� !��9��%�W'=�s���0��s3�%�芔�O��a+��*��ט�Wv����3��玡1��Uk�n!���H^~�"6`y7���1��AҦ���3B!���2s'6�gҠzmu�gt&�K����6��`Ps@:ݷ��M�2I�r�mԚ�L�-X�P���?�zo=u���2�=��%͢ga�k��+����S��)(A��O�.�^)��E�@�2ψ���DmX �� ����ɚ��LZr���C�G�[B�;��	7�)]7�/<n��	@�����3�(�;c%�4͓k#��^���#{O�WŚRH�R�^�s�=8����g8��\d�$m��o�M��Y��dR�Ϲuv�ʾ��5��Mp��Kx��AR��k�*V�uAs�Ci��_�+F�i�N���Y*<G:�'�����
7S��>�p�5�Iޗ��D3G�TҎ���T���	l�V��������?E��Ф�&��z�|�8vNe�ۭ�X `Q�z�<Rj<���=�	"q9��9Zo��2� �E^���>T���۔�h_��=�g��\'C�  Q�hM����?罋� 	o̇RkYf���Ŋ-����A4��Y��d���&��f=���&����Qũ�,cQ�iaJmE�O�\&�ǣ3�f/�^+7�O[|���5=wg�~��<�w���qF��Ҕ���!�%�k����r�m��4�����@15�� ��Z<�Aҏ��иo���W���yXD�'.���(�=���/��-rwrh�xr�1C��Ay&�}z�Y�jV�>�8�ڌ?'k�G�i)Y(�`� 2���o�|j֟.�W�X�vp����N:�e��]���_�&>�B���K�~u��+�$XZ����ܠ|��㗛��6�m�X߿{��ӺX%B��B�����Ӌl�4ӄ�e��Y���Of�uz�m&��UV-9��L<��9_׳�%;��������� �0�|:뫬���ZW�_躀ʸ�!8�=F�]���Z|^�������RLe�&�(R�,�Hte�g�WC�/vT��Ax�ԨΦY�dI*"�E!��K�>U�fM+���pߩ��j�r�1b ��񶫹Y� �G;�r��+] =PÙ(B���9��_L�$���tQ�yֻ���d\�����m��J�ӊ`�x@#E�v�fAv��v�#m]��2������\��'nX�)��x�z�� K����y�6g=�"�It�.�ܢ*�𔷎@�9���ao�h�j��'��4L�
��nAɥ��SQ�<Q������̛�f�f����	Q��+$���j�\2��=�����mU{ho\�ܪ���i��i��PbyJ{������aG��.&���nS��J+�B�ED;8#�Pv��DH��l7)�\��m��f8�%�
(h�2r�����K:�F���_F���b��46�W��R&.=�1cb1�W}.����8����4�ӍV&�0��\����;jJ�6�66V�8G�_\�^���)q�xh9��[� ���1���W�4��Z�QU�oy��8��A`�����H-�����Q������%�F)zE.�6{�����3SZ>�Ҫ���`
�:O�d@�|����-yVI�KN
I�r)��	�sR^S߭��t�2&j� _h89\��~�%�!ԗɌ��(V1�,=`�&�mپ�[���\J�6�:y�Ze��[�����ڛRn�,v�oʎ�\]e�-�	1�4��/������=z��E��0\��"y^��$�
��v��b3����X�m	���]�� �"cN7y�����qJ��ذ����ъ$T#��"^�۫�V~���5����U�,����?�a>4���z��#�I���U� )�+48�E=1Bp�Ӫv��"kIIv�Sn��s�O1�:��@��i�Ok�̛�~*��G�u�W���9g=���������ζ=� i.[g��N����d��h��'����cm��8��X�϶͢+��)xɳ�œ���]����l�%�mκ�h�^�|�ULTDgNk��/��D��q��	�孤K��|�}ԁ`>6�J��9�5�-T3���P�ؤ&Dc������7hβ
~ߙ��O^w�Bw��ۅ�F�L$���G"@��������וT�Iu�籷�1�V,�8�-��`�^G����WL}^~6��X,�Ӟ�0��av�䈔dyL��[	�����r�]���kE�7�d$dPN,��F�;0�΄�)�}\�q��Ky-b3�L� iA \b�Mjo<2�����0�mS�b4�>!=ݓ%����7^�-J�lrс4=n���L�"�<����W��hʉoL�Z�k�d#���_��A�=��y���52:�)JAs�E��z�<ܒ���ڌ�$\e��(�7�̷L>l0�7k�!"�7�F{M�dsmt
}��(�z͘���2��P`;�adn����}>�f�⚲g��$���Gz����r��b�҇&��"�N��f�ٸ?��x6��آ�:Fo����\�X���rx��,�k��2���2knh���g��K��y���u�{��7̵٨�y���N�_A�Gc���{�o�7�Њ�)T+,���G�4���(��j �w��+�y;A_.^�W�(P�t"� '�T�.��wT]ƪ �4.�f!�G��M����Z�m�_��'�}<;�ǂ�Ժy�g;)�\��zt�uYA'��΃��k�D�'7��'���FU/eGE��$p�H秥��ѠM�n\�_Bb 7}g��f��\it?G�<�?-��c��/U�>U Ӂ����D���8��EUS{;������M^�X�v{�J�`� ��&���>�"���S;OX5�e�x�u��d����V\h����5�=`V���r�i�G��~-�U��%����1�eņٿ�Z�_%&���7+Z?��uWm��,V�}�F��NR:
lZ���P�5��R^�c-u/w03�N��in��y;JJ��)do>q%_��e�м\��z/Tg���xa�|x~��;$�"K��%��B�n.��DRPXcl�69vY�j+&����ru��v.n�&���QD���Ye�11ü=~��;���N[�W���h<�x�� �w^ �@�έl$��}�iT���)��-V�Q�{Ь'�*���Zk\�^��ִ,v�W��{���åb�r���sU��aq���J��y7ҢLX�K����f�ZWʗs�ck+��Λ�4��':���x�2�.�:k�f�ͷ��c�*�T��D�<״z�m����$�*��Ơ�X��Sӓ�˗ E�(����`"������8�F����/�W��O�T(r�������(�x|h~�Ry��CZ;��-�~�hP���$�h���U�U��<���s�c[�.1�W��8O#���L��W���eM��<K���6v�,���k��|⁺S�0�E��Ŀ�s��-�
��sx�,i�H���J���N��	�#�8
�-���:Q�-;b@5fA����3�����P��縲}���-#p)�@�[VQ��g3����_���}�2�
�z�y�,�UY`c�h�hŉ���Xј��_��������%<K��C��`�S�h	�-w�q�s^�:�YZ�&�3Q��+F_�?8�l���!��ѫלڹ��>_x�v*�9��G�g7��K�p������h��YS����pq�{�JE���Zl���ꃪ,"�Җl�w�rݼ�?fIF7lUn�a��5�ȕ��K��^B.�)e=��7#�H�J��-�
뭢I�����5(g&�r�w�O�,5z>�~q)Ƽk3�#X���y�~MY����v�~�P�E��Os˓˲��gm�y~�?��&��%8�M-�+�?>XF7<v��1_fqS�Iz O��gw�e�Ie�^j��o|�Nt�ξ�oB
)�5u��7S� Bdd����#�W#���T�q�e��HX��þ3�Z��>bb3M���l��$�bQ����n!V )��z1�D"!��/+)"�mG�
,�g6=&����n������Q���]sU���tZ�K/._�%�(���� �@��|�:�	'Au�g%��.���F%�f���W�?����r��˛��0���J���m���oP�E&�Mo;6XX��@��,��*��[�y*���L�,r�n$�EO�:DOzf��B^yPG��zkB��[��/��}TI�y��N�?��0E � *�#��c+���G^��$�{jZ$��d!h��%�۾e���M�5��J��gxdo��g�����e�{ҽ)�̊*���a��\���j�
5��\� ���P�ל1=�R<) �3�륗�=E4�5��7�!m#��V��H3\�L���Ԏ�:��_<���JjbQ<��>��Kp[���_+嚳eQL��o�AO�,_\�+��hh�_PJλX�)=~�=;�R3���`���s)�薇�!g��^6_��ꪚ y�?hK�Г�؞U��YW����:C`7zr,/�r�s�������Vf��$���_����q�p�I�r-A	��ƙJ���R%c�c�yV�eg�5H�j<��kK*����Z��1�i������^�R�{��dJ&�,O��B�c��Ǉr�+�e�e[/��_�	M2�n����~����T����w����%o�s%Kʼ~�T@N��No�φ��v��z@~�we���9���}�4��{�kl�_�]�+�e�����ͿIM������0V�&��������𵟌�A�~��S�D㬍��^�7��2%?6�a�uu�}��wnvZ��?g�@*��ƃc>r��=6q��p�.�a�y�3$�j�+U���	@fb\K��d+�7S��S$&5\������y �u���� �<�M='Wծ>���ݦ��~߽��q���9������;����H��f]��M1���.CA�L/�m���>�����vc}�w#�hn�H���v$$�E�� ��Wg�n�k����=�O,���OH�Tz�W<��U�e��d��SRk��fL!s���Ob�&���Lk��K{|�K��{���`��%�$�C�������f��/�F����� j�nRw��t>�9^~�R[n�fFE���i<�77:KZퟎ�ݦ��b\�l�`t���pvL�K[#���e�������ˀf4�ŭRr�I{7p1��0xd�>��z��ۙmh��~��Th,:�V�7Fwf�m�$[�ΎT�p�A:�f���������������^��4r��v��~�q��_;��@��~��������Ӱ�+��u���{���!��!��T��<�|��<H��!I�1X��%|���F�C���6B7�C�rG 7G��ֶ��~����y�2��<8���Jn�V�y$V��<.� H�O:O��4��m��Y����(�q�|J�����z��^��c3uw膡.�H�F�e}�Z��׌�騧�����e��䊧�_�V�����Z��ɂBM3s�9�5��yv���f�I�,��mk���g��,=F��#�<5���3�V�䲮A!�t</*#|4!AG��Zz�S �{B��1���t�_�N�z�$��\�I��Έ��Hw8^�r�R�Fug�M�&tYn��<;ۊ,�>��z&kN��ZG�KܤW��3���t�3g��?�G�<*�'$��]���e��t!�z\vs����B��m�@����هټ$ݻ鐶���w{�*ݰ$�u{z�]�x5A�
	��ڜ`]�F��3���*��̟*ۗ�F�
 �'�Jo<��_;��Õݤ�k�K>������� ^C���H����?[��+�x��
��V���Ǿz��������u�p�佫����X��hC5K�/��Zf�`p�]�?SAҷ�H����R�[��"`��_�FՌ��ו����$A�����%���h	p�����%�6l?}���ο��\4a+�b�㰒Z�<<�'�	����O��z���K�1�a@�]y�ԅi�{ޝ��t�,63]s���rxJ�V�䴼*o2��Q���"��{�=�V�"-����V�e�3�{"1�ہ'F�Y2t}���s!g�Xm�*m�$�(��*�k���i��/;h��?�i�i�Q�U�5�o��O䬇&�.'y��I�6�y�ٸ��Ug�6nP}p�W{���-s�n�䔾-��Q ���=��$&>��#�k�����{���dݜ#�����/+|_l�ǷKR�MJX�Ahu���N�[?���!�_���b:W��Bw�5���o��(��}*���%^���V�j#�/�˿�Wq-_h�n�W[���"�n���q7��>qN�׉��P"^�DF����?DI�"�u���������R��	d���VF��>�I!f����������ÖCR[�+2æs֊�d����Kp�c;�td������QJj��r/��;�ȓ 7&rN�?��~X5'mBF�s��e�=��͜����{������iH���q��װ�D�RW�~^����� PK   \��X��>}��  .�  /   images/efb2c8d6-2df1-4fd1-b4a7-6ff478b87b86.png��W����P("MJ�zA�4K�/ ��AJTZ��*`T@��.�I�MD���v������ι���?0�1�H�Zs������RWG����Q��S��� �r��0��=G`}5ePI/�
��(���7��p�<�
|�Q����J�X^W�2`v�una�R 	q;���Cb�_mcs_�#�XDz��̡����JFI�{��6��LtN�O|�oz�\��xec\�۾��_V������~��ϗ�/�0S*`=8��?$��b��H�9Þ]{A���R�����i����Q(�{����i7��}�9J��.��7�<�����N8��?FQ��z�Nb |S�?���� <�?�@��� ���;lW���'�ׯ@'�SB��g�(�����G�fz ����^�t��c=*!��(�xa��?F������A��ZЌ��y�0�VƳ��Ê�XH���y�F{^5��B���t\9�?��]��8m0��m�sU4�y���׽F���B�����1S^:o�:Ӏf5=��V����h�@�>j��L�D�lQ��K��F���Û�_������8��d:��UG܊��z�?�ۍ��J�|��T8ʮv|\8l��tRѻy�9�%�&ߪ�q���쫛�9���k0H��R��E���"�PG�W�dt����	��Ovi|7;<Yv �Rr�)G���HB����V=�tlRw��'���j���wc�xh	��QR&+��I�W��9J��C�'�.M�
I5Y��Q�s+o�D[D�"5y��.����y�����{�<<5Y�ƭu�WD#�x=�N^Z��{vR��dܢ����%k����3�后����=��ګ��L)K����{��q�Z7�D(�#��P��
h�X='�,"�8�={=p	�=ł1-�t��1Ũr@�a���"ZL-1�����'+��On�YH�Bsl�d����t�6'ܔ�nC;D�M_��j����ՂVd�R�3��9����J�a��X����_[eɰ�/J5�����0�6�V��Le2�,w�
�W�������%f�<���t���ԏ?\�V�ԸE+�B�K�39�����ɓs>���!d�>~DE*���P����Y�.?�6�X99��}��O\塽lF��������5�u�Y�p��*R��QiE��i9V���]Pk6���ጎLj�荍����7N��b́b�=Y)�I����]
?���D��0�k*b�����n��f�|#�j�ӷ����4�"����&w't/�ZL:V�'}2���	���2J��5߻Br�qz�?/�<�	B��X]c��Ȭ� f��������ϴ>��>���W�γ���̟��
m�ϐ'%'�_����ܢ��Ҋ��lj��_���
�+��	nWw9������'k����u_�s��u�S��0�ޚܐ`�ecC/�2e�/��1�`A��9D�'.xt-h|�mٛ���*��]��D�)p¨��o�z���|��H��0�b�!:�٪�=��`� gt�"%%���-t�����=a�сi�;&�Hj�~�)j�A��r�+���
1E�i��>
��{�I�v �J-���ѴN��0)w�c MJ�3GBHde�׫�'jY�>�>j��9(r@]5�A�+�ܹd7�wo��K\���n�R��Y��׉Ӓm����Xz�����+����No��i��-�ʸg�pn��39�G�vNb9�3����%鹆]����5_��zz��_"�|�n���5���Ժ(�Y�&#��N�`AL?��	��̞'f�a�����!����5����:q����A����y�]&���g>)Q^#�ev
���4Yy�a_q\bg����}�p���֊�)*o^IV�D���mȉ���}�.`B�A�N��s��dd�`�h��eiG��a��a�1?����ފO��V����k���nq	ݶ���M���-�{�?��������;��[�Yad/�h zC�P��m��.伻t��ʟ��J�����?�NZ\�`F�<.&Ls��el��w��fT�mP�Ϟ>3:V�����F�DYM/;���+�6c^�(Di���{�
��k4]�(��]�K%#fb�R}����E�K�k�i%ߪ@T^Ŭx���mԃ�x
����^��$�]��7�G�G���h���Ha�ٕ8}�&����v����2X�-��W����� )0�nB��p����"1E|KB�$�Y@쮩3Cx�$��s���h3=���=N��cl�ף��0�@4�m-W "ܗnaVv���&-d�5��<��Ä����
m~����vŃ����>�>�-~���$��vСt
�wC�T�����J-��p�ɸ<�Ʊ�	���u���s
{�b�}���?>�e���Hl`���Ւ�b\�_�*o�XK�@�8f�G#>A
�/�
fO���[�I����dI�+�GF��e���O~*����bT�?oV�/L?��w.�B?��3����n�7�]�	� U�w���κ�p�L�^1_��LŶ�j`h	LA�Sa����r�*��*3~N��rQ���w��\���=# 4���(�P3iQ��k"��t�G:DL]Ie��F�S���,Ϯ��D��/�3�[��J��6�oRғb��#��*�?=�r�����3��y*��z�ҧ�/����d�sXq�d�vy�y�j̶�Į��qXm�r�����[��I XD	c;w�����Sl��#�s��~|$�����'�֯he&�'*��7�<�:x_��ʭ�f��P-����9i�y�}�w��^�U�_��FHno����.Q}���i��t8Ќ�5��B3/��_\�Ҝ�!-rvs;�f��U����ֳ�����,!Pz���R�ɷ��ӹ�Yﶾ�T��2Ի�ۡ}v<�E�d�m�S��x�Z3ÑΒ�ӬI�@Z���1na�LpZq����_X\�W
$�u�B*����!���������#:���a������sN�j;�6	��@�D�0�,%t���_,(�|�UV���*�`c�-���{Z��k!Q���_��A��p@���G2X�)�ՁQaf�=I��ԫ�qT��,4�X��x���/QcqFvz�/Ց���*&7u�J�F����S�����C�V+�w�2��~�����fΟ~��K}��	�8AC�ݸ��}�ԍ�a�[X)J���J�	]�K�\���_�?aX�߹>��qMHtÌ��[�12��	���Es���@$&�S�%��M a
Q�îo5(A������5��?<�I�K��@�<^����Xφ97����WxJ�Is.߾���B��R�[:��&m�=�/��{1C�eoQ�ޓ���x1̊{�]����2x��Y9X?����TE�'cy/Jn�6K,�T_,^t�=ɷs�[{��F�KШLy��{?ȵE[�d>h��舡��N1ej�����X������m����L��L�FP]�Nɩ#��9#�W�ڿ��1��%5���x�[�I����_��jl� fזħ@�[���\�l����>�z٪!���Y'
2�2�����O����up��K������]
���2ͷ�c d����֖n[�]��C9;%�ߋ����O��bǮ�m.z��::�*�3p�ܤP��ϖ>U$�����?��c+���1�5���|����4���T����sx�;X�a�2����m��)谺VTW�Jz_���f����&[�KHE���T��;f��Rse�aE�2ݜ���B1À`�b;@� @S��Pr7{�~xL����_C6q�acǯ.�ĥǈ�ό�P�|+�D�x{#��&(�~���{cB{8��s���B�$�1t��R�mΓ:5(��z��˥����/e���RģV8���e[���|L(8"t�����U��)�,�8ݶ��ۍ��%T��_��z8�	�a�Y|�q.R*��t>ޯz[�'�!�%�������\���}��?��5�]PD�xҺk&)�-��7��R�^������~��$�G�.�0���g��4��R@��[^@�o���v�E����������6j��5����NW�do���N5%�<��JR/��Kk�ؽ3d�;XzT���J�
�~#b�=��HxV	/���i�m��)p{K�
#�N�ǥbn��L�����w0X��s��#���M��G�����h��#�M�o����*D+�R�>CŰM�'���|���>N�4Y��y�a(��/���۾&�MR�C��[ɫջ�?��Z �E:Qb������Gjڹ	'���k���!k�}ٲL~���pXr?�l\x��z�Y>�ܱ+�z�
/r�D>O/�ѧ�ge�\������76ޅ�B55rߐF���d�j�p5D5�D\�|��B���s��4L��T�z_t�g}xM�P�~��K����� 4�W�z��7Ma���d�k5����(-��� �ο8�X#Ďx�|m8&w���dȹ�#g�V���6��~]��xTw�C|�]Go7ojW���5��Շ[=���
�I��j��b^1��˥)v�a���{��>xe}�ל|]e#6�	)��b�{-\��{i��0�"�g�t��8�O�X�l�d��ޝ��YҴ���kIJ��Í���]D�c���Pnx�0n��w��9�|~�%�+���K��>)	OW�zS`�.*x!�;�T�t��A�4�bK�$R3)�kx��ߚf$ػ�L�P�2[(K��J��5+��$a����m=���=t�8�z�5��x���#���f}�b��H{t��%tm���kB��qS���}���Nݲ�s�XҾ�3�-	�PO԰��>{X��P��;��tr+n��EG�O{niВ��@�{6bsd����%}lmtR��K�FR�M�c�����D�{'��n46�;�(�Dl���mE�!R@<�;�����L�H�oT�&$�u[���bf������!������"��j�5=xU�E���9����gf�d���waK�^7�v��l/����Ǖh:�h���"ƶ�r�"6z����I`R �?�}AS�Eb�+��δ��a����A�+o#R9A��GԲɂ�d��s��Ի���>3��-�Wi���Ա
m��ݖ	�I}<"y����߹��k4��e䖵�}�+��cR��2A34H�H9u� �����4Z���Cb�3:�������)��篾�Tc�7�D��A���sqd8�@�����85^'�wl��|;����*
`��B:�h�u��k��^G�J�|Z�j��Z4�)3��+UWoH׏����№(��äݧ�
��!�QCP������o�9R����w�JWW�L�R�����Ċ8."�NK�K� �¥���N0w���� Ts��8�><T��Du��p٭���m��8{�I�Wd�/_���ِ��k}]�Y���|���s�����S��8�^(f��R�?Ft�����ړ��z��f��PVk��a_���}0����������e5�&� �q88�b��ڤv���I�md��&��H�[���3��/���P�}�L��D�.�y�SI��;H�Ay��Y��*��L���g��^ǭI��oݔ�_��mqB�*�K/rїϞ�R:F��7ż`�Q�W�#�t�%�q*��xI���m7�q-�w�Qr����V�{����bo��']�d/F\���syn�B(6���JQ�/k�Ӷ �r�dF��a�;�`k�t"���y��hD������2�� �����l6� )�VbdB�RP�./�u��«�oV%�T��55�k�F���^}2O�}��V�o�[O� 2C�����"�<,1R%�����>ju�tyh���Y��nw�֘KfP������.��6㇆�Hm���_Z?�i��5J��A�`&�pr�.i� ��)
�~f����P��v	]�gJp����G��'ι�A��k�����"2.G<�D�ob�*�7h�g�"K��f&��r����ۦ�M�.��Ó�����[}kp�+A�2%1g�9|�X���r�e��H��AG|ԩd08 O�i����}:���!���'�����cr�j�������KV�O�6>-W�wn�\�>Wc��h>�
�r�z�) n��4�m���^+��Q��OE���([c�T
�;�[��X
'=_	AH\dF���#�L�(M9�%��t�5��ʍG��f���~�G�,���b��~�y\����-W�����pf�����|s����bp�:���o��u�+��Ii���қ�Z�"/|?
%/�����R`,�>��2�.c0��jĘ���Fj�ώ'�-���O��y2M�o���	r����9%�?�QfEJ�1�NU3_���8��X�Ђ�8���o$�%0��S�3����Z��v9����d�����+H��2���
S ��9�8E����G�ݭnk��ψ/l�c��,�7��"'��oe�J��d��2�~��Ű��;�A�]�:^���@L;�S��%�;���p+;ӏ���P�*�L!�A9̥I���hU�T��S�3B~���s��d���F%7X`���=��q�}R��4��Q����*&%�Ȁg�t2eT��M�≾&���*dJy�L����T<�ur��qb�o:�7�-}2���O��Vz~,ZMÿ<Uaԑ���%J5����*�$��E�ꍇ2��D�L�4��j�S��&8v9�8�R!UN����+�ʫy/�d�ߎ�5�bd.�m~�e���=�la�h�i�FU���A������JJW�w�KG�~��O'WnT'x��'�&""vl8̿W��:�v�x����P"�9�c2����B�$B��>�qwV��k���鍺��W��>����ɗ���(��h즮H�b�?�^H;�{̢v���t��Pc'M��&��GV?H['�~�J�X�9�f��H@D�(ڳ���_�'�9uJS�J��d��xcA%��(YP���6]?<bQ&��o�5<�.(�^7��w�����Z9�t�Q2-�Q�ac�|-<�o9"n/������L����^ڑ[���O�����o.�Z�C���F@�2��1�hV?�����*�?�@H�%�싞 ������q0R�;xz� �|�ۏ�G�*_kpz=����އ]�� v��b�"|ˀ���f��6)�p�9$��g-+�>�~��Lbƃ�IX;�:i�����/r��̼�1���߽��"�_�=1mZ������T��,֢�ȗl�B�5(Dc��L:r��jln�>��O�i�4Ji�J�W/ �{s�����9}��"�R�����^�LG�4A,����ҥ�0{�����Ȥ;,QC�����Kj����6s'j��j��.�qH��
=���Rz�X^򕫞�t��-�ρ�}�Ӧ|�Y%h��y��y�LV�rB�q�n/%^}�Pp��ܦ�߆�M#"���;bXeuq�'H��3���a~�0�2=�Bn�m
�EvQ	��>��Iu?~��Pҿ��S$o�П��O��1|�W��%!}w�ǿu�Q�7�۹4gLջ��]M�#<�%�W:�
eI�~���=�{�?N��1�l�:a��h���)����.n�-f�T��-��,;���8�Q�
j �Kiz۾�i8!�3�/��T)�����$�UU	4A]&�Ls�i� ��\���\b�e�*�K`4�:��c�����}EP���ǳ��-�:���������o����Z�R罖+	��/�n�ܽ�D�:~.���'��V�G�/�s�d�7�il/�=&���(�S�n���}\��h�g�����b���`^�i���t� ��2u313��P�t�\��E�f6�hIB���sC	��/y���O����3Z�l�ʉ�����Gjg���h�\͸�L���a�����}y���|\�KQ��	�����K�&�^�vO^:1��ELXn|�FAF�2+w;*pR�?<�V�����!��s����j�I8�2
o�i�֒���r+7h����FF/+{:�#��N�̓�7^ȊS��J���m�6�% T2��]�1+�I I�*L�	QH!%%�}��nQ��
�������/x�wV�9���i�|�(�*���I-�>廝�8����%g�cA̩�����
�y��(
��P &�����Ƶ�>�D��YS��;#�,I)��s�{qS8��P9Lqi��Ue%y��)Q;��68s��"�Ŝ�U���$��!���r�;�ԛ�o9�ǁ�p2U3���!ۈ?��ۋ;��ݺRr���50�eN,���o��ܡ�¢�6���A������(���,a*`������Ʀ?k���x��u�)�ZSr2����y�����7�b�d��}E�JӃ�AB�Ҳ̗��h��� ��'��1���F�|?�֐=�Y"H��ۈ �@L���0�Q��cQ*u�0��A��l	�O%'�n�1�1K��/C) �
�ȱ�����i�^FX�KtO�@���E�X��D
��e�&H �'Ե���7˚{�hpŶ��)c�<VP�Cr-�>b��Q��F1g��?�kek+�"+6�@�~|�˷]�ܿH�[�y�^�Yj7첾d��QJ*>��,��k=]%�N�
���+������P���yK��jQAA�m�FA*`[���|�x���j�lέ��v�T$*A�J�B��o�����vK��ӧB������E';�>H�.O��q T�i�T���?D%�[)���]�./걇'�� Lc_!�W��E
s��Y-�DuG@�';�8�c`qb�:X�/�����̒|%�'�/��0JJҚŷO�o�޲S���pi&-��O�������(h܅���ޅU^�����mh���Q���+�,n�q>9�KF�)��<>�,e`��a��OQi�}C4�	%�y|�`�%@���
���<���V�4�,����</ā�ԯ�=��N��j��{��͆!_w�F���@)��'7�/ב�Ar�q'�B�\�̲�yu+��+�`S��NJ��_x�����(�����l��9W}M��%O�`_����Z�׎��m�x `ݵR�Kߧp��ɢ�<2q<��Nl�o�~ӸE/.�[�ҍ;�[<�e�9�m����F�8"�EQ�R�%MV��e�$���)Hrٝ��[�hf��,c�7z����,��U2W�q2�i�����-4�v�G.���pZ��P_r?���?�Vs����m������}=��i�� )�~IF$��=?H\�h���0���C���
N0q��K�6n�7�G�g�e���fr�&���F<��3��f�ؘ=2zy����Q4�),�%W�SVo�n�����K����k�^x<��ߏ$�أ�_���(���??e�����
���פ�j�R�-�Y,��[�Ck%#�to����[�-�VB���W
;+�v#M�?|�շ��-)���L*�%'�@,�ΰ�n{�ڢ�cV�{�⫉Oψ�7�S3Au���sC���lzb��Df{ǉ$"{*@�,�?���UL�>��=�,�)A����B�}��Phwl��"��VK�
Q$�P�Vtp)CT�B�Р��Mks�{�9��:H4n��>I�������*�̢��6*��#�/�(�3=Z�d��3f�~�.[t{L�Ȏ^�j?�ƥ�Ų���N��c�J�Q���4%�neȳb
�M��$�ώF����.Ց�ڠ��чR��Rs��l  1#�H�ֈ̰�?i����A�׵i������"d�Y �NѮa�Z�-��q�������%�u�� �
"��-t�>���`�g6�8�6�Xu���r�a����F�_&x����l�(�`��ђ(1�h�f�ba5S�1�=+����r	�AC�e�>�>��9�$(K����П�W�l0��Ax��=W�Aͤ��o�,�/��eG�:���U��%�d<�c�tu�qUy�|߃0���a:<���ho�~��'-�l��$��V���Xe��i5�1R!�u���>wT�L/���K���������'�-��,�=�:[�UEh赈S)/������v?$�V�.�}Y�|�v���3hB�ݐ��r_�ο�����gM�%-'+s}������%������N� ���<�N�<~l��C����������dt����|B$���RK^Ϭ�#P*�D������ ���.��7 �#9R�A d��4)�s�t�(��T���T�uw���!�g��c�^srb���o,c����2�3���Z%֋y@f��J_�P�`Y7���jd,:����sx�m6ĥ9u?IpCe!�4��ha1)�Qp�wl\��w�x�Sh71F0zX� C*]\�g�ؓU2?�!��+/���7�������#۟���/{_�4�"����V�Ć%�xx{�[�v����f��aM���L��'��;��"���s��p#�}v�҉�y�2t���b�N�c����8����ԟ��'� \Q���ׅ<��̎��"�AO!	(BD��)�6��@�f�>B�!�$)o[��+��s�]w��D:{��l�f�"��Zc�����8@͔!un�l�&#����R=���aL�	&�l���������>�K)L�p����\|��#��J�ݭD��4l���`/#�h�i��A�t0Ec�Ē��$\��m���A��5dcG���ߢ��i��|B�޹���)����2���|�����$��m�<�lɞ��ؠ�br���~F1�p�Y�����3��		ckC�n &�)ߤ��� �@D��� |P�!�������1��sy���p�S�T���N�Pн�i��q�{���	Y���D(m��e�1��y �hͰ���о���iG�j�8y|���[�8�J�:"�Gؾ��!qK~�E6�Q;[h��Mn����%H��KĖ���LV��L�s�;��w�� OW;�e�
�0D����gr�I�	�^6&7�1(h��(1l+�q���.�(�*�Hq�p)|�^Ds��O��%gj�R�j/\jL�W����|�'����ήU:�l��}O�	*�U�N#{�����F$u�قuӊ��M���_�O0f}'<�b��T ac��&8�>U���^<�X���ԗ�G���6@Gf� (���N��Ƌ�=�>YYN�)2�k�LO�2����爤n��cALjD�R�4@�)\�5yF,2rj�3���^��vy���\!l3:�P�w���CyXvs�i�+!��i�~��7Tq(�,�����/���Ċ�m��@���=���hךgG�`Ǹ�Y�==N+]��K�!v�lh���F��;����O������c��z��u����#�'IK�rbC�߰�����Ǽt;	=5$�O%��.ߕ���㍧�rpv��)��g�,�O;t����<n�m�.6�tv��6�o<����✈�~����Ǎ��e���{/m4m���cN��d�A���Ȇ��i��}�J[�<�H�j�Q�D��^NA�u�F j�%)�_�p�����+xU��^�V�ͯj(�UPM���
�[bj&��A}�v�ݕ�7�Iܭ{xq�G%܆��)�>��F�C�A��7ֲ.��`�N[�����+�V��c���Anp�WtQ��0vh�NJ/G�nx�Vpu���&<j}&k���2����~s�0-��|�F�����AX���td6)fɽ���"�"�?O,¤o�m�@h�R:/�[�|�0`�F;��b(Kb���(�6xgV����Qil�bHܗ]��F���.�PI!�M9��¨�,��),$�X�����a��t�D�xNVu�|-D������!Ww��&}L �<�b��$0g�����Bd���6Q�\ZTv�*>�Ȥ���J�ޕBC�jѐ�)R�^�� 3~ك��ڂ�hO����h����T�V���6�c:�^�h4�U�s~�-�	���sh��u�E�hH��B��p��n��Xa�H���ι�_�n�<cQ��I��RDC�*S��^�Wi9),�t��b����R"��.}xa�'��|�FP�,���?~���3�<]�~R�N��"j����0�#d����~�|k9�q=������u���9�C��>v�h�������7���ߢ�
Q'U8hG�& ��%o"�B���B��k��W����^�~у�
�b�#a�/�KYa,�:���Ґ����&�$-�*�=����̶Ƹ\E>�~4�ǭ"�$�>�Ge��e"��h��LU���IԸ�I�Yax�~���aL��%��R�񅅅�i-�g(0+5�a�8G�=%d���.N% �9���������>Q~��,���x� �W ����6'��ym�Ĺ�ȼ���FZ��j:K���h]��ޞ��o���63�۩��4����#��K~�HEo<w��Srlx���e��$p�2�3�t�mC�mc[bTlV�Q�,ibw����|A5P� ����l�ٶ��]Ȃ�`�Ykaa�}�.�7m�����C(c��J�y(y���A��9*�v<������{cayA^�Q�-9��#ד�A �JԘM��)��!�Uu�-�fNz��v)��]�+lo��@_����;k\>��.F��r��|t9Lά�<#K��#ǃ�b�g@xCEocn�HS2EK��}r��r�����,�Hɤ��:�L�m�S�7�� O��4�C��_>y�60$���y�/�V�D���s�#�m�<j�����yJs����`�E֣�	xe\&�{wIq�a�6j�"_�˝q�����=8��cP��?��$t1�m�_�R�ALR�GG�u�k����Ͳg-�~��u �k���e�$�=\8���ȩY�̡���q$�Xc����.��o��|��oUE���\�J�B>X������H�g��:�(�Gi���}��.~�d���Q<�v	�ZR�_6��CB.�<�b�d.����<fnR�a�:Y���k��c�Ln��@ӿr�"��������~��k�҄|��8Z�YD�Lh�]���� y�W�}��~Y>���:D�1�gFID�)��)O�C-�n�ͻ�}���A��A0��N���L ��.6���K���ke�E�z7ZOtL�S�����֯3$�IA�=�މ&�R�A�|��Q���m�i��i�@��w����G�jY���Z���$� E1�Zl�h��._Ω��q��q���Pݷ0`fU��k�2P�������\,,����F�ZuN�@����GZ��Z�L&�A�l��f��1�v3�G�QD.�%��A��I�Ă��2:X����B�%�߈eK�ߘ�Ԝ����7�%kyh-�]�k�O�]�����ױZ�U4���ˁ\� ��>-��6��E��[��N"B穒�{7=.~�'���˝����P��a��>���M\6����ۯ����MB �sS�6؝\'f[SI?�����%<m��7ޓf�^��`�~���Q��U�?�1�$�Ǧ?��Z�K�U|N$����Od7�L��;:��#�6x��ֿ��6�H��N<�q��{�c�jG�w_��?-fP��b����2���܉.��bS{�x���l�ɷg��$�u��¿D7��D�����n���:M&���2E�̞����Dy^����h0����:mp5���9�|�k��\��������KQ"�F�����_X���|��7�C��dU;d,�i|��
��\�/+�'j,�I����� '�,s=� B�v��/�3k߂���0�c��X�Fe�1�#�N���s�(-�J���U�p���V��l�v6���*R�N�Y��~���˕��"~�R������H���q9�f�`'/�V���l�������E�G�d/I����ᇞ���p������#^��DR$P!�]3��Y����k�y[�RFX�.
D��cZ8�n���Ƚ�)����'PW#�e
�F;GH�/f|N�wgMyb&���*�Gp�}>����2BH	Kh���s����Ў�%M.
ț���N[�/Z��͏��X��/�����T�nZ1��_E�����2��q07���V�����˪���VL�7'I?I֦|��G1���k���uk$�,�WT|��#f�D��Ԓ��cN��ڳ��Ye)2��_���k�%�5�n��2��*L�:*������v��3ҎokJ�:�	2(��ʷ�D=�xt��Y��I��8"gX����&�f
��T͊��$[ƚ��>M�bB�0g���7)*Z�\ʍۡ�2�9탲��l���y�����j���|�k�z����;���Q��������ȿ�*]c���}��:sqK�o�)h�]��8�,5pE�츏��˅�C~󆍀��s��M+u�{�4��7�~���
��m1܈�ԜI�>���_�P7X{7�~f�L5��q�|u蠫[�uvY�E&�M�wl��;������Շ ��ɰkܳ��w�b�S�(y{����6����!����'k�Ġ�D�6)��x�����*����,!F6�AE-���+�:.��'��2��)2�1�ӿ����X��)v�8IQ�uU�}]���ov{&p��4���o;kk������)9p� �����XkV٧��������cAGet�F|����y?�#�����~��-㦢9�vg*R�Ϲ�~�pM�zA�7x���ȫ�Y��w%9�����a�����&8����$h�ѝ#oaă ��,�L#`��Pb�7q���v���e���G_�����k�z���$*�+ac�M?�	ђ @�s��&Ǡ���ۘ,]j$K����ȥrw<�d�C�>j����^B�r���SX�WS�����g�^ۧꝩ�B�#��V͟�o<�viX.�;���>�� Za=�����bS��e����X�g��.�;��?��?��3��Pq~���l"�<��iBD�c��C�������Y4^�o7p-<n��@/š��Fͷ�2/�=;i��L�oϩ"*T#Ya &b�u��e"W�����X��A�Ǽ��4G�FҚ��dȥyq\G��ʲ�ԃ�E�&�`&���I��Qe�cY t�iiA��U�����s.KG"=�3W�
4}������B�MBx_M��L�>/�q=sP����
��F~P��Wl�N{��k�֔��]��,bAk��M>��M��[k��ח���O_���M<��K�Ɉ�����X�o<s�KH_�ç�R��z�����^���w=��r�t������` Z5Ԕ�
8�]+�����:p	r�j$�S�
!��ܑSRj��� ����JuK����a��cb�T���}��?�,��x~�]X�)@F �����&6k�;�?��ޚ �Z7vj&o��"bS�%��;�I�gdq�rx2H�"��h��}zٹz�X-S��y�Ӥj�F������l�aӫi��J��P9-�]r����t�w��N�ϋ��j�4��^K�����'.i(�f�,��L�Z�@q���o��뤲��y��mɠI<&C�x_B�.d>[�\�ar?� G�ڜ�f�-yaR�{�`��ܐx�UG��OΓ�Z�GMC�C�s��x�[ܷ�7���bޮ ����:xJD���ϱ�,�v��\@�ӨW�ID��B���)ݡ�8����Ã��#�٣��R�Jb�<�}noL9U�.��>��y�}c8�M������nZ	�7l�\,<kߪ���o��6ʊ}�0�aCt��X�!�Ek�=0�9�M2���;���|�u��,žjܪ,|h�=�)5I�����?�Bفr�;�b��a��!^�I�I���L$�?d�ؖ����G��X�K��u|�c ����'��!��J�.�AFl_��y����&>[�L�br��j��d�@��5'���A�m'd�ݣ>5H��L=�(�;��=۶<��k�̌����Q�&�ݕ�êM��;`�ah��;.���ˋ���?׏�b�\$�8�ʊɍ,�q���%�oP�A���d#��wk�$���������,�]��i?�d��>�_���o"PUu��U�>|���Vs�K�a��%[�Q9t]���D�ʏ{u`�uE��(��Ld�>��A��GSeJ���z�)<1T�$��y���~����%��e�$N���z��!Q���L(�%�2��/��6�L:��ٜU�4�`{y����z�o��f_��r�PƩ�������p��5bE�6z�_����&,����Q�v2��qɜ;y������O�\ �e��n�w�67>����ȵ���L�e�%LD��?rÿV\���v�.�j�#*�4��} �����ۛj$V��d>YjiI��7�sF�)C��@�xuE�����c\�k岙��WH�o�(�UIɃl�t�x.���*0ټ�α����h�����|Y�C.bi�]\�� �y����i��C~#�A,0��*����)S�	Ќ{ݷ̞ս�++�6q��+c�D<��~3���\$��l<j�m)���g�Y^���0�y ��^�y���ёM���_��OZ$�fx�nI�?Q[juF=T:]��ĩ��7H#H� 
�\ZþԶ�I9W�mP�K��Ё�O�?�G���Cv�4�mAM*@��E�u�⟋
)5P���7A &��C�[�Eս���H7�R8t�tKw���]C
H� -%50�H�t�H�;��?��2�c��u_���v�A~;w&\�%mHQ�}풣���}&��g���S"A�P�����:$���u98/5<a�4�Р�/��`�H;���0 X��x&���:E0`�-�a��v\yh�K�����7;�v����7"���Kd����|8]�ē��O�'�7ʴ%j�ꪧ�o6��ie�b�x��	4ks��d�Z�����!����Q�_&��*��$�9�`~��j��¼����Z�
]�P���[غ1�_D��&����@6��&w�B ��ΰ:�a%֋h�W,͉
�x��vp��> ��S��d����5���x,���l�ֲ�EG_ȼ�A�Ǟ����,����2� ɚ��e���3Ĩ�n6���z
�ښC�,[Ę�&�?%���Ц쮰�N*��i����G����J��?��E[�]7�$'�7][F-D����S�.V��������V����p��C�]9-av� Q�U�n��_�|<Cl8a;�iϔ&8�8�r%	0��&�_*�lP�}Jbz��O9Ԋ\©+�J&_���y0�B�]�*[��cQ�8t
*���� �s�v~'Ӷ��w��P x�L��L[�b<	��z
Nr3��1^�b��B;��R}s��F���u-%�M��)<��?��Hg�>��H�N���ZTx�W�a��~�P(s�1� �R���*#�e���~$����G���fh1GOn��&�7�um��2�vA���,���ϛhG�r�ؚO=�a�k�L��y�����)$'GP�y+H4�-��Lڠ�LE2��6wN�~��UTvTt�}���dX�ʒg^��������uk���?��f�^�ی�&�;0�YC�?��f>���5!���sω4��6  ��܄V�����>`�Su�*�w�R�䳲 ���O�fzhO(�_�O�!�ceR��u>���.Ngp�hb����1���w�OB�ۊd�����G��4��ߊӞ<nl��m��9�Q>1H�֥��,�Wn�O��r��Z��2�rC��;�ǣ�����kw��ٶ4��8`��XjfHJ*��&3��Z���໡b�Hn��Œna�fq��4�n�[]�d^�ӣx%�A�8m�09i�����/��8�9��S"5-f�b�N�VE�{WT��)*K�sH�gO
�p������� m��^!(���O�BMU���+=�ʃ�����y+��JFw��^�)TnO�T��l3{�[z��H)�6a���j��$Dт�p���Nv��@�d��`"3�e�B�<Co�����fJO�E����\{ؐ�
a����G�tk��G-p�ۧ������e�@r�����ޟ������0����]_lD�~�ih�R�3��D��t��!�eP��k��+ퟱ�����ul�/@�P������������5Zx�z
�oSH���J:~��~uT�*���w�:������QW��� ��ӌI��ɦ��wPI���3g��� ��Ѥ'sm��w5�(�Ko�|�e���1.�k0�d�[3;o�����ъp6�yd 1�V�tV,�
��܌�A$7_J08�͝�����w�M����1I��n�5����Oȵ�d��+_�q���l<H}U��]M����MN��A�vݯ#M���r��z6����]�!��mB̈��}�ߗqڏo�^i�GKf+���5�W���vܒ�H-*9��A�L�X�����t'�w�3�S�%���J���C�4 ���WOP�X�Sa95M�,�sp��R��"iy^(K [��=��V�J��A��L8f�3����K����ݤ�A�q�����k��sЊÔcM�9a��|WΨj�F��M��������1U���L�j�&��A��'}Os��d/@�\S{3��pW��B2���.f��~$k�^�����{̏�&ĔV:F0mX��/���k������z�瑾�/�${���S@�����7�6��X�Qŝ|;���P�d�-J[��!w~�<3Sv�Q�˥� hg-�:������7�'�f�!��\���p�ĜB���9=f�7��D��%��{����#/�|;�.O�8A��~}���Q�P�d�%'0�j3�ɗ�qR�L$Ϡ������y|J.<H��ܰ��Ӟ�շ���=}a�g����amy����Ԫ,i%y�^�,y����uOr)�z~u6��o��4��x�R?`yv���9���.��x��*��(��` �iV�RV=>��Zd����f0E��*c��o����D���G�
!���<�A��U������%Ŏ���+�W�(�[O���~�\�|[��L���=ƌ=u9�eA��v�<N�o����	e_	wI��P~�9*��C���oͷ�b�࿃�8d:��)�h���L��	��w?^�!醞v+?�}��Ab|�H�1��%ǔz=����_>@���`D/�}t�G!��	��y������TÄ�S�f�� e��k�_��߾;�@�aJm��s������vS#V6��l��V����D�`��%�� M�>v�=
���Hb���ӹ��y�'?�4)����7�eD
�<���t������0ǂdp�w��~�fJ�87,E��xr:vƙ�Co��.<XY�$O��4X:Xs,hr�/;݄E}n����]�R�G.��먌`g�>`��sB��^�*���/��͎�Q�W9puCh�F������' "�X�!�p��<�z��79�0dP�D�]p=X3�w�)���9)�n�d�Va?|+U+w�b�~��DI￲2����dԬ�V7�=�7�:߬��C����|'~g*{�� �ߒ����͓�#�J8QK�ă`�g�Ďo��b����O���a���.}z;��(��a���xy1kA�{��3�~_jA���xE��L���ї28�]�/��QF
�^Q�6�Xxf2��ɪx���F��4�̄�%j�K�k;8�%j-N��nr�ҽDv� IU�*�y�D��o�Õ 
J��Qz��hH�o�\�^�N�]��U2���F3��ؓ����sW�s�G����N4�Jwi�@���ף��D �({l�t�WؓЖ]W�r��qj��p���ׇ�H�0�c:��c�q;u�MR�� V�Y/
)U�<�0��P���x�k�|:���K&m�<����7�<\���5�!Z������Z�~i�6����S��|B��X�d ��9���5�$�Ƿ�bZ�3�8J%j�`��<W�G�H�Y��s�/!s��뱄�Jm�{:�*Y�����"f����Z}]]߮"L�.`� �X�8�����)���Z}�d�����U�Ě��V׼(^�zp���\�PDZ�{�3n�dD�>OZ��eAyxs�X��z,���`�q3g��=L�C�3�@9����;��B�	�0�ݜ�<���R%�(.�O�01�&+ �+
(���zV�d��`,@�]r�~�ۼo��bS��UصP����p��\*�w��w���	7�/��h��u*�/���5t��E�3Y��T�ߜd�P�3��=��M>�9��ĸ.��6贸8����R��n�����Q��S���&�JsC���=P���DR]E&���r����lr�pGa2ƒqw�׹�le��JY����������Y����!R� ����2du4h��ٵh�n����q��3�b��e��7���N����$�ب׼ۊ��o�O��`���sR G���&�Q�H^���bh&�0��e�����bf_��&��bŭ�� �G6e�]7s�lV��&Ϝ8 �����]�N��.�G�]Q�g�N��d����v)�r|�C����4<9��,2��=�:�aS���!��r�)�?�����~�,�cJ�]�RE���Q��;�9�6����"��j����ٿ{4����Z��7�w�y��b[mGA�tO��g�}�T	��g����8s�~��7+{�����f�B������ʉ�*~OX�η��N�S��1	?�+��������^G��DP|����������w���D'k/!ϩ�g��1-$x|+���0s�Jh���A��ZЭ��dj�(�<բ��=O�����^-�f���Hq��o~^����`ȇ���^�)<y;�S�\���8�[�U���s(�r����O�u�*O�d+e�+ew�B�@�i=��2�Z,��Z	5m44��c��@��R�`��Ƅ\�3�Z���r۽Z�ﺁ�G�]E��C����2��;�
ޭM3��)|w?�JE l�8?l���iLiZ�l:�
>��7
>0@퐥E�Q����O+vi6R��\s�$V�7�����Ȟ�% & �\��]6;v�����t���R�^9����P$(d=q�?���&0 &#U����C��q��H��a�ɦ޼�XV �T�n�W]�pK*n	��	��Cg��'y8���ۑ2Q�g�+�	טd�b���;�JS�Y!���23B�2�!���ـ�?�AL�������2�X�X]�`�l��o�^*��Ĝ�w�$o�MQs�w�����M_@��>���!x���b�-����.�S�`�#�Dq\��+LK[{�
��� ��ώX�Ӂ��n�@J��	�wnZ_a�;ܮ���b\{��.>���:�X��ʟϼ��*�a��\��">}�p��'��|��9g�G�5E!�����3�J��[ȓqD00�vY|�z��5��3�oi��1� q���?�v~RY�h�L���x�
��,�`�tQ��"+� P����2�Z��{��F���O�՛
Q|���^���=(�w�79�����{�|Qx�ϼsᓹ	�T�lA����5��֢������lz=Ty�w)���:��?xp~��a�m��x]���@�yte�ت1>P<Ƽ�x�|���󀋣�C'���,Εh�i|�h��>"
�Ř;��쏓cG�X\4�S��.�0�&�)t���HK�tǽ

FB扎�,Y���f�{��/����_'����`��R�������}ׄ4q������Zʍ��e�|�
���K����mš� ���?� ���IpC�P�hg�J�B�`��zo�LV!�L��Pa��慻/�Tܨ�B�z�4y��=�G��J0A���3��i�`Ri��Q�v01℩������\;�d�0�.#1f޵�(@��� ta(����7��P#4�t7����1�4�[ߞ�`5�m�A޳,���+��#�҆���-Y�4��~kJ/Q�hi��	�i#ĐKR2ł�I`	������8�7{k�i��nm5������YNJ�o���:�[��=���]�-:�~�7k��^S��:�iĢ�Ŏ��ެy���S~��!�r�l�x��Biii����&>X��? i�"��UX��2-,�ܠ4�I��Bސ��0�Y��tQ�"��b��:B/�C�'���Ju�y�~���vA�����@:A�� t�h���4a�8+�Y�{{osk�뻲��Ad�o�H��!��.n�B5�/���v�|�t��I�[�M�o�+�{pC�+/��2ȍِ,*\ç1�ߣ5Iqi`_��%K�ޖւ�Qɀ`\sA,�V*W��q�_3H��EC8�S�ƛ�7#ڳ>��k͚���Q�r����m��7Z��Vs��9�a�<��xHtb(��&\�]~��^(=[��Ė{���[K��澍��'}r���,�~o} c2Ǫ�Z���9�L4��4pNB �u/i�PC��&!�*71J�8�:{��:hk��Gq-��j,}���h�B�e3;�=���V\��F�	[E>A( �u�}�d����P�,���J�.����Z� %��'�(⿺-bN_6a}��FnA�����k��n�]�;_��i�g��ݹ?�&g�ZCk�$��c�
�y����)�e��*tP�ZA��.��X�J��Ɵk�6ب���I`;}�߷�3zn$�Yv��6�%�d0�b�b�3w'�ԏa�<����*Y��]3ፂ>���nX����Ɵ��I��r���V���A,�	IK��U:@Z<�Q��Ut�A�5� '�T=�u����-��|+_J�2[��4$���n�P{�O]�1a�SYX.`��m87v(�p��	�8���5����K�Ѓu��k�e.��p�!0*���!n�A*t��J���g���jϚ>���Z��x��x��)�R�����$Q"W���j$!}��l�Ǡ�~.��f��y*s]�@�����T���bU��C��� #���<nH�O*[׺�5���-�l�p��k?�9��£A�4Q���?Z�M[������˗x� Zꋭo���Ǐ�����_\T�����>��H�<݈���7�m�  ?1�Wp�1��Ɠ���h��3��X�Q_�B}��eq;�u���b#�X��\~}
x�1u ��vQ�S?�2�*S�*��ܤ��5�%I�*J@чr���w]�uƧ����7r�O�ήO�Ď#g�
�lUur�WnlV�B�d�عfD���r�q�J��&X3�� CQC�6��[b`��A�a���\1ފ%m��94��V�߮R�s��G'A),��N�X�;I��-�B�yξ�"�faR�Q%����hJ�:o��\��%��մ���	���G$���_\ļ<���'4�et��ֈ\\�C|ܷ�@P⑕�|�ͪ�}_N��F�W�E�X� c��	^7�iGH ��Y�z-�)�*�K�މb��xds�QGǄj�0kD<�O8ޯ���O!�c�<N0k��|�	��J��z:�����J$�Z�m` �@2�{Ij��U���`�nh<��K������2��L��L����w�2l���Xu`�<)��=�y�"+�U���q�K@Z���I��âi�	�y�������KI���t�I�h���h�����\�6"���+2D�:�"�5k͵lő�\^�;Y����p�2"̍A&��2@h�G}����:HX9�������
�J�/s�1�A�q ��]9S%Ƙ�n 2�mZ񎙖�G����A<��E;��Ix����t��MВ�ס����g-��(����<CEK�B�S!p|��Iڨ�	���:븝z��4<)NJ5æ/���_��h&Ӿ��^RU��v�������|Gw��{&H�MN��I7������t��)��+~i{�G���X�R�R��|�����H��f��H��l{y9�L8h"�����&\�ڇ��������D��:88�����D����l8��R��ɠ���\>3��!�.�@W}2CB���؜���[Q����q}�N�1�9c@s?�h���^��j@��@����?ϭ��������j��yG����,���g6j��׼�߼��
{���Y���&�
���
+��ub�m��r�^MU�
b��ijN�gQ�L�����ٟ-!�$�[�T��t)�y`L�����"δ�Qp����-Py�h�Z����¨})�
�H�t�G���E�OLd?؛�M�=c�H�4l��6ID��5-B��!!������^k<��Ց���8���s��eL!�l0¤�{�P<ϥ���A,�U_'����yA�nB�u��o	p���0��.)ó��C�j5('�V����5���}�n�̐O��rT�Wh}���I�Z��r��]��\��j�K��i�f�i�ɓX!���]��faۧ)��uLV�G+��v~<��q��]��ff�]���hK��tź`��	��Q�}�ފD�����#��nb�ި��z���ҳ�2��:qC���2�	�[��� #�� ^=����R�@O�R���5��T����K�$	�x�I��GWC�}]�D��\F�pv���WS�jQ��Ј���1���<s�H����J���\%���~��]�"��
��뫔aqZSC?��U�v�ug��Y
��,}�Lj���������J��έc �s����l㬉��c*��HǢU�0c7y�YTq�+��ƆYw�q��?&�Vsc�.T>v��Q ˕n��4�F,qg;�'��55=]WN-����n4��m��1�U�P%�K����h8II�h�R`���݀*b�n��R�66�!��3���^s��ۘVz��ag��<	Y[�7T����=C�q$���p�r=A+�2,b�
̦����0�jrf�O�&TP�kmv��FI1#:�п2� #���Up#�0vX�A�M۷>��t�]�u�*�!��#j���L��5��si���7�1y��V.��a^��
*�c�����>��<E��ٲ���ԉ���>��;k�ʞm{$�4	h5��}�q��.������Wk���H��n��KM��&a��Ec�{O�#6]�Y������E�J5��Ҹ�8�rKmɓ
�$���}=��}��֗��;��\h�U���	�e�ڷ�X˴��^�~�@����t�x|~�����+����K1*܎UmO
Y�"hu3�ry���ܚ�={f��)xz%��ƥ$a���kU�afN��ds)�������q�3hP�[���	��yr��9%;B��.�b��Z��@�C����ux���T���RZۯ �gK�AN��1q��c,��F� _yrF}�7 ��C����:��܁x�o�'DQaĲ�	�xқNxEs��V/�����ޅy�vZ}֠�2�8��q�a�k�ٍЃ< Q�%Ĝ;�2;�o,Y��>�c͕��\�~U�}�.q��k�[�2���~bb�N�����P���e�2�W�}��"��qG��>w�n��1�~��L��������(<z���9������()m%�"=��nhTk?�>�%19����>��1��bI�&��Htm�hp=��l*�����w\4���� "��Kˈ�� �8}��{�ZjÐ�1@����)� m��.�	�"�.��\�E�\�#�Y6<s:<��C�Ν����^iX8T'C4����V���$lOV��"O8W��߁���m�{Fu��sc�ƿBXˤD-���t��׺>���֌����Oi�����&x"��!��qk�r
ꯚ�q�9Z/�*���A�|��?m�\J��}�"[''.!�����옒�իUUB�4��,	�y�YL�e�:��C�=���Q��ӵU�ׯ�(�&,ڕ�'zE�3���Bq��mH
����[W����+�1���ɕ�w?����$�@�����Y�^�d'��5�������:ACj�5,�q���n�G��Y�u3_��)����N�����ݽ.�0����!�If���1A�,x]B���p�A��P�[��@�ļ��~({z�HC���m]]�O���u�p�i�<�u��ѹ
�%�P[��ei�A�@�F���Sˋoߛ.�?�b~�5�p_b���UU�:UU�9N��a>��/U3�tE���;�U^���^p�����Z�wxu�������&�t������h�1�``lL���Z����t��u��|�a��9�c'�t��d*}�,�G���-z�<xWd}һF�5�˭����T��gO��E�#|����ެs��\�&��K��O��vzR�9 �<�X��w�|O
��z����]mf��԰;�}�X��	?��x����S���B{����7�S�hy���<2��ҒKe�nߠ����,�Rz�M��c"�'������JW勮�%���b��z�g��55��8�؁���an��O�$\f���~����ŭ�U��0�fk*��%������N9�"XK"�Hq�DWD[m��=�S5<�y������a4���w��޿n�vr=j'��t26;��ך;>oڌ|�|���AL�R�&������4,���ԄgF��͖�������3�+.�G�=��=E�RJ{ٳ���h� L(�${��"�����͓�*�f�x�\�'��u<*.���p����s�R����^�㗯��s��.6y"�+
=��˒!i=\hv���ULo�Qq�"'pl�����4brS���1�}˭�RF��q��`U�9vԩY�d������W�?��U6�s�'�4vvw1f�����'���y�t�.B�O���P���^(S��փ�Z>	S�Xq}��ڭ���a�AH�%C�[<��.�G�N3��\��,�X�Oϐ�O���FEJ�A�M����L�:eA�MM���&�#h�h`zB��Y�nF?YrN��\�*|8B�+U��9�k�c��[��rk�o�o�r�1I.�S$S3�`�:��)�W���w�6��'�X����pc�+1A��k�,��,*�1#|���m�>�9�����h��nB\]���bM�'�ݠH,���}��ِ ��`�9���\3*�p��jB[�	��!/]���E�ȟ:@� �	��c��z�+��+7���t���o�"}~��7t�h�y����&�������H��æ�k��F�#��pm�I(���n�mK�A/���6��^�1��{��Y��w�m�h������X�E���M��<�����s�痝���,��#k���I̱��埥���h`��1�A�ӯp͜H�����������޷\� ��A�P�X�G��ys�������^t���V�9��鱯�P�2u�d32��?��r�^/��,p�sA�Q�[�c4v.ʞQ2�]'�t��fr���y��Y�l�Ж���J���ql�RQ}�mէ���bM
�5Y	1ɱ�^��!H���"�Q��rO�I.?f���;ܕ���Q���n��B*�^���Q?�wT��Ȑ�<ĵh��znd?g��g��v�ˬ~���U����nm��Ы=��v_�`VD��sW �c�����7.��P�7]���_��zX�
O&o_��QW?��.������ꠉ�E���4'_���)�E*��!��X(�U`|I
��b�Eˆ<0O�GY���?HG�!�V�l�K�x��$�~�>��"ӳ�����
2���e���&b5������C��NvA�{������c�Q'����G .ڝ%_���Z�K
 *��I�Uɦ�0��2ɔ`��@�"bq�Sd����5��6#�`�(�����C��]::ar�T��L�}�JxX�G3{�᲍|w��#M'ړ�i�;"ϝ�� ���'��S���5DP���pj�S��<��M���ǢY�(�'�e�;N1��l9��^��m�C�%A٥���������R����V3ˆ+m���mu���<�GlU6\/7:U	?�0N1���������[iqy���X-���Ǐ��r�`KE���v΀�Ix���9Ud�UA��z��*M�g�o[�oL��&v�9^hL���,�n�*�}�:_0���"��|k|�˴7r��ik���>Vc)�hk��b�G����A�b��jP?�\���<�H��7���^F�{���}��`����mapVm�e��Ɖ�д�%�aVs����_�p��ݷнm-ҡβ�s����H��Ӽ��_v���t�����"�o�M}��a�ō$ѱ��f��n ����9��&+=�g���ղm��PI:	ƴ���K>��I��3�慻�rOv�@����t��0<�|J櫆�_F웾�5�#�!�t����g6[�f�Ҟ�#={�]-�G���
 ��pX�9�X囲�2��~r���>���wԑ9Ӫ��m��l��	q��,��Z�d{�\t��~�;�\J��9#Î�L���f&\$�{ʢUy�]<�@/��n��?4���j��4�����j9S�^jU~�t-�' ���Z��ݡ���l�H�8_p�RZs�>�L��!��CG�
�G����_5��O(m�**�,��Nk��'��hp[�����í�A�q:�B�����\�g��1 ��k�o����Z����Q6����(�Ŕ( � ������5X<�Y�ݰ�}w�B@v3�X|�G#|�9�>Y�q����x̲��;��ݽ*�~W-~v�q]b�ݻ�L�)�hE@ת,QP}_���/���X�'�u�<��t�kP^尖�'c�s��p�v����.�+�v�m��s�k�Q����!�?� I���则3�u��C�z?��fHRb"�oߎ��"o#ھˆN�	s��yr�<��ͦ�����~��{�(�pRdzS���N�}-K�^|��^������B��;?�O>�8��S��U������YR����y���myE�]��G���M�HA^�?��Q��I4Gq��{T�5F9� �����c��-c`Th�[�/.&�����uMc�o���͊�R*��QJ��X���Dx�oE����mZ,�2����'U؈���,�1��q�5�`�#P���n�;jTq���Ȳ�Ĕ�n�]8���j�<��7EE��y(�$��E㼈5.:.|�S�M�1������#��f���[�S�� ���ϕ?�Y������R�j����R����z��gq0#B'�y6���N<��]i�O#x�N��9��gԴ_��@P~�&�3��%�|�Ҕ��������??�F������ə��LEl���ׯ_gk�Y���`/�|Cy�l�ϟ/��ҋ<5}&�cyY�E�����Pz�eDS49�׶�����A�j|�5��f�ú]:::�ƅQ��)))�53��ƳG3��?�%�3�K��Dwww���1�'�ݜ�w����R��i�X(sM���e���|���Do�R%�*�� �_��
���acZ�7�������lS(����d���w3-./��L{����ף�v�m����89���G~~��k�"F�z$�h��DTTd�
�ڟ�}����@h�6���*�=�#ԭ�9v�i�����i��1t���5y�K!��5�����:'���O���|�u�up8<\I�؜��VO��ko^�lK��m����ʢ���ĢJ�V���9���Lp)-ՙ��X�z��H⊢=��4V����֔��"�$R`%rww�ߍ��V&K�k�B�Rg�Tq�׍����&c������SyC���H�O��R7Z6	޲��x�s�z)�PȲ,,-uM~�"}N(5�����Q*=�Q2�Y��u��Y[;|��#:�\\6�-�*�g�����w9p���0�����
��n�@����8{���ޞ�	�A�3���5�ʏ�Y\����̄Sv�L�n��s�Z���<ecc�&�r՘/4��
A�����o��q��HEU �� �.��@�=m��STDd,�4�l1[)��ɀ3^}�������!��֞��l�y��ɩ^��^��G�d�?N���%I�
I� �h^��-t��k�G*VyDA��ƳR����S�ܸ�����j��b�Gѭ�����[6/<jݸ������'�4��eI�{{m���u���>�q?��~����v��7+�~��3j���ڪ�+/�&LM���xu8��2�("��sg[�*�)^ v���Dh PR���mұ��{>i7�������C��8��8;[�])P ]�+�>�\s��q�%	]�`iD�D
��Tq�~rW(b�j�P�a��X����F̄:銌��I�"�u���V:4%��3�xd3~D���xA��ȤB���&F�{Y�r,S��޻���� L��6"�1]���aE�Rb��A��� �%C��`�#%��>��I%��^��P'
�11�y4SXAWIkL2-
�$�#r_Z�t���X�M�����zx���@^�H�|�%ݮw�Y��m�} t[f>�+�d���|K��˧�����ZC��pf>n � -Y�
����I$��c�f�7u��uZFQ�2�h�H{]*�ϯ|N��x�ʲ|����_�]J:�#+1?�f�����^�\HZLO���]�x�|K���� O��"�l����}���1�Uo���J�������o����������I��o��{�D7}/�`5���Hr���d�]�9HoE�q��O%T�OC���ꅄ�:K��	OC�f�7� _S "�������ӀY����ub�D����LEF�������׈�V�a2�����ΰ	C�������}�I���p��+�A*���ԘR[�.��pQU���|^��e�E_���a|�I֘����P�[�~�4��Ĝ�G�X�>[au5R�9�"�bsJ]�B�v��i����¾��I�Uu�j�
Q1���h���������r|3=~�Y69n����8�B��Ԫ�8�Ņ���۹	Zu��|�2mjTnZʥ��ɳ��&%B�o�[��Cx�p[|��p?�������m�m�]����QНGF�A��b��w��{_��)�v�)83���2�ǥR��n��\������e��X �:=��x˄Ý�"���l��xr�s)�GF����{{�Z�.�ת2�Gx@�N®3�|�a���0����͝�g_�;�B8�0��o����m��Ǆ�$KZʐeT���R}�5d}1@�]8<�uF����߃:B�(�Q4�9����,����?�[��H�<��/D��3�
n2A����J�LM}Ml}�ܷ3�sr
bŁL��~�9e�\�+��o�LX�&�6:ܜw������8âv�䲵����N��'���7�q"^�X5�1����3���Bgܘ!�:�av>�,���7N���B�)�@ѥK1�\o����@�N_]aݔBh_C�v/7o�y�k�sz��?O!�.�Z�;B	���=��&Ukm����ynC���&f�� ��~~~=����l�����*���[���I���=G��P���%�7�巸?W~:Z�>1���� ��l�T�k�p�ت{�Dt�J��[�'6�jC���w��1c"\�@Єu*{�&�]���*n)#�)q�}�ɼ�~��ʲ��K趏��9d>���m�]ʹ���Nb�(A<���7}ik��^"�Xș���J����A*?`��BvUV���򗇼NuY��%q���ˀ��ӫt%B�H�y�J���@���Ⱄ���?B�C��7t_f�kS0��}�z�����e������%��JW0�����E�u���������:d��9g��6
�)͑��icŀĂâ�Db�����N�5��Ah��ÇKicc�׫B�?c�"��Oչ�d�E�C;�(>w�s�� ���u������u0�<c$�SS@�D
 &"T���X�sO�M��Q��ב��&�[�(Eߘ��.S�7���ӷ2��[5:�9��������������9s�sgӺ|	5�Qb<Ak����nh��pw&������~��V8�ҳ��r${�w^�:b�����p9(���#�A���9�5a��0�i�W}:��cx�݈�72L����o�B�3 �ά-1xt�_ۦ�Yo�m����#	�ʖ��G��.�F� ����]��\�4�7��ׁa�aIT��Y�z�|r��jk<�}(�22�����F*��;�}}铯2=35i��V��?Xs���@��Y�t�����'Jh�l09�/�Z���o��_��� �%��AN���Y���^������2��2LܠK =� �O��lV�P�L�����_���ʔ�-���%��U�\g��?��Kv��-�Ƽ��EXc�b�̔O����f�h$
��Vjp4�2uh50BǢ  1��4H5�}��`�D�TE!�N&��X��l��o&�O�F~����= U��AC�����J�~c;�}��
�=�y�>�2�wǲӀ�Z_�]Dr(M�.Y��u#�2���'�R�y��<��OQ!>�Շ��M7o�3�����������+B�Dmh5Zm:8����X�����p�跙Dn-�:��?�?O��[��<ܝ��vFHt�����5��hZ�Y�R�'=�溚ۭ��p| ���Yȫv��4~
�ۧ8!�x��RH�Ăv��g?�.1�sF�	N�X����.���Dn���C,6њ��|��ֳ�.���G��e=�h���oY�m|Hܾ2�ު�%���ݿ�&�V��V��Y�{A�srq��lh�E��1
rY/(��3�56W��I���ExL�;\�H�Hbbb��O�}i���?rPg�`�݆���U³Bi~���pI%%��]���<����32E����V�R�7
�|Kc�J������k�Q�Hh<D@,��o�B�/>"��V�^e3o���o�HSjo��<|������2ڻ}*lĒ�����1��r��hh���*����v\ r8O}~ܨy����S�MXb�k�����_��/_v�c*��~�:
q¹���(~��|���ϯ�~����;a�ML� ۓ�j�aT1��W�2����9�Iѥ\~_]]�Ъ�F�L��YdC�Z���_�ct�g�,N�����Q@/�nj� m�6�qP@9�HFEF�t��Z]ݸi�3��w�$���ŔG��Q>>�( ����I�+ub��锫��]:w���� �	/)k��%�U6yŚ�-�4�M�n�B.���6(z:����9���n����U�#Ifu�>Q���v?�Vz,bTN�r�?��2*���"�%�-��)�ҝ��)   - !(=t���"���9��s-���9��}��8]U�������8Z�N=��#X�u�޲��ku�e�/s�Q��'e%|��c���C��2���h�YP������J��%KʠU��C��JiP��:3��_�yu't��� ~���X�>9�V0���z�h����oT��Du܁��^���{�y̔����1t"�jҎ>���-O��\��ѧA���2,��]�w�ص���I��á3��@������u��M7m���״2�j���b���ʼ����	�����{_���XI������JWy,�Qa�}�caT7�:��H+�.ueM�#�y`��F~�i@m�a��ɐ��0��zߡ@.z�Nf��VҔ4Q�u�Y{�y�rQ5g[?5��t73���K.�m�gY�uC/|IG������,���L�?<�-9$hQR�����c���.���%�������מ(tɴzƩ�"p֤^��Ӡ"5��C�]�D��!O$��NVI��ǻ�M
#�lz5�k7�ji-}_Ry��/4���C'-y|э�ᵈ�2��dnY6� ]b�wh�rJ�9^	���̈H���!s��7RCx&U4���8X㕚L�<�b#Y�<n�5-T��K̴h���vƩ6�M��sA��E6>7�Ȳ��g!�\́n�_b@Q�:�l�H8j�ˮ&ʡ��>�W��c�xa.��jj����{ �a�N�+�4�Mu~���Tm�/JM-:L��M�[Z��O��Q*�Sb-���/0���R#��m���4d�&���oBt$�P��n�~���'�=;���E�ak���]Ր�OJK�_F��s.�C"�-?dg�ǯW5&��-ׁ�R�� K�}e	����rW�~u �p��(;y��Z�߮N�t�2����1����i&-�v���z���7U3\)�sy��L*ް�i�4��'x:>	'�d8=����Z�|}��17��#��+$���],�`�㗃�ߠ,��� _��#{����ʓ?��z8`^,YWO�z�������׳D�f|������(�ZW;:���f�	l���j��dy|iW{���T��ѕ@�a6�[~zb��?��9\T��\4�ڵ�0j��nb�hH0���b�C���ĭ%�����k�ј����jl���°#��48����uAK5J��b�cY4{;������ikн ���U�?<�t	��(��&���4"v�h�
�^Z��/��ɣd�>{�tӃ
meR�6�4��fԊf.�]��%@��m��4��3u%�L��x�o�{������d�*���r���SY��iA�0Vpє+�Ww|�ڽ��z-���<0�/�E�'����(���`��@��"r�Yؘ�,֠����"Sr$P�s����krK���Qy��!�.����8���b�nq8S@�"����g��]yS	�t).���{��_ʜ����-x+�v��b��n�X�4�W�8 �����>�*`�n!�af2(���1(f��
P��]�0+&�m�I�n4�d�b��C���.Կ��,�����*T��~�:�7�\�Э��/_�r�r7����;����o�h>���I�����������9�r;�O'�?	�`֫���7��'f��c%Q��Jb�:��U*p���5&�<��Q0(##τE�h��,�h'3�>S���˗/7.BCA(c�[�vv~�^����r;���������)�h�=�8�lj�4���9���xY���糝�l�r�|�AU���_�<������ ���־(D���K� ��P�bqwPO�y�{8�k(�i5�`*�.D�299��"ZO̍�[�Y��B�sG�Q�#�0�K;�|�5�:�=F���L--�WuA���[H�Ĉ�i[7��1=�{�o٣��r��A���Ɣ��X��������$2�$�z\$�I��qr����Av��w2H=>H>H�(��:8��tt��a0%�kiq���Q%��Bmb)J�Gu���ڬ)��R>�����2s[�@��Ah%�ڐ��X4�S��m��y8��}�r����'Ko�M'�a� �Q)#.�̿�8d��G�yv�Y�x�5���GQ��y�[-hV_2F;!Ǒv����r}݀*55?�Ś6E=V+r�*�[G$�L(ߑS��)�i�Db�~"�)���."_���܎������0��,11���� :�!�����-�b��W[[S��?Q̆tr��Գؗ8�E���<�O��?Z��~}�jV��)F� ~��I�;�U�+-��(U=sr�V�{Rg���R�V"�hd~�֬��Y?�S&�Y�绣vX��F�����ߙ�"#@��X��8�Б⍛5q	����a��n�
KPåM��R��K-�iݜ����F\6��������>.Ů��v���BFYb������4� �H�$B��A�d�� ���=����G����)�3?��@w:|�&�̨�q~�Ov�~qOnn�	3~�󊿂,�t�)WK��=t���u��*"�6|��^:R���j�k��SOӝ���A���2�@��p�?c�#�_��c��H��d�х�b�x%��ʝ6H5J$J�-��D�z��BK�;�!���� gݭ1~��ʑ��@������,
�nܰ�Xl}|������e�%�k'\���4�����|L~vW��y�=��<9�E\PS�EHq��G��ÆooXgN�r�ܸI�) b�|d�2�kF���|:��Wln�c����_A)J�͆�Fz9i�"dZ�<���G�A��3�r1D�RX�Rʩ 36vd�c�p$�U�u�j���mJ��-����.n<	`�����XoDozma���~K}{�!	f�O��d����.�0%�#I]Y�T.&x����yA�����C�{_v��NmFaٻMuאw�@�?�$��l�A%��)ה�,�7k�t8M��"������&毶������4��ڱ&6q>K4·<�jE�Z���בp�f
X����a�P\s��� ��B"�Y~���h���"�k>�^�']���J")>�i�&��Gh�?�i�^��5��>���-�O_��t �]�t��O�f���K�I�"�E���#|����VO�6g�L�P� IG^�_���kg�R���4�V�r��#���ۃ�F̘�|�Omՙ�k�k	��A��[�����pڏ2�o�:'36��ZK;�5 ʩ8��2�WL�8q��!�a�UK���P/cGW9�1=A?X�	l�+�0�n���ļ�(��/�^�5#��'��n�H.�'i �m���I7�7��fO�>wX�<�Kd�?�w����/(���[���/	Ǽ�ב�K$���s�����G�)��K����FGGG���u��@�[)�^>ջ��2�D��������qv���J������Q�cdJ�O��M | �0To�f���~4�mv�-���o��Z��N/|D�l�s�iH���%8Y�س�.�:��\`�������p-�Nk>2A�[$SbC$˼l�-�ml�R�[o��W�K�U�C��\-���]V��V����������H��) ��^����Z*_�<���'3��4ߑQP�Q#�����d��e5Z�xB�w<�AD"�:9����k`=qs�#s�к��|�\�b�o8`���,E���[�Ja:��~��N*vB]
R����(I���ɩ�⁪y�q�*�.�o$=X�7Ro偯��-sx3�V�vҷ-v"e�/����^�LT}�B�JOE�MT:$H�1f#j�A���Ч��Q���W}��� �>���]7�S�e!U�T0��O�4S0�Z:�sd��'�@���^�?]��%�O3����cL�f�l�'���QV�r��&�Ef��Ԗ��g�t�9�q��n��3��8�&+���pEq<{]�h"0�8�1��i�9��tK��!���7�5����effV��ߌ���4����Le�&F�=�nklL�rN�����9���:�}9;>��]t��#�p{��Ȱá�*��
�E�|� ��J���M;����k���ڸ�)�`�z�u��UU�.z?1c�]�(t}�5Xr����pc��6��>~�H��	�_D$AL���wM��{e����q��B5�}lʄH�s�æ�+>b�U����w�+�xuK�J�ȥ���m��^WW�V���K�;�oØ)m���U�����*��Q6��2�P `D$�
4%�fDșO_�ELs��Or�X�@���Ei��H˕D�����O�E�(o��:F�C1]���W�η<�I>lJL���Y"�[�x9�{GGoO��+qv87������p�s�6�� �%G�k�pJ
�px�������<���S�y�k������Y���ԥQr�yI��]+j͚P���T�T��*;é��(���R�>��S��]K7A�5bg�GW���`{���46���J�����!$~晘��C^�X��a�D(~��)ic�)��ٳ0�����j�'+e�3j9�]NI<����x:/l��i�\]�v}��O��<;;� so�<\L�-Ķ��3)j�-�?�?�g���4����XSP���~J܈5E[Z��M�q�w����t�4�{A�K�a���?����]��K�-#*$�R���^��v�9,��9����
���i;�����8U��� �5��,5��9ݻ�Y{�o���������/�Lma�����ʪ���V��	��vY�D���_�|twQ��z�L�F�?xDP�Ӛ�"DV��̉�ԥu���'+�F�8����%�t~�i�Ȋ����N~1^�l����`�7p�C4]8�	�AB9��\�潆���+
�9���(|�_"���W@Id}
M��>������kU|XP#�񌀮EA��@�jU:��I�E⮵
���1�^ab��] �466�.,f��e��1=Ɂ^%Z����/�H|�!�e�K�h>���!����ғ���D!�a��C��p�%O�n	֬:�C�"�e/^�������F4�1������"-V��w4���8d�������_6�`l�A
b��j��zf���g�g�%3�ZS��I�<;*L��(a���C�%�`�q���ѫ���׫��/Tb��h�l��W�m�t��0cp���$}�䭹���'!!O�Fh��,�B��;ߒ�_�[�w=Ǐ��2~s���g}O�pc�H
?dT&��� |#����lǀ��%�T4�����kp^��*���^P�5��t�@��t�m�U��_��8s#�V����D1g���{�kr�1�'�o{x|:Cy�@�|�wD�����ѿ�p+Z�9�I�`&��w������
��[���O�}t�Α���F�Y���X\�XjQ��뱞�F�R����4��-��y�~�tc�1��-��#��'	[^���<����������͙|U��o>.�( ��6|d�>;��ۦƸz��u�e
�bM%x���FFF���5� �2H���!>q�V�WG��@0�3S���NrA�VC֔�H�7��H�蘟T���*Z�"�g@����� ����G ��zU!%Y�&W�QX�Rx��=��_5	�t	{�	��0�E�`���K�{���p4�gT���)�>i�5��{�K���U��U�/��B19��-�K�đ3ȥ����:eh��7��W(��s���wk%7G��)�>3�<P�-���\���-_�A���^���pc0�e�?P^],s��˺�1>�ý�[�D!|6���>��o�kAD=uu�([\��G� Q�k<�5�l�-���?r�,�P�P�p�e� \�ʸŷ��`�}�M �ݿw���0Lq1��N*.f�3.˓�}�� C���ڃ	��<����#Q1�:�v'�=�2Lӵ��KM�����r���~u�̪����-���wSc�`\q�N��w��l�lB��zq���b��г#O�t*2���'A;VI����7��P31A�����Ce�V��T��-�~�~��g����eP&�бvv欷$RӲt������%�H�z��x�� J�,����Z@�J�,J��K��CTjA���Z�aUwb�m��Q�(!����]|ݚ'��L@i�%18f;�>Q �8l�g_�><l�$r$��-ƷN�:R��� /ooo����R�p�*K�A��~ˆ��|F�T#qw�'Wy�>���.V�\9���B���K�����,����M�*~)Q�H��0���P��ol@����ź8�-�}yq1LFJ�k
�e�����^�e�ň�U�<̞��r�A���ں�*�*��ጉ��{����y��Ly�S�uTİ�M�{�	�%I�cم���-��(}��>�ǾF���JQ���dL�cP6J��
Wa��: �>���;/F��@�?B��v��^�r�~ &�bud����ր��4]��J�7���%
�����>�k,n�="�:��=�Bs�V�x�^��f���_���ʖ)��R��U�ktA[Gw�8����5C�W�u���(Kq�k�`�i#��HxvrR���v�����-v���WDD�P�y���j"f�&����D���j0�޽q�2\��͉Sc�wx�"��	}��,�)����m�vt�4c��LKy�̙j]6��bn< ���iX�f��Ԝ�Vf�>��5���U�Ya���U����o�0�,N&eh@d��{���t���M��Ae�N�=��u�� �!{K�Y؟#���&��W2w|!��	�JG�M�[�&xЪ�T��]�����犇�v'��r�}�L�8����G�x�)�B��1�;Q>���}$�l�.��2+��o�p��d���w��r�B!��W1���sj�,�n�Y��r���t�6}�w neB�L+Z�\���r���7;g0����I�|�zDx/ڰ�Vq
������R����T�m=?D�:��c����XC��ڨ]�C{M��ȼڮ	(��$��ޛ������?���?,=�}.�Һ(�w�����.a�Z�]LL�B6̷��$J���%�S�=Y�9��UY�A�s�;>�O�l&����� b�YU�䟹Ϧ�pc�o�a������]��e�����Y���/�9�>�s�QHM=%� Ғ�[ہ������?�n�^S��� Ρ %��ўXfG+aOLs�~&q�3_2�Vp�_Q�ڵu�\\;q��s\i�����vQ�Cԉ)��o�"�a-����J���'-ˑR��确���'w���̹H�8Ҫ�Gi�翈B� p�b'<��Ѭ@G��N�;�� lV.��,�L��П�_W_�T���ji�Ѥt�r�Dwt�i�-PD��^;��p���}^%���߸6TRGg*������?��o4�|�w�4�&�B�5q@��� _�olC>w���!�h�u[�L�e��l��q�Yc
��3��u?����<�CKQ`h(dR�^]v�ZH1��W���H̔�8�c)����r�III�S;wp�����b�[�c;�H�h��ձC�0 �w ����s�z� -�ޟ�g]g�E�8\f�V�0%:���t�?��*&&fz�Ӻ�HT&����e����z��t�8�֝�xL�˷R�^�:?4<<,�6GJy��`/�GJU���V�@�ש0�=G<��ǻ��I/��q�(�E7c]qY{�M��o��u�:雉^��љ�D��C�n���@���8���ϵ|���/sp����[#�r*�Eя;;����D��(K��J�,��V>}|�B�|TF���v��|��ĔCj��`F�]�l��ӭC�a�?��c�C�>fP'��Iv�eƗr&"A�
 NA�6|AZ�mϽb�����u��\�b�V�t,�� ���E�A��͞�xB{�!�_��;~��9J��<���D���	��#�-�3�u��<�/d�#J����HJNC-�c	~�4��P��@��0F��2H/��]#5k=`��53p��!���-s�#�y�;$�'��7��T�g��t�}[��G�}:�W�\$��/��Ջܔ^��F��M;�w��@
n�5��O�~�}ǈj-��Y5w�3妵J1W�cHy|����(�$����Tg�p��6�t*��m�H1�t�s	D����(Ƶѐ�X����B~lg��O�B�cc_�N�`��Q>�F�{(��ս�Ǧ���kc��]D��˥�Ռऄ�-����Y\���B_K.�F�2�ě��f\7��R��[��Ŧ��/*��)˯�ܵ��bO�?lw��0e�_;�}�qX,��tq9�}�z�7?}�1.έ��x逑&ﵚ�g����C.��`��i�G�N�Thi�=�3
� �����Q�'K���:q����iD~���I�<k����)C�>\ ��4Aw�|�[
p�M�x0a�iԷJ���پ~=ι��-L�Z�Ö2`���bji���cT*Ǡ���K����gM�e�VT�OLLlF��	�
_mGW.-�h^ �b��ۜ�0���#{���<U4œ���a�>����G�F�w��+��3!�E�C廂q[B�+x��m�c[	j��-������&C�\׻f�ߎd�og^�;eg���1
H��nɕm�����[�W?�n����W�ߑX3��f'�`p#���!�B��JE��"����H��K#U�Iصr�	�/�}��d8FSѨʲ�;���=��y�%h41����R)m���w����Xz������n�!@��xyz��F�)�;H}�j�?���5������}�k��1�Y�k�TrK�6>�t�m���h�Q������Mާ`:�(�����t�'FFF��lj���a��f�}��66��Uc/�7����}Q��*��:Y��(U��ٍ�bѸ��3Y�����vb �������r_��W�.AvUj.�3>rȥ��1����@pCĤ�!Έ|���@a?U��(Z6��n;e
�.ϛ�~�{�쭘>�ɹ9���#	��_�0Oz77'��D溺�_<��\(�Z�c��=�#~����M�w�qaI�_��zfQ���8���	��yt{�{FM�b�Ư(����%.�m�[n���D �b��"�=lM Ox./,,<��-I��=Yf@]?�0|��d,U��p^3UVޭ]�SVXR4����T`��U�Y�^�2�DN�P��?�N�p�3 ^a��c��Ų#�x|D,��J�F��Wh����+5�����������$�	��r�$...d�t^dc<��kj�\Pz��]J�_�����]�"����ֳ���[.�F��
��&���� X��*4�h���h%���$Yw�8c9wwB8�B��M]:]'
Z����lLxY�I���f��6�}�仴44r��u��Z�E|ڌ��1B0��%�J�ׇk�aIn�E1��\���	����s-�GF�:	kD�ƥ1M�i�":"�9g�6�����V��҇=ޯ�>ά�Ԭ=�H��M�h���I8V3ƃ��=��߿k�%D�rG6fk�%F��ϐ�et���!��峛�ۻ�`�����D�	Qy>��W�q&Z�Ǻ mX@��{��JOZd33�Ϫ&%&�N�[�5rs�!k�)�k^���!'2B�7-�m�cI�1��[Y����>荃@I^uZ��p��q>{�x5��i�^�Ω��������y���:S0n�&��V�`��輖.�zXCF�M6�W���fG�����y,�}�e��[��`�}� �8�z���www����bA�.tڀTX�(�.�Ux�v+`�Ǉ;j�M/�0L�˞��������Ņ�KV���1�&VH��U�ｋ���I�_K�Kڊ�omK&�i�A�����g~��������b@��3(�{M�؀E����InR ǂ�$�f�-����\?+m`G�G��qw<8�f��B��kN��lT�[��<�x��"�G
��+���,��f���#~�����F�^Ͱ9s��.Vdڈ=f���}��ҷ�]���=�8TB��t���b=v�o�S˴���K����H O#�77��^(E�L��ss|d�mE�����z��؉�([W�hY���DC�ifn.�X_{A�E�����x�����W#�����ES; ���$T�l�]kL�7����ox�ڗ3 o��g
1�K��c�W��h|�����QgCN�оȈe◥�QT�]\��,����N��Y��+�-�^S��"a���.f�|���<g*���H�ݧ~��s�R�w�wb�^��oX[��0q�|R�mj�M�3��F�6�q��/�r�"e*,�1�1��R;V\-��%�E�_�	��O��'*��݃7���v���E�ŉ�/1�=U�����`]�^����s۞�'/�p�{]�&���&S{�?��
Q�����Q
��A0#���a�U�(O�k��Q�~١������O*�hܑ�&��)�Tj��^�>[���u���$����2���!XK���ew�X# ��e�H�B^�\3�������h���3Ȃ�6����/�=�ט���f�\��ϟ�`����������!'oQ����ׄ��M�;T�����a�	J�
�!��jP4��U$\����g���of*+�_ǣ<z��
�'�i���}�D,4����^�k��	\������_W��V�;m/�;�Tmhgo2���{<<!��Q1*��M�"6����a(�������3�)�a���\u�ν�Я���:�'��2��/�������+�u����ć��{E���(8T��K�[7��Z�2�Iuxn��+�"�[�6}֙ȩ�z{�G닯�'J��C���^=S��n��x����%?�Vv����QYa����#Jrr��	�����VU�����&�,��Ŷ1u��1 �('��.}[$��<{��N7�D�9P�;����_�ЮC<2L���޼�ռ��i A�K*���G�L��}� >mY;�q5$�2� C+���`Pl2I�6G�-�mC)�E��Ө�ro�3�hY[���C=��{��7����& ��g!
q1RuQ\��&�,�+F�iP��q�T�	���l�1 ���mf��{k���N��\\eF͛�_�S���~c��Q��ñ_�1T�j`+[�WQS[Z�S�����m]�
h��Z�g�ށtɊK}g ]&=��W� b���w���L��݆�:Z���t����(s�a2:F���Wr���^p���sb~A�">�d�pѦ�,���˔י�Z��7?�X�s���<5B[(0���jd!¿Ņw[�=<��"�5�p��`),�Ge?~�0T���n�>:�tk4�D��VH�~��M���[N��oF3ᇓ���0>��㬚�%)����f���,�.�QA�_�x��uy/IX0�����rT�ux���bo2�c�)�$����aC8�,B*�ۣ���0ыo�><�C}_۽���t���.�|Dq��T�F2U�P	����g������B�n��/Eh � pK��V�dXK�_':0U�Z_�5��Ǔ����Μ]g`�7x�D?�'&����;��a݅��SRnD���n�<�X]Rb��{+��g�1D� Pe�ayT3o�9���{F���D�%��^K���񝀆�Ǹ��B�@�t��Q�	�q�7�	��5������䅳�"Ñ�/�٭����`�!�a�R������$�/���;��=��G4�P�:������;8xڃ�ݩ�������)��N� #�e��{�!���Ӆ�/�-F�rb��zV� D��DEE� A��]wpp z�ʵ��ۘN1��D��0@_���b��E�T��~J#��PM�[)�6��E��״�q�D�?��l��!�-L�>Q
{��'�=����?���J���}���WRsp��2�g@�T�x1��y,~Vzm=v���[7�c^�|�cc��V��8�=��̊�픸��'&&mF�dM {���z�:�c�{j�����X�F���M�>���ʞ��7g��ol�������X~t2*���C�\�>�o�k��S��w��W��.�'u nn!�Cpt�`���V@vn���/)��u�T�}���o�0�!�E��c4L�n~��$;U�^l�87$
������l1*JJ����9��2W0���b[���./ev|����4���*k�Xj'�}���a��(���'�������3Bd%��<�FFO�|˓�`����XPf��vv��{�ìJ��\g���~��Uچ5��������XTX������/��F2��k��,�M��o�o�_ӧ[{��gҠ�~��A���'ؑ]ೝ/&Q��Z��3�>���Ғ��Z���6���\R�?��y�, Lg��xY:g��aVkq:'�I���Q̆��F��Y����a�T�¡�3�p��upnXʐuu ĩ>8a�8:��1.]��u	���2�V�*~�"D8=ġ�:|>&o�45YnT�~V�:�2�G�.�m����Nf>}�hj!���i�ag�"�dIB�����{d|Ҿ��{<r����B�M�u�m�&uC�A`N��������0�i[�IC��du!���W��m���k�:�S8��޾�>��Hdqxb�����}��ѯw�f=�/.jA}�c��Kt�0u�_�|y���Zc1p� -;b��W�p��O�P��~��5.~�p-��3�R��W&&��-{��᳀���������f�.�/��(6�-��`�_�3��L�D�!���?lk�����AA���h��D��=1v�x��Re�(�sO���7��hW?x���BI�ȮA<�ّ��`b�8҆q_U&t�����.a�e����[@.���D�Z]��"[�=}�.���Z���.YDk��t���n�\G���L�O)���n����`e��s9N{6��sMU��]�^��%��E*���R{��@f�< L�j"5�#���@��v z�z��K���9��D����(���dBW�$�hܗz�o��O�����s�uؒ��\[`h�T�ؤ���I"@<X�����-oLu�+�n�Ň��(�GtD줛`>u83ߠ��z�2ޅ�S�c�B��R�g9=��+Q\�H5�����sQ>����;�kNy�:>�˂<@�T��:��O�A'l�x�k
>�M귴ww�Φ{�B����ϯ^R��:aX��spe�%�d��3㣵t�<j����?!l�&�g�Y&��-FU�'N�l�5����pŸ����L�\���O��a�6I�e�jK&����t�.�
�1��Gm��'T��r�/.�J	&'#k�>�
�Id�����-��T=#�kt�%
8�_v~�
;.C��XH�m��q��7ޙ�\�����券,�3N;�z۾��H阓�0F��qv�E���F�����ΡW�޹W�|;�2]����$�Ѿj2�7������a�x���Dg\���rv����!^P�ɮ�|�7��ůX�� �(��dje��p���8& k���`�&�,���j����(�����9�"��E�#�f
^��5i�Oa�V�u>����_o`�X�vQV���?�b0B��`�l<�];�ߥ�b9�{����ʬ�x����{jj*��ɕ(T��\����N=���2vwv']�i�b�W�=��5���������G�HQ����lN��]�"�*M��x>�f\!�{���^V_���@�DMI�`�5D~-n.�M%���p|U__�<0������3
/�LMM��9��dN|�U�t��#��ؔ���bz��edd��ztA�G~��>�ğ�
ښ���8�-�K.̴���O�^��5�#>� �Q�OӒ'�'����Z�A��Ş�.4���������*T�[Z:�@=�x�8@̡MMMA���L}�K�\M�kz?[ �r��/����v��8�N�_RH^N�>��ؤ�����Xe�o �㊫/�*/��>c�A�*�mʺ� ۢ�{��WV�8���w�L<}��}M��P�w���S��p����?�D��l�VL��ծ��j OmLOv2�wt|�-H3�ͱ\�I_S�gD8��d!��
�S(sX@
D[��-��蝊'�Wm#���Lgg<"BH&O�GJs�r��<#�������|Qقd; IP���I���8�R���y+ů���*���#�����A�n�-It9�Λ��p�r��d��7����s�����.�#T�K�5���'J� ���M�W��!��� �3�Ձ(�&%���?T4���7 �[������V?JjM�k��fg�K�=��s��dC�/M�[��*?{�yY�:p�gV{b��x�7x�TY��K�B�W�W�)it��g�B.j�v��M5�'�r���A���@]��v]���9���Дk:R/u>���Ǐ�ϣOE 7 �A�={p���o%CNN�"Doe���0��Ҕ"ۘ�S= �^do�T��x��f�QIurm�{������͹uw���`���YۢF���a��ODۇ *��UIH,Н#��!�	R����zt�~Vx��#��I��7��-����Yc�OV+z�Ǔ9<6;;{�W6y�(0�>��KXدvp��-]�K���N���_�
R���������:Y�r����QD�Fc�:��CVE�#m(�������r��[�n/R�
�p��������D��j)����ڷ��C�����	؅� ^IS����c��rM�^Z�}'���ׯ7���J���/8]��G��9m*�R��T�E����"���l�=�_�h��Qq��K���p��K]�e���KC��M�}0�J�Gש++wss�hxx���~v@	����RI����:�Gl����'(��Bl�m�W�c4��1�5���vX	X��<ǅ�瀱��V�ՍP��w<�E� ��(�3���<�H�GY�f����gP���j/ahU+�.������ܓ���V�ȼ���5׷,���7��r��,��n�������vov�r�Ǧ�����JN�&1R�̑�AVc6| �feyN�]�\��5e�҆�G951>>y�/�eoXgV�ޓ�^`}1x&w��a��AK�y��鍄��"�>�*��Gú~�L{O����������8���s���'�^��a����r����@�27�7��pe�\W��\���A�i�-o#�N���K���"22ypQ�Յ����h��;�k%�T����;��q�>sp��uuk̭��-��`��r�:Jv�H����{G�FU�e�SS&e,�vs:�y�M=�"�ˀ�qj���w�����n5g�N��3Cy��GB2�p�+&c��p-��N��~˗���63�Ņ#]_�oe��X��EE�Ys�ށ�T0��/*����I8K4w4������+�{�Gv��6���9?t�B�`�oL��E`�5!!D�	�^�Ŷx`8�9��׹ݟN�`04mЊ�é2�SM�Tv�E�%:{�
���u!������cB2��vN��i�"����*J��K�o�k��0M�ɀ�%�5�K�'%�Y��2�/��8�5T�]Z�)�;����"B�aIW���NY����Q����Ft��o�i����B�͓���#�pi�PK�D�Q#����`��'K�x�'1Sy6�do1ۗ�X��.bbbK�W��΀a􀺂~�'NZr��ɨ�+p8�>�HW�2�� 	��j>���X�L����i|'�;2�3pR�g���@�)��I����6��X�p��o?p7��i��Q|Ǎ@X�/~�P1u�0SaT�iS{ �]\�M[XK�U�9|D�X�l�r%��%�P��6ϽɊ����!Q>Lబ��TP�x��Y�#G��m	B��Tϯ�ڹ�v;[[�����* ��.]�Ɣ���
���{��\}����Z^�9����	����q�%�˛����t%ܥ�\�1���4/7^leu�邥��K��)�xpyxx��� �!�����M��%���,��D��mX0��S"�$P|)����9"���O94ZddbF��@�/����eZz��w"d��['>�Tؑ"ӘJ�ݟq���ut���0 ��%��)��v��W_/�ns0;�G��'��
�`�%�@�)F�u�.9�C���\��J����5R7j���T����LT6���̗.G��Zz|�@����<LO�>�HaM=j��(��]��j~��z0�fO��r�}F����s&�w�aw�I��Ɉ/p��z��Z�ʣ0���~_tv� �?v�"t�1�.� �<uds�ч���^Q�����U�[DI�,]��� u�I�� ��d��1�qU��d��K��ɸ~.�����w��$��#z�'^�"U2���������8$�N&wt`��G��Tɏ���U.:�	�;�U�%-���/[r��Wp9]$/��"P��c�73���[�;e7bӊ����v�5itڈ݉c�r�<� 
������ozH��������GD��/4_��@�&5Ԩ��'Y�9֏"=;�1�\2!<t����k�c�����;�tA��AD�)���n�R��@�F�4u��&@�	�o����q�,�����}�.K��٣y�@��\d6Ms��*��b�З��?KיD�_t]*��������ML�O��A/�܃��8��$%m�}�Z��c�U�ǔB�I�qC�~���M�?==� �F�J���Wt�Xy��.�3
����E�$/��҂ک9��K���u��LF�#s��t<�^���z�9�����~�i�Έk���� +\{rA���$����@-��h�ª��4O�e�PR
Q��%
�a���S�[r�©�5��"΁�S�A��5���l���J��WP�Jl�w�"Z��q� �mqj��V+b�l�"b��;F�]�F�]Z�|^9��^��'|]W~r��������<,](��B��r���s���̃���-"����-�7������+��<�+��/W8�롿*SR��x��Cq�\�_���+6�j�&U�H����#����؃��?������./���cDxM��\@r��:�����,Z&%/~�
����pg�b�^����@�^���Ƹ�k�A�B�Y#[�i������IU@PE�'C� N�i�\1ZU�%ƹ�|w�`���]$�'}m�R<a�*������~_j6y OȨ2퍞+m�@<4��Ê�c-�,�� @�}�Lg��iV��m��Ŕ���]u��͵��Z�]}�+�DͨC�Xa;5�|�4t�,�fК\
����+cm\ %�	�!�J�Gg�������p���:zi�~�ONy����5�n��&i���;ݬ�����f�NW��?�]�z�`:�����!FH�DFF6�
l��M8�,�X!�'*����zq�E�BNV����t˄6��+G=��� g�ů��P�r+�mF��*��6�������WI�gS`�m=+9��>�sF���	�")0�y�|(���r �P9�29c�)QgC`"�J�˻��tXTl�r��d�¸n+�e�B�9��o��ּ������Dk��Rc7��q����g=�W�eX�*��_���?����+����2X�4BtK�a*����0��jy��|mY��Y����2�VQ�Z;X@����&Ͻ���HR�jZ\X�a�p5H ��CJ9�%^�h,f#P�y�VK�G�mm�C{��c"�1</`�1ZH7��V)v�6Uv��HrI�>_�}�KD<dm�k��S��:���������a����y~x%�оQM��Fh誢���C[[�JX�an��cn��a�V�� τ�sVJR�J���N�H��8�6�U[`�X���鏇���Ϸ�0�+�}�ZX�R��t�[@�8̶N�	��5�:���l��`�M|�sn�lh��D��
��0T8��xUP٬l�������t��O�dׯ�3��К�5��;���Xp�9��@k� �!�w'���+��"�Y+�Y���'9Hu�Y˷dv�q�w����u}��mr��_8J>L(���L�"�K���������t_=��KQ����jt�7��a��̬������+����ZF���Eh�V�aDQ�e�����7^}�Gxd�����g�0�A��I-QO�>�iS�3�4�Ghwvw� �.�D��VzX'?�G��n0Ie�b�'�2*�^^ ��nvQ�3ش��.,��c!h/u�w!u�^�K��~0V|jnnn��#n��S(ɴA����T��m���5��(�	KIM��`��_�9�^�;ݑr~E����]�F�����-����น�L)޳Q�e�os���u7  I(d<�+\���)orS5�y���W�§��!��T�P{�ߒ���th����h�������t[yl��!�rԊ0-[�fk�f�.[	���o�/�9�ţ��]�t��4rn������`\�C��ds��YV��-3e����ceآjv	ŵ�3�:0����x��i�#�'�],.;c�FVy�1G��+!�V_�.��ן�G���\R�d_
u_A��H^Jt?|�$e��������{%%��f����uuu���^2B�^Ԅ�xׯ_�mY����#ǃ?!��[J��DQ0v�Pғ45=��EQ��1��7��Ѕ>R��
�5�����X�,Z�������/ٛ���:&̣;$	Y4�[���W>��?�g��"Z�ėvg��i{{��'_�SÖ`�:��J .3��AZ¾z-�W�����v�[�c����@�{|�W�D(�-�f �S����f?U'�������Ը@��8=����� �Z)ua!�� 4{��2Y��]n�fp�q8lw��M�{�ȕ(������:�ހxD ��?�_��2�y��6��@l���6��l��qm�/ނz�HA���=���WW��M�&�E��7ۜ�-j�(r|�\�Ҁ������>����1 ��J]ⴍZ�]��k�%�XJ�%�,�vD��_����:l����"4��M���w�M�s�Y�u!hǁU/�Y���dǳ�B�ONX��}A�w�	�r����@�[��Y�&����,�Լ�n��VEl��%�3ü��φwcإ�S�E�M��Ϟ��{�;>::�/��lBB�"���*#;'�U�^�}~��$-��%��x����D
�"�]��X���Jy���=�v�5E蝘��	���o�~�	cRi|����Q�����Z�+����нg��D�M1�2�\��IB�-���{�H�M4��8p���;
x����7�0�8N:L�����6�u��tÓ/�w������'>�t��<ώ���x�A*C uP�vp��%�$�^;�t�.��:7v�������j�/��o�s����h#4́y3#�����M��Bn��A����0\I�.q��y ��ҞPИ�Vq�_��ԏ�i�����C*!oi���f�w�N��3)*)��3\��a5i�R����5�0��y����&~ߪ�u:�˭��\�cǞÁ�m����{?&���(�+w����P��QJ���w�㙑=�-��q�#��m`��+�W?��[9ڥ�%��-��{�k�Ў��km�+�fN��w	�A$	�P���i���g\�hXu!��D��p�DMk-jՄF���
[+��&�#?�,�Ց���7�2��vU=����]�h%�%�fѻ}9�;�rލ�/�oϻ��Bzc��]mq|v�]�_LG�>7�W��ٿh��'��J�n���ݔ�QA�;I|V�xF��(�F�чnn�|��&�;q�!yࣜ`�� BzRY鵠�|V�S�8�˦� �L�!�ӓa�#�efo���0ȸ��P[�i�"�Q�=���J�I·G�J���HW��p���r.l����������N���v!V��<��ܶO��2ao�ߟY��Z��T��I3��^9�dOf�r�n�����,p��,𱺱y���/�8��`':u��ղ畇���_�Q���Ż��fX:F=��2����B�.��5� 1�9�͖���҈	&&��!���q&ЃYC�LOߞ������t+j�U!h볺����O? ���4KrP�Dѥ댺z|8�R����I���55�+/?R��d;�^˚I�C��bz��:3��EP;�5���wЊ;�����mݔKk�'�S��ZB��
���0�Eָ�=U�� L ����߹�t��M�_�V�9b�H��_�0��JIs�W�u@�G���s���477��x8��{�EBB��5�I�Tf/�pm�,�w���pY�D���='��p5��F�o�;R$�J�GR�89�8�?u�5IZay> ����R3x�n����L�$��t�"ԳE�-sM��4�z@��'�A��_�k�BO�'տl齄�I��0ɉ*���X.$�쯽ظ�
ь�҈������ϧ��]>�;�ݻw�ǔ�4(3�h����$�,�QI�WW�b7,@a:4�l~;��Y{\�m�|�Vh��l	c;N=�-G�g���m������׍C�� �\�!���@�l]�gZ�MA.��mNNN?3��B8!�I�)�pf�K+�6�Lx�(G���ֵF�JG/��	R�H���~��4��-0�AA`���޷u��^�yr4��ӻ.�o���q!�LD[�`�=;G�B\�_ߤ2�)=��&�e�CW��qD��A�Rf�,����֍�d���i�$Mά�H�=~tbbb�c�ne0�EZ"%b�d(TM�v�wL�[{�zFi7ݲN�����Q� �ۇ������|F���� @��ʽ�O���V;Bk��ٹZ��ː��F�����j/����-1�d��|�%�gڣ�i�+^�3�J2o�^��I8��ne�8���L�J����e��B�91Z���F�������"~�k!xzjbw$3�!LڇV�qڍ�N+s��z�R`�c{�\v_�	.���q/
��X��d����f���#��^)���SB�����b�U��S� ���d(4������2xY &��~��8�c���Y�������1�E�K#(�p=+�U��������--j����j222M[,��ބVƫ��3E�2*j	�"̔Pe�
�p�ǩ8>A�@{�K	t��Q��QZ>+e�������Ql��#UϚ�� �}��s���>���uTB��˨(z�ɔ���v?y��A�����wĝ�|9@~�3I� ��+1v�>>S��I�x%��9p:�F��.�Ԩc:��P����҈1��W$4��K�qV��9���#/�ϼm>�(��6 �;�H���o��'_m�e����sF����F/=�E���w��/U���d�%�KV�w�p1@�T�I���d9�_����x�J�l_vߡ�]�b���D��*�S�����g�>�h'��l�}�u&e�7�����h�+7.���Es�{F�#>�E\!�DRV��3_/�D��%���n��ˠ5I���qɚ�R��t���~L�%p&3㾮~��HS4����r���V3ǝ[�<~��bԐ�~�8HV �;WiS���P��C�® T�#���!/6p|�Yf��UzkСV��6���l,Z��§ٺB~B>��Dˣ��%�5Cv�2#���Ҡ't�0���&�	�Ԁ�
���N�p�j����9?c��j�ٵ>$��)q3��"�S��Q�3���sK�K@�g�9�{##���9ù���k} ��-��� �Xq\.���p9��P{�����L�^ɌVњ���f,�]��<�]+�)T�z;��ڑvc�9�KݑO�B��%�m��\Ȟra�p�÷�	m"��{�����/���{O����M���.-��(�{��t_�{���K���#D�Bw>L�!V0 5�r����k:�����|�e@=�vww��������!h���iD���� <�Ah	uu�Z��Y�߯��{�|��`���j���&�clNh��?����L���Z��=v�y�'�B1w�IP�k�W:����ơ���`3��[0���+�~o���`���j�)� ��UϞ�oll���OB��Uk���o!�	uJ�>\?ߖ�w�GQeJ�	U�K���K��1ߐع������2F\�C��M�Al"��>�z����y��lv�ÿ��٤�0�r���p�G�������V�ӋTpn\��ii���'�4z斟��#��� [g�=�jp��49:�� S$��F��l<�~��nR2����n���1�N(�`1�Tkjax}3AGI��`����%�����y'bc��^?�(���Ȕ��/X�WBCb�9wy���s�%����9$��QV��f@&<���t%[�q=�b��q-�,�d&=���e�񝅘ZN����E���{���6
]_��Ʉw?}�tlfjJyqiI�%�h������
0V
�݄�]a�8�)^7���iу�zh�����$ÏI�Y>����ץ���9w�[w]��S�>�M*3xЛ˸|k��մ���ʉ��"{l��7_��_�x�#hM��p�w�plJ���X�yZ:���n���W9@��JE.��A�US[e�Gׄu�'�"�H�Nm�J�쪯���d�#r}}x�N��R�祖�o��Z�.��V���$0�J��_��Λ����X&��:?Ս-�����?y�a��y��!*H6�E8]O9;�3��Ֆ���]o�=�d"�`^�9�c;�7��@�6�L�ߘ��o\��A��a�c�Ԫu�\@�u��w4:����K>0Iwc����7i����n뀶����F��7� Y�ƪD��\�^� ��IN%�m�fE0=�y���t��P��szKz?z�R�g~gA&�z�����>	�9��i&�&��aco�Q���<�����T�L�k��	����� E��z�a"��2\�4U��p��$��p��:�O=�ᆪ��l/��R�̴�d�YRqE�Si`h��]�'�`Q%qAG5*pG��B�yΰfq��^><�.��C��K�K!Z�i}��м���	q��t��a�3&/da�h�{���n=Q<a��`]J�_U��k��
���CA�H����st8µ棖�73�.��<J�/��X���=]��D���le3���}�d�>��^*�ف��i�Bb�_�ٙ	C�l� ��eJ�W�(��mn����`pW�6}���ОX�Kzs�j��\�C
�\���J�X���ڝ|�h�Z\�U����]y9�(J'��p6�P��FK��s	�향���0��N���r��ba�2�N�>/�Wkd�9�� M-���a�N1_��&i{jζn8��m����E�op3f�v��禦��ʿr�HH�������|odV� V�fk384�[P�Bd��v�m~⦜��n8p����#�ZLP��K��U�&{�@ǣL�W1�f9]D�fE��w�X�an�������A�%"�I�|uk2߫S���Ȼ�λ����P�p����E��Y�q�r��JK��x&��vk��Cp��KP�J��*׾3���t���j-��8
pG������[-���V�p������8^�|aWKDx7��Ol�z�C��Fe���+�X##f�^��������8S��mɏ�@=~F#���I7,���#�
����b���n�>h=m���2��ֈ�l~]aD�Ƕ��3J��ȂT�K"a.�Lp"\VJ��"�ڙεQԣڅrz+z�,Ì��zF]v�SwF�n���r�{)���yj��a�(�e��0���;v�5�|�1A��<��(��s�Kj�#��?�����{���I���)\A-/��t���7��O"G)^�߬l1�Ѫ�PCI�F����������Lx%����D(D�gA�(�!�蒸y.ӧ]H,5����@�h�Eh��Nk�Y�^&�E[B��{���CU����3��b��0V�	'�/�3�	�c���G�4/űՎf�	 :k�����:������z+��e���0������R�� ����ԍC��A�Av��!�Fwd��o�w΁Pv��$�6�6R��K��Q��A
�z����yjR� ����9��[��!=�'��C������	wي�#;8�<��sF�Ŋ+-��p�S�)t�aN�;��{�fG1AQ�*�D�K`&���7{�����]L���/a��@�Z�* ��4��C��Q磛����Ӱ:1:Y'e�Z��V����ƫ=�C�n*�ƚ7�w�~��힗R\3Ҍ�th�b�y ��^����������k �3�yn��129Y�vDi��)�}ϣד�F����J��1z 5������bӔF���2����)�I�ѶD�?�wm	I�f�m����A��㳋!@j�f/GN�{��dlP�;��<�l(�K}Jd��O�R*�[;3�VU�p-�-u�	fGʲ/ޅen�!�3x�o��|#�e�`ל��3�������:��g�N���/��>b^9xۤ��ܵ��>�W=:{�i8��r�G��E�� [[��ǰR�[����/��e�-���Ke"�k�z�;C.{d�v3��%c�=��J����RJ�B��#Tg�D�����rе,uY t8���,��!nʡ���4�Ƚ[�D�4H&RDVX�L~Y�=��av߾�E�@�mJ�"���\�G��9O:P/�
�,o�.�W�=*� �
�ä�����ǍaX����߬\a�K�~���� ��]��`����kU}V�x������	�.}u�T1=*6,�](�l9:�����@��xR� ���&��>;�~N*טe���8���@�1�H������8w,��MJm��#v:Y{\�K��� E^��w*��lW��C���k!vj�3�E-�1"���F��N�ׇW�f1���y��t���`G�g*�V6�����;U?���*} �������H"Hf��:�V��b�B��NΣ��Gz&[��8?v��;��EH����&��n�6��1��ԃ��c����еҤ�M��x
(��N��)t}7*��a��)���s"q�Y�,�+Q��</59J�"���a�/Y��ʥ�-�bF��3�eU��u�e��W�3���v�����F���y��/3&F�1�.;� u&��i��X����] ����!?�N�s�j|��	�w!�p�m��M�3�c�t��A��{Hބ�<,8�&���/7�5)�mZA����Te0z��3��xw�٧.��v�cj3Vb�Fb��n:��)=jnc��+�Pj�������]S��4Ҩ'�.Ru�;	5{�k�֦��Z�#�0�����#x��Q�O�(�?<��w��߼4��K(1.S���������k�%�jH��a-]D5���S��O �w�-����w�\�@�̯�9�W>��Y"`	�8����0�(����ɦ���a�	玦��C5kph�e�K|)����9@�XH�=`��[�c��=����Ws�,��K���z�G��C�H�`�La�+=�Khw�����>;����Ʒ�P���+	:TCN���i�ͱ�쳎5	۵��gfL
���7 �L�k�3%�Ŵ�9��Uf�1�5R[q$���P�m_�m�|�1�N��"��n��w<��/�}xxy�d1Y����O��`x�g̒8��6K\�'k��۩��0fJ<��w�o+-;����] ��}��o�����ށU��q�˝ʮ�:	�����.�����;��MQ\�������7q��b^o��}Gamn��@������r�X$Y���K��^������f��;�My6^G�Rh����0 ]:
�ĮL���Y�Q��v.�T�L��.�$C�>
qy��O��U�v
}�8^O�gH��ed/��	�h*�7R�L�G�;�X[�B�-��wR�l0M��	y���nu�Xo	9��-�lၚ��JS��х�GFvF2-�t ^0h�^��GC�U�L�m��xr �wl_��{�&="BOe� 2Ę)9�6�R|���H�ͺe���ڍ��'���BY����q�#�py�R�0�P�n�f��B��<v}Aǜ�!�,���u0t��H���f��ȱ��a�MY�l �E^����jx�l��:�RE�48��>��n��q~{�R����o����O������3�IPQ�����X�8�J��=t��0��� �:��u�2���J��a2��2�/"�3�,'��Кx�_��qj�e��ޥ�#��Q�y�B}��{U�}�]@h��C�6��ǎ����z.����O(�۔.f���'8B.�i��{I/q��o�{�~���c�C���x�f�Ceqv�b��՝<)����Q8�	�q�]xHf�"��ސW��V ��.y;�p�#;z��K)>�e���/�{C��Oo'�3��H�s8	��bڵ��&�X��u�4�o4A���>�pW�-{X��m���<�)�`
^3��'�G�S*sHy,C��HG�_�(�:�sa������pܺ�z�VylS�*gB�d�a}������2Ό ��&/�H�٧P���׉4K�g�͔>!�"N8 �s�p,�����;nhܙ�LƔY[ ,�Lח�uI���kG#f���531=�fC!棓���و1}����$Dx� ��������vh����넌x�7��ۖ��	����_<{�os�~���������E�q�D�E��DR���B�k0����e��E�5�� Ǝ�N}܋�_$���B>,|�@"����h�l�'�� pV%�{���W�"���K��9�I���H@�*�/��%��IG����H`���?���k�d~����D����}�*M���PK   ]��X� ��! �3 /   images/ff7168f4-0295-414d-88fb-5470e87041c4.pngd{eP\A��������݃���u��%�BBܝ �%�Kp�`����߭�����vg��������5�1���@ ����.��!��B�	���TwC/(���.��^�%�����7[o?O����������������	2��� ���a�A1��T=o!�Ŗٖ���A���GT噧cԅr�k��,����vH58Q�ͤq�������Å3x�HI^c�P�~Q{��gxei{�v�Jv�"�����pI��í�m��͔	��8�g� ��v)�Ep+uc�aʪ�b	D���� O��8x��A������#�֟���OQ<#�����F�[�<Q�kU_,j	����},��php��E�l�z���:^)�����z�o�FR"��:���y���B�	��.���'�җ9����l�휗9d	>��z�w�/s��#�Ү?��@��C�]��s9�����D�z>�RF!�Xj��h�G��rѩg[xq�h��2�i�����$id&�`EQ��R,楚�Pĩ�W^ }��ƽ܅c��??���`.q���d���/*�
�9S���L�(���{���8��j��ѹ���b��Mҥ�����U��#I���ջlA���G�,��ϐH)l��̑�������Ļ����Ĳ!��jV�H��`bG�ϻ�2.q�",̮����H���r��1#��OVp5�-A�[��%��q���H��]���<9�6��&EB�(R���n"0��_�մ�9Z	b�@���&�ghk����������.n��x�}Z�V����!���UT8���<<
]�`����s�ǔ���{��x:_�7�K�!���B��Q:9ځ�)��+Gг����蒖t��d�E+�^4j-���?�|b઺=hzQ�w��)!�nա�9��
�-�W�_kVg��Qe��7et�R����edע�g���T��{T�q�O/dՐ>�o����5c�,�����}xW�$x�)o��_���ƈ�8�2�z�#��7~hP��4�h��}�/���'z������و��ޟ^r���}pCY�E��~� �p�J���Q��[�y�f��� q�+FO)#�$���9)�Y�����������o�*�*�����]�{�3���Ji�<�e�y:ɣ{��U4�bf��߮	͛ͮ��e�i�<�#����~g��Ro(�8�EA�{�`��A�������ټ6JńY�-+��+��ȤX��o֚˙���6�J��}�	�`B>B:�_uI*	�����VB_@�q��������r�����l�����7�t�<�D�ë�uD�Hw��jjǢCS����t�H[`}KL�O�38����݇���R@AzE�h�"��n�T��Iy�.���.���^y
?ܲ��f�;�i�3SU�N�Ä��	��{J��� �z�@�������[s}{]�,�i+E`ЙV�:�y����ïH��wy{)N�o;���^<l�~Ic�
�������w�Z=%�^�X	�ů���NWD
�j�d<�N-ۮl�
{E��������|����=���?}�"�$� ��#���(�vG"����
��P��?D�zr ��j���`�����l��0e�z}�~X��q��S�i�Qʸ���A��a%�;>�l�5EG`���ul$��̍#�EOC5�G�>}�Br�0��8�"=L�o�]x'�^���wxz��~�S���.��NA�d���Z�p�~4��Y-Ƕ��=�L��q�̸WO�s�*{���Qf�)%��H�¤��:���� �K25��eË�%y��@q���	K�"�ŗ�c�/���4���oxY�[�	ت���"}?>�eF2��(*8�@&	|���%/��b��$�m�
@V"�83�`Q�������c��D��Fx^,g�WeN�R^M6Ŷl �j&O�DE�^���� ʍ�G����s��Ʋq��r��xVa�*x=�^�pEt}��҂���k�$/�� �K+��v?I��$iߞU�M���2�;�;q�1��b$��a�,��[څ�f[c�Q��Ř�(�c�����ڲw!&/c�3�������Tm�㉗����nW��7����-��r瓚'!�`B���
���>Pb�a!�������M���p���u/pz��Ӵ�s�'L&2�&�R�MY?� ���B�֞>/̂+�]�����`�R<va�LZȟi�*i=���)z����ē1|Y�D�"�QA =�3�`�2�b-�����r�/Y-	G��tk+h����^&Z�b3�I��/�M�@}uf/�ሺ��:�b�Y��x����ǳ��զۭ�^`��<II�L<�ۖ@��z>wD�:I$1((��{������}7�.6鯿��XdYX��J�;���h����0�1LO�78
�����������5u	T-���?�œ���Z����Ya:r%��<��W�S���i��e�0�s9�hi��I�)���OU��t�u���6x���zA���}��l����d	�1��ˀ��7��^����S?�ʺk��O�bG�����3{����⬰�pQ��Z��'�7�s����J���=������m����$�Nrca��Bn����٦4�cЅ�(�nTTACz�� bg�ϠU)�n�2�g�kƹ$��_�ߠM͞��T�u��R}>!�s�U:��9�����y�QQtLEc�wT+,����W��s�7��4v%:#JmiD�ٕr�2��S˲$�U���E����5�C�e+2���B�&��P�?8q�ʘk�`�0m&9����9Ë�Zﬀe'P{Џ>�N~y�aܑ�,���h�>��cY��E-�D�x�'�Нv�O	�T�u-Q ��$�(Q�4-ZI��ړKI�J�ײ��Jr���.j�Z�L�#~%�J�s��&fEyq��yjB��?rO}�i2��������Fz��_o��(ŠId2;�P����q��@�Z2&�ؓj�F�^	s-��u���^ �xG.?��d�5���W��+�|��-�^�%{92'��z���K]V��O{ou1�N� *�,
�0~Ca�(%�?��-fx��*�b�= ��i�<M��Kc�z�J��b�'���Mw�d�3�*@�&G�_��*jW\�:�W�z�"��hF&�--�^�6:p�S������ͫ�N։��KL����L���e�R���2�� �GǸKǵ�^�^ u�H���EJ�#�����V*�	�g�m�����9���"\-���%��d�/���#�F#ˋ[6����t秫�wf�ӮTF�ߟ���+�G����H�`�mW�9�X+:�K�25풮���_���8�a�
&�G0�Ac��.hP5�_X�Y���b��]��0�޳	�K�#a�54K'�
 ǂj-F�}�z�
�totIo�/y����b��5��!�h��T��D�������N�݌�r����ԛYOʸRnIJ�ym�-���g�:�n�I��.WU6E���;m������6����T=Wb1igG�ԍ�~�h�8���}�����D+	�#���Z3	�w͒��U�^Hc ?�jn��p ��|#������% d7$�Ю*ǝ��4\)V?TP��PbW�mN<���'ؑH�ZbջH��,�i�����!�����]���� �c�3*��Z���tG���pؐ33dS��Tу���1��s~�>fd���+�	����_�ӓc��?�.���b��УA��;+�����I���J<��am'La�l��������;���dͶ�!u���
x�]��=sSq�UVi�Qb_�M3��Fv��t�6�J�Fv-���fki�B�('�Y�FJà��s�kiW���P[�p?4		�Y9��.������֙x>>V1�0`���TNLSd��y�0����!��#�v0��E��%<TK��,C��z$�6�}�����V��A
W���y��P���������W�G�2'r������Я!�Xǎb���o�Wﻈ��1FZWi�\�Q��_Κ��JFQ�{�׻�:Q�܋�>�?ny�"*�U��#��?��r�FJ7Q�D6z��5���()��E*��708�J�}?	�`:�O�4�4}��1�� �F����]�@�Lͣ�L��ۊh�����|��F�4��ݥ�����O-����-��誰��!��vOr;͇���1�0�o� -:�l��\d!���+'֗O)���wͰ$�L�S��Z�,��/`���@��{�@@bA���9]��q� ����Bˁ�7UeݭQ�YG���s��=�J������GN�w.�E%/���v��/����hʡ[�"Ek՞����Nt�`�
D�������H!�GO����S�	;�UP��t8b� cL�A�=MG���' ��T��-KH��KG���:)e3Y����������Xw��mĆ�����x~�����<���l����M�}��\�`�i+��M�gzu�]�ՀA<��Ԣ���O��4L��⏢����cɋ��7�$_%���W�
��n~Jh�/:H����|�')7?���'@�|JR侄)L;����R隭�����0�/��n���W�E�ܢ��&�E���{�Oo��|d��MM��'����\���c�H�#�c���?<�2�Ua(���}^��"����>֫�����U�k�nK��l&�K�ۏ�F�2�fc��$Ǿi@}�c܇��.��)��I᥃��И�a�s�-������ƿ0���9��ó��_7e �rſ���!����U� Ds0E��X)e��i���-�8�b��O�؅~�1"Be%ݼlD�\^��|�4��E#���є��uV��"f�_da>���3�!�8������|D��_;l�"Ҟ|�>{z��m����I���i#�(Mx=�5��рA�Dq��?����7�y~.��C�����!�j�q=]O~��^�}��-�L��eaI ��.����{��sH}aB~"�r(t��=fW��u}�z�{f����t�΀F��r�ZHWtB>s�i��#�b~�L,z3ܶ�|31Y'�x�k�:m͕Niɩ��)�f������O�3��o���I�"T[�J$���~U�oh�B\�Vx���X�����LK�����T���'���V�o]���܂�ECM0-zS�d��EM��c��â��n�U�A���]�J�w�sg�C�}��P$l��:�n������U^Z��P���&���o�-��w�6���W�Y�Z����|�jU<W�|r��:,�B8!vcբ�v�#�		�d�a���)pۢ��񟔡�_1B�&~���e�shF��.�®+��!|B�y������R����/4�L~Ws�fЅY=��3x�/��t������߇@_��kv���{�����@X�˟|���H��1����
w��#��ݼ1f���Đ�dv|i��47%x�������A���a�=�K�E��\���Y�?�m»��A��ju��Y�eD�vE�~���&�1�ްXڏ{�s�tD�y�ῗu�mK-z��廪��ɛ���L���2�fd���Zb=3^J�!����Lzc����#���	C@�B:��η�Z#q6�T\Z����M�f�Z��υ��nd#YX�$�󀾣��V1Moa�<PB.o��^����%T^�ڣ�JVSmC��P4�*��󒿌�^9A��Jbw^�6�滚����]��M������4��A��S�y�)��.�����j�+֌�2M��*L���X��_K�|&;�^V<��,�~cͻ^�}�߇����53��P�ճ�Ɩ�E;�8����Sr�KJX�\����.-g����i�4��Tp�"��@�M��)K��mR��(���I�>��]ރ7��?z�>8T��a�N}~���HU�Jh�WX�a��LV�C�-Q+&w���x\����[��b���=|nu[IFӒ�����g�q|/�n��G�^�	X<|�b��o�w��n�'��8llC�h�����I�� #�Q���`�����Ev�y�̫�=��v~uRBu�-\z�$�zf'!�ی�KP?rZ�J�앯�w���k����yH��'��K��Eќ�G�H����@'��#&�����'�R�.��Lb��(1���)79�aq�!d���`!�m��<��S�ו5�dO-�E��\��P��4:��O~e��^�͏�Z����x�pW�]��p���B	������-�%V�*�z���w�����iiy��{�Q�'�c'*���W`2F~�w�]s��`��? ��8��+���#����~GԷ�L����fm�ݝ�e���C�[��4�_�����0/�Fxu�<j�������Tw�Rf^��i`4f$ ʎ)��px�CNW�)�'����"6� Y�� �P~�,�,����Ik|���I�0]�5 ��҈��t�d�d��m���<�q���C9�k&���;v��K
�Di��	o��Ĕ�;"t�̥��߆��`D6�GB�R��g#?���0-���%M���c����8N�+I���FH�8��M���QGr��1�9���M&4�|��<1\Ƴ��S?};�(T�QRմ��������Kj�<UT��w.9��Ƃ��W]|s���մ�`�ѣ�ܨ��IB�}o9��}+wa ���)A&e"��S�f]^}ɸ�'�i����kw��4��Sek�L\�_1W6t�Bo��_E�X���~'����=���>d��$�C����т��uj?�KOԬw��Q=�I�H�)����4��k�Snc?����0W:)D�Us����.���T���L�Ј��א_�`�x�9U��*��?ކ�n'xe.�H��IbG�bV�Y��bw%2�`ǝ1�F�ڷ�����QKV�
{xd���ț���Z�<���\5�����oY�\RWry���J�UT �5���X�EE�	�ӫ ��C��d�� v�?�k�%T�bu�����ܪ�� ��*E�4��ߑ�]�dIPۥ_N��X�񸓼�n8��6��7�K�j[�G�B�]T�W��N:�}�[�*�1�;����Y3�;��.�Ru뀟�"��~-3:�ug<��g�L�#�I������r�C��"�<�z'��뙼�ET�(g�hP;\�8�q�͵��9 �%!�Y�O�����W�I�0+�"C�v���]�K[KLܽY�h	ie� ejf�He��������[�C��]E�� �99�>#ۍ\���tq��fW�#�������p;�[?蟓XmA;F����awjM��w�A���+t��!���Y���nץnt�!�1�b7U��c��.��<պy6�)��3�giQ
���T���+��k���J�v� ��[���Iǌ���!�N{���zQV��%L��^������@�t����|1��� ~a�}u�)��1nt=��2�#��N���6�9������Q�IDK��\��������Pǭt�η��}��v$�_�[^v�bFKk�Ƹ($���ͧ��e�'�6�x_��9�F�ږ���,/IBI;�lQB�N>@�U�ȟn�i	il�mOL���#u.��[�^����:��$!���^�q�䭭Er@U�P�+fʡ�/��Ao5Y���	2�����p�Y8
c�#ؼ}�h֙�bH&�p��ޢ-���O-Ufs�G���-{�8�M���c}"T�d���} 6V���M��u��H���Y�=13~�����*�Qyu�v.���Կˋ���T����D�����C�ώ��ꂴR���>���c��]7/�e��9��L�g�
Z��1�h$�q���V}1�60f���I�ۃ�=37}����E�vtT�W��Lj[�HY6��f�cG��f��=x$H�La��ub����.���y�FLR�|�N-=��v��_T~?q'��9GnJT�޲}��D$��m�rb������v3149�(w��ܩiyV������Y��P���)��RĮ��*V��[��_7i���8E揷�ڦ��$���(�@{l�"Z�]�#_'9�lO�o�cж�T������gs�)�LH<ұ�����g�����"X�,��Z���E������|��ղK��0�}	�17^�z���mVq�!��?]��W��2�rhT��Ր#�`W6��TX�Ҧ��mZ��ƅ���cn��Վ�<��O���r�|-��,[�,
6Hˠ
�#�|HN�w��W����(>�-H��{��c�%L~(�+��J+��r��96+(�	���hל6ͪp�H�{��{�8��E��B\_(����t�*{n�6�ݫ���
91˵7�Z���E�6����ܦ�?g��՞��j���PY]�~��_@��囬���̒�<M�{D5��{����J���[� �!��7��񛔏�c�ba��}N�)�����j�G鶬�1S�٬L�a�%Ҙ�Ť����\)@����4��������lV؍��m� �E�"9/�K��b�eC��K�qw�t��}$�W����g��{�����;����x_��'kf}�u��e����1�U�篆�k�7�|<�+j</�I)����P>d\�����	����ڧ4Eq�xvW���l�t(�z�:�H��=j����Nf̉��F�F��͇��o�!C��q�" �'�����4�5�[S����w+)�=o�ܔZ;
�9�Y�Q���G3����W��a�PV�	�@%�z- ����&¾�gb���*g�i�'���$#�i����_�J�|�u�;��r;�T��G�q�u!p[���v0���ܴo�%5�8P�L! f�k��z)|���o4c��c?YP
^����M�EHg7�o�07y_���2Ƕ��Lj�w�S��m�0�_�Xk��DǴ+��v�
���m�KO�<S����U�_�o�3i�FP2eO"\絴Ay���0���4�86y��QW3	���J�s�zY�����8*TX�������0=MG����(��(#R�q����a,���(��۞�}�0��6�wC�ߖ��0�F[���(��ٹ����b�'���j�[�y��k>���Q5��mqVE)��:!sC�[�3ʸ�_�4u��K������(�C���`j�V�
�����J�4�������<~�O뾋�cl�v�Xt�N���~Rn?���`�
�RjHV%Mu�+"�2�����d�K�r�eF�)A����nL�5d6��q���m��ʿ`:����N�g@Q�nqF��J��}2,�-p���F�.�t����^�@B�����A3(�������j�6���@��v��#�Ƚ1�T��P�J�q�a�	Rh@�k!��mNR��*�V���Ns#�;5T�K��Fd����b`>]٨(��5��T�*����;���Դ��.�V������:����#����vO�1C�M͗���1�%R_�O"q��;(G�J�5���c�y�1
"�ԑ�K3���]"�F��1��gM�f����E����[^[������xݾ�z]4�n��������enNB�>'!���KԢ3��n�5v��#~�L��aJ��������R���5�[�^��Ư#yJ%փ��[���=[9
��;�i&���赏(��>p��,�]vV(����DV�kC_w]&�!��.p�8��8`��-Q��vũA<⢨Ǻ����o�m����=�?�~f��2o�+Ĳ5�ب>��`*K��~��X���m;�ʷ��n��Ն�6w̩���a���&e(�~��s���KWf��0��ϧ�RK&�2�i!�zڊ�ay�H���\�R5k�Tc���Ц^	",�,�h<�0�7�����}�~/���Z��H&)��5�IY�
��� �hDY�F�E� ��;�m��`1��⌳%�i���o4}x~�Ti�2.�)D/�]�U"��(8 -�}�\5v���i������:�80�,Z����	�+oXJ�Rs'$�;$?BE�i��y\�ZL���ۿ�������sn%9>�^����p���kt�����M��'�₳���T:�~R�Jz`'$ŏ/����S�	�9���=�{*a��+Sd2���S�Bbmc�q�	�/���*����k�x5��%_V�>Ӱ/-�n��#�ɠ�R�W�6�����23�9�l���N�e}x���E�˱\�,��K]����YG!Ʀ��آ
S�xu�H�-Ȫ*�!7�L�����^��
��xS���PEl�Di�
�L$v�N@���592���$%EKEIדi nxC�pϯG�~U0�)�"�me뫪���T�2=F^|������Pl�������)$�^�!68XL���!]���N}\�j����"���0qb��T��K";�?�����E��Q�l��DĲ'�pމ���v�*zH�n�R8k���n.e����%3O�(��]�K$�8���`���@��X�嘯���=v(�44��3�<�q6��?���]�:�M�����#�(�_q��0"�p\����+Q׷h)�"�
Jf�Dr�B���J�Q����x]2U�zUO5��s�
���v�̣6��m��5%>�BA�m�ه0�*�pe��e4-Ҥ���RW�U?�DN�F*:U$󎜠��(�?aj/rG��dۊ���)�Ψ,w'D��;��Kga�i_/K'Vx�A̪R�����9��J8���Cj�]�^����|q|�����N��5�}�&@/�M�"M�>Y���]�Z�
�V�ZU�A��u䔖w$�$sS虳'�/C@�s-�ȣ0p�Ԋ�H�6�q��ǩI 6���QW���"�	r;�}�9�ϰ����(V[�YG�RZ�K|���%~?Ib����@�*M���㊭�3�iz�]"��:V�q\J�����al�t:|>�8��V��A�u��<�$�q����@ۺ�
��9����ީڈ֐��OQ�~&����?!Kۛ�0zg�)�n����`�Oa��
��n�O��}��B�?6c��G�8���1�}@������!�9E�e����|�4
$ݲY��j�D��I��@��K:ڱ��0�5?F�}|�����#�k�a �p��x�;d�z�<Qf�O;J�| Qj�
n�=�kOj��.���[8Yr���(��3��&L��Я�_�_t���T��L>�rR��'���ӫ�몢�4`>Ja/�GuI�A����B�S��!
��!2wK��%�,!q�ag�)e.������׆@�}չ�T�nY�a����7��oUVGl�ӱr>^�T:���O��8=/� �78�{׏P���:�^i�K��u�`޼�*[�*�����t6x��d��\�WQ��0��x4TB�C�P��[*�Ph0�_���o�g�@4NE��*�:!��6�=pVLp;�����i#9�!RB���!�a�lx�g��Hf���J¹�8����L�e�ƨ���i�D�$��gQ��r� b/\�8b�-��)�.�!Yޑb�~�Do����3��?�Qhّ� �' �a�t$l-���-��HB�R��T��*'�p,�^�]��Θt:��-B�rroMd���s�rãx'�~F���`�S�"��͠���)#L�?%�!��E�E��Y@�)�<��m�-:���>E�z���̩�N#���A�ސ\X�-�KBTga#$���V�����f3���Sd64}�v�k
�29�QSҢi��e�:z��B惛���ՔOi��

Csl��9XI\-��̧N���e��1�-�oZ����A�Td���7�+��0zYn�/c���&�48g%M�X����jԄ���=ƱR��d���ypS��zHd���+r��Ƒ�̏��|fƍ}�du�~}c���&q�sZO���G���7
���S#t'�:�ہ<ǡ���-�f����8�!�	x�\H�<��0U$Y[���8�k&��z����գnY��R��n�f�Kjv��wh����b���֏����(��/0[PB�)���%>��i|j��BJ�k�sM͹���v����Nj�s�/��68�b��*ѱ�!L���Bt�}iZ��n���J�W����v�|��㏁���K�"E�M�LT�5**��������]����;<yVC�!�����7�;�@&'�v��s �U�7���9�EI'Vj
+!HUYZ_�$���/��:��`���[�~�MU��U��K���f�e��vO�!S��/�N��6܋s2���X�z�:���͚��3e�':�2)��My�y�<31�� x�N��g>�5�5�v&��_c���0n����4���4?i��L�L@��\���	`O+̙��H����B� !��m2ݱ߈Ǧx]��X�Ô��QA8Xd�d��g��w#���޾(Z�IP'��ܕ�Y��՞cv
�A�yq\���
� �wb��=�L�I��y� ֩��e�� ����
A�3r���"��S��j���
�����W�9%B���^Y�鵏�Sq�HHO�����Zx�Z��C��I���D �͈E_l�S=�=Sx�>cp��|�h�®�D[�=9!K8]Y�F�� I�-M����\u��8�h�wЯ��B�|���ɭ���D�ˉ@ 
�3f�����1(mO@�ĥ�����ئ��@q0����E`1���T���L��qK��`\��/}���^n�` ���i��8BO�9��Ht���m��%^�^ݍ���j,"�	�+�C1�� ��~4���J����D��Rrʋ�{XM8(�f��|W��X<�ߎ�N�J>��R^"d�rn�n��;3��(ʞ�Cy�K2�Z7�I ���#�c�L�g`��#�kݽ}�`o����#�G\)Ξ���"�������'� �j�G���S�_P�#����.q<Z���џ�Z���dȰ9�	��n.�k��w�%�sYn�~�-Xrs��j�M����e��A&�Q��1f�M?�=�J�� p)��9���IV(�b�J/?�mŮ�J�6�iҒY�g^��	�/:z�;{g�74���æ�q��ӼtY��4��hϭaI�1��řD;w����?��a,۷�V�,�ݞ:�;�q4�T/}�X���Q�+`?�QgdoJ ����_�Y��>/স�Ce��iդ�����0��n΍i���ز��m�*�UQ����q('[����|Ӄ�f��L>��]�J,��3I���S��fN4�Q�<M�A��[���V�����L^|��� M~-˩b�6�`�ɾk��R
9VE����a�9�,s:���H29ֶvP���0>���ۮ+�s���;�ͳ��]�Ԋx6�<_Ƥf�
���-��eu֊%������?�A\j۷_��K���D2��W��.�5a��%EII�]���	�u��l����xO�{�|�KM���ۤ��A�>V����h؄Գ��Q�r��uq���`�n����]�g���_G����������<5��ޑ3	�(��o��G���(�uS9� �����v���iY.f�C�Z��z��h�=��4�/!|$Y|�\1�l_�+!��I�lp���]j� U,���E<z��y�P���}c_��Xo��"��R��"Ķ~���,}�J�ː�k�nl��f	7����-E6mN)P������$ F�(L*v�T���w���0g�[/��U�E��h\�y؟R�Ս*w�T��������};+zF��<���JBMޛ|S;5���f򥟈CFnCH�)8؋	\��&X8k� Bk���l�ec5�{�r���{Qek�hf��-!҃t %1,9/�ڈ�{}�6T�!I���JxY�C�����>�����ֱ�sts�遌
�H�c�5���I6�c���G*t�lRՀ����q1�d��*�:���ⱈwG�2�ȯ��D&��Bs��Ӷ� @��E�����\�?�F��w���qNN�R��>��F5ل��<�|8�Ve�fHK�1�:Ǵ�X��"j��y�����B�k��&���_�(�xAE�,��NC�䞫02��|w3�;�Zg"�Ժ��kQ� 8���xA���J��=�O���Ob�zst�2���4<�ӧ�v�VH��3E듫¸���&����=���[S���f��an�-��We"|0�6S��'k��oJ!}E�I�$3w/�Ŵ���t�a�;U�?��Y/c"���4�N��op[��~^�s[�����n�8D�)�mNߍ)�9:X��Y�Q0kC9[MT��f�*���;�joUTQ����W�X���8p��'0�$˫%�d	R_��<��6��c��\)�l�I3gn�(tf��!
��j�jI��(�~��4���]����S�)�"WZak�a�|�����Uv���'������c�(�CKNP�/�[�;��ə�5�@i�Y��'�F�{]�7Y���l��������\I����!�N�L(��̥l!ϫZ�W���;�@K#L����7]k\�2Q��$�y��sZ �ȅ��Ϲೃ�Kk������ҊSk���c*qa�U�j9n��ϖ��=P�u��b~5�[�@+X��|�|ۡm� qx�r�e;�<��������o	�+�:1Ӽ�ӝ��MS`]ڹ|�u��FB��+��)���7�C)�����q�K͵17?��X�I����[����䭣���]L��k+��M�'Hf��"���Yq���Y��/�6q.�����E�*;K�LJ���߸�x�o��u[8���<X�*{��H��J�.����=wq�7Ҫm���h�Q�(`���k�@n��i{5�n\����[�Kfa7lg� �MVU�L�ʺP#ޫ~xz����e:�����)��w�f�Xd�{�֍C�߆6��i9�-I�te�fl��� ���0��G1����A�L��H~�0�V7��޽a��G�s�Z?��Js�	�i:0�&\�{�~s�i���d'���ī�m���?�2�8���K����O,B����q�)K�|�Dv����Vsd�w�"���]�u�26u$iO�,�y*p����n�݈�b/���p�ݛ��µҎ5�Q�d��V4��D���b;�9�E��痤נM|]9@:V�E>��S,>�x�	��&]���C��8�dǑ���|P��`+?@�1��S�Ԑ���`۳�6��/�����wQ�5B�p�-T�q�;â��d����yս؂Ui$�)V(1A}4=����.�,{���t�ƭ����%�Н��g	~�L��	��+�^�9�ןo.p1��@C�*�b$��ς��B;�ՙt��7�G�G�ϭb���/����3����z���@�&��\���"��"/`*Q��Dy�]�艐�·�M-u.c1���ԁY���v��P��0��	�ID�j��SD���	��zy����
JY�!�v�#$��֝;�5�Gb�~V�{�����,�{w�s�].��>M}�e|]I�h�\���i��9{ ����-���!S�g����'}Er@�^��*6௯)� �vO�/��S��S����d,s�bt �&yc�hH&$�h�,��t�=���R�y{���f%�m�fh����=k�z�wH�W�F�@�w�,����/J]0�۩��GP���*,R�Ϗ�G��I�����9�`,��Ѓ��E��Ϥĳy�gn�؏���+³{��T��޹#b?�� K1Ж��.!����|7Ϙ598�[r9�yU�꺁�џ�54�L���݇u�I۱�<	n�6DR$5X=.�>��� �4�Au��懎|��V�+.�s��6t�D��,�p�@��C2�bj�C@��(����`����y Y1���eim_g&&0��w*V鞐�?���_Y��QsZ6��|�T��u��_3�_�K]x�G$�g6�8g��몎ݯ�#�J|�.̯�Ԕ�&������X��cn�'[�G��J�N���J[6���_�$Lo�>1�J�;���[�/�$��ZL5��
�O�,��RP�+�s��y���y���9z�lVr�G)O�T;�B��%BOM"O�n���N6V㈮��d��&�k[b`d�����ǳ�v��B��Y[��5՟Ȑ�ˉR�2�E��U}d��	�8@	i����2��B�N[I���=a���$���S���.�W_������b��jֈsb�]_]����f�s�Ur�dr=����³S�k`D�\~B���Y	����Hǜ	ъ���aL�s���#-褕�k��%H�Խ&%��I���#�K�
U;t��Ŝu��*5�<N��r+D$C=�������y���z?�#dP)Μq�K���J�8��n��ə�N�4�������5�5Ì䉏 8ž���n�o���ܕ�	6R���� ����~|	��C)š:~�����5��Uۭ&QqZ}���8#k�;0�H��������C*�ﲾ�CfQ�vkC����"�gY�����[�E���CI�� "  �4�"��"��(% !�]R���H�8�H=�5���;�}�s}����y��b��^�Y�z���g��'���0��f���:w�tg$�	fV��?8�q^p�/^�f�ym�!����/K�h����-�*���^]�l�q>�Rܲ�����a�I�¡|dKT����������)GQ�'Z�X�
�aY5��Y���QV(}˝�{�5)#�	���k����E������O΅ì,V��F���	[^<�[=͒a��ǜ�x}�O>��̞���}�y+���_i���� xI�8�Of^�=��R�#����ƛ��G�9dD�7`��z�4��8�3P�!�Nxވ��/R�>S����+$�� �.ġo?<�W%	ݘ؝�~|�q~*f������p�Ʊ�Js�M�s�4��W��\�+7B��xc��婙���3J1�����=ϩ<��͍��,�!
M)�'-���}���zu�9�?*�q�x_��D�.�R�A.-7�$��F�]�CU�� ��j�&B�C�ӓ@0J7P�=�+y�M�����I�گ��>5������sx���������;տ\-�"@�k]&�^���!W��Aa]��F*�]O��T�����:�����ٓ�����k��4�}�
�r�r�zT�G��/�d�����WO�i���~��|�<�v�l�?�-����w+�i�]�=^�Y�Ԕ؂`��_��_�<�<���Kq�����>�dm���h�C!�u��/6���gM�Y������`��������}�*G�.�|��~&��u?�MG�R�����J��#x�z��+kF���k(E��<o���_�:��x�智�e��ҋ�����������i�N��g��.�p4|����g�C8y��m��k\��oK���wAB�<�Ql���׻h�3
�����f�3I\�����DLǌc&���:�>7i����	�O>�i��9q�A��Z��m�j��ǴRѶ�$M�>��7�'\�V�4sW�-��!.Fx�.B3g/���~��d��[��!���9�cZE��:RC��8�o?~ӽ�����s��g8��C�[�2�4V'����u�i��.�\)��L7;±!3J�>�jU&��^��=$i��Lw5�_��;����qr��s#u��]�m���"��U����^�_�mb.P����������+Gh�;�%�L���Iy�^Ȉ�v�<�Bh����~����諴\�y���܇��a(*nrc"i+���2N����mځ�	��;���q��^�i5G	ߖ����i�A0����1�������;�>�^^<���G��x�
6kZn6����E�}^����H�P�>r�@f�
;D�gԕ�9�>�dL��#Q�xN���h���W�%e2[�'�>,�g,��
J;�ӘG��?}r�N��0�AR@�Pa"����)�)���/�*ve�P���2w]�>ؙ���]4�M�}y��?�e�W��{���$�9^�8+P58Ny�>��8�j�t������s��JR��I[�����E�w�^��DA�`�v��p��Nwb2��P�����?I��=�ťxwf�}����eTA^�T�7������q���33����x�Y2�� +��-V�aՇ$_p~*5�e���uw4p~~�_v� 3d��B�pPk�%�\��T�<����yL�0�J���]�L,��zDH�ʚN�`�'�G�Jc���IF��3���x2�+�l�`#�~P����U�E�'_OeT��O��A��ʬ@1����A~�'�I�f
!�n!Wt:w�c�|7��3�!�+
�z(sRH��sS�>~Od����x��d�����su����\�/��f,)�ψŉ�H�*��o�u2l����������Ē����u�x�9xe^_Z�W<#�S>�{�G�7`�_f3��ə1�+_��b�]�7������~��L����`�9��[x��Fő`���ٸ�I"W�p!�gx�Q��=�Bd�~�퍻����|�t�,��G��fV:+��*}�U�=?�!�<�	l՛����BaQ���H�Wrи�bd�<e��ٰ�>d�Pr�q���}JdΣ�w���D��C�q������z�~������.?�x�<U��[�W3|6W�RCX>+8�I�ֳ���b��Bw�^�$�Ѯ�t���7yQ����������*��1�5x72
����v��w��;SN3����}R�*]�Е�ӳ���+z2g����E������׫(�`�kg���+�"���0u��%ٺ�u[Qˡ��ʳ0*���j���_�A��'�|_�~�1x�Z����R���U��|`��>u�Z8J2�񙸛U�/��^��ޝw�<kmN{�!����òؑ�<X/.�����,'+�B�P6�佺ƈ�������sm�@~5LL�ި���/>�5�	����a�Z�Ltlg����"����k�5*�R!�����*oK)a��(��ߨ8��F�����7{;ڽ��s��I��m�֚�XݹO�uwv���~N(hμ>k��+5d�[�͋��,˫�����!Z�f�RK�����H��J�ӣqVvȗ|��ɦ���Y
���1��yʭ����hH_�>V[�<P7���a1��a�����.wIN�����'e�T�N1"�<�&�Gz�Zc�=��6��Rm�N~��,-}t�M�ҙSt|].�5������=�I�7�!��:;;nWD6b��n��gh�c��3����3�W��lCms{!r7�Y)Ũ��mZ��n�d:�������a���Y��>��풹�ϪvQ~zaG��^�!qe�[���O�uy?�2�� �?�8tx�E�+��xK� ;)q޻��GhgX�ͫ���0��~��f>�WT���s��	z/,���[�߳}�v]���X�̟�0p�ZW񁏦Mχ�Q��}�n�B���|��K�f@|��L^.�zά��Ҭs���*������yO����02��%�$R&F���
}*���F�q��2���lr/.T�;y ���:�Q͗�϶|��R��xRn?749_��+;�Rϒ��A=��1w���.����)4،���8��fC��r.�uи��$JX-"��oKY�mn���{�=��A�qͅn��"ԙ��l��*i��:��D�4������Q�5ߍi������n���h[�@��O��Δ}wĖm�`_m��f����V`h�������C�����w8�n|̽J���.6-����y?L�8�m�?3e�9g�H>u��|�H���R�~�{���4��18p��dC����V(,��-32�xZ���p����o�2���IB�I���庂�+�:�4�OPO�
�Ŕ&�>pV���*�L�FyZ-g�Vg���F4�"uTD��觳���ԥ^i��M1��<�d�,u$o�g����Gh�_ ��7ܭ���Y��8�0Ezܾ8o��)���b�W��}�k�j{�L����H��ݨ�{�Q�kˇąuII���
���[���Wδ�5B���G)V
���O�fs� �2��[���m�@<����u�DK.Y�����&j�s��=��d(.�/�yA��.��V�X�Ϙ����+j��]vv~UȜϫ�0�D�{����p�������
*�=,F
�'p�X�I7�9�A��^�R�P��y�f��vך��Tp�u:�Ή'=]s	�T�Uߢך~]1�F��5�Ԛ�tC��l��/�߄�+FL��~Մ&�3�3�IM�y�*��V<�[J�$Pa�Í2MW��j�����Q®=��R�	��1��_Y&";T*ag���Ψ�4����㠒�eq��?E�V
憝&�%�x���Jx�,��"gv>��-�=>��[M�zHw(�V�\8��q�ҽp� �i2�����.U��<i�%7� �y����=GM��3�.��MA6�F���H1u�b�z��W��a��r�FT��9s�w��z�X9�A��������j`f��M�؈��
SuY���l��!�܆V��wLl�2ڙ�c6ɓ�9�̹�6@��*�L���Βk�z�=��:���n\��a�<٭:*]�<�G�[0�*����S�R'�:�^�����2��㊾�����l5�/��N�y�X�.�0�v��x��=���V֣��zkL��=��ъ:�W����D�&�S,��4Do��Fz��n�r�	�ӡ^�ae�63��qyH+�~�$!��9��j2&|��-%�x�So��J���v��,���*��s�� ��T��w�)>Յ�9��#:��a�fS�j���:�S����7ɎH�ڡun{�����R��`��7<��d�R^u�����9����~��P��\NY���M<,��l �%4�#1�5���L�=��>,�T��+�[݆���<�{(&�^.=�+1����s�ݨ�*)���;ߚ��T���q�R��!c�rI���I�<ϟo߈-
��,��	��"v��j
!u���!��n&��<��/�W��>�څ�PK(yY?�p�v98K��s:��Tc0vI� �(�0�ô���o�P������m�+����/5�Ա�>c�^���������&������\o���d�|kQ^d.Z�X����}�u!�2�؀�,��܉�Z ��V��=�/R|��F��hc��R��d��Ѭ��Ng�!�Jj3��[�%vp�Q7\�A1��9�������W�K����f�uF%e�.*�$�����I�\*)Yeٔh.7K���(dGM�ΜK��)�\K;�â�0��ץ�e\��Y�xK�]���;�e���q����%�x4Vm F��n����/��$T�w/��1����r� ��"*��i�\*���#3��)�^8�J�F������G�_�l�:%��hE� ��&R
ȥ��~Z�P���f�Y��S�%גU*#ZW�9]T*�5m
c�����2����˖�Gvg�y+adL�e׏��T��2"��g�$J�~���1<�q���A1]Dep�j��"L�J����}�t&6�Z�<�}���H��.��~�n���#�;�eP�����+�u��#p�&����3�_���r�}�M1E���6"����c����Dy���YX��2�G�W����R�(/�?���0��j��Fwp��.�����n�������ƈ]�('��8޶%�h,��$�>�a1�c���E�_�-H�/T�,��Z�Zp7�.��nPW�BZȐ}��Sp��]g�h���1f�lCm���ѯ�<����Z���!��3JGz�Z.g�D6IX��o/��/��kf.���^�q�C���g�E�%u�g��);eNx�>�E�̠�������[��$8����!fĪ�l�u�zDt���VMqbYX(Z���Ä ?�%�r��}��CT
��Ɣ_Pv-O���|�i;5��პ��:ūJ������r_o��-;���.�؏�h_��xI�c ��ٚ�;_[�<��b��ݲ�"VyCz��5ake|~����p0{�O;��&�(/�g8��'����O����U麐�r�V^e71����w�jI6��Z������}U9���i�7�t�=���H��`�l�\�}ww�Z�I�'`�x�o'�٨�.q��#�;�q��#ŶO1�h�~yd�*m��Q?�6�5�i��u�:k���q��S�ѿt0'��A��i50_��J4�T�LݹshuWMpn����F�(�?����0����GC=sઃw�a����@�h{���k	/�tE��[V�P��Q����0��\e{����t^�e�Ѧ�p�R�\z\vo��� 1@p�n$���x\����e�˻��l Ā����A�i��D2J��]��#�} ��+ϥ�Vv��h-YSTI�h]���e;;����ߤ���.�9�ת����T��H����@�(�A���,= ������>�`:�5�9'/��J����y�sg�0w�586�g0�@�u3�'�t�����DO���Hk��kw7�� ���?YG���(�ue�P�Î5ߨS/��Q�1��e���]�-���%��`���j��Mc�f�s������.��*Z#��9�����֑ ��xvz]�i���)��[������h�S�+x�w���&}[�T��0�!дylurH)��"6/��A�U0��/�W���[�)�,��H {o�e���q� h'���1$AV����V	O��C�H� ��Σ����]@9V��g}�Y��x{鱭i�(��I�-���X�x��~�5-,��)�V�"���5�a�ZFj^�}�)Q��e@e�*�5׏�q^k"Rp{^[g���x� 3�ο&�������M�o�*��:��p��^�t����\lj�w黍۵����g��z����Gbp����H.Յ�l֥�K�4*g����yuQ%Q;H�y{�FA�K�T)��.�7�k�g�|[<�/+���;\	5�)"i��.Ԣ��L�p23��|�ǃ��콸S�����ގ�Rj�e����\ʦ���>��
S�|�&t-�^��aIbY�+_���	6fh��u�h�ˈi��~�\�E�5�V�.g(��)�������GcaO�^a�g��1�t�����F%��κCP�\O�?{��&o3Z(�w���e*�H��Au"�c�<�T<Z���%w+�3�?���MJ�6%��]���\�x�����i]-9�{�{z/�w-��S��؈p/�dM��/�h����uV���e�����@�[R����.��2m_V�������.=
B�oe�'�p�������(<��u����o��	�Lq�f}s�p�Cr�}`�f_�,V�$\�|��@����f6N�.�s�d�=�u��֠����s�N��ĵ1��Z���p��ý�6�X������TEu8��?�;X� ������U�7^����luU�B<@�lS��l�@p�k�/8�6S>�ٲˬ��u�{�{a�n{_�ڢ>��Z!v>ؓOqݾ^��K;>&�#z�	�J`~Ȣ�pVf�/�}f��f��$
����(�/47N}���,��=�nR[7}� P-�u|v~�����1Si�Y���=R�����͌3�g���5�U���8�����E���g�(��M� 0��+7�i���_^���s���]��᪼-�D!W��3����<*%b�����F#�,�Qp�P�'���eO�8.�����cjs�Km�eώ�/�=���4��ma�qN���Tkv�X�x?^ڟ�fe�(�!����*��FvrgCIġ�%�u����%�((���5V&_m��)�4+�SArx�����L�\��N�ѷ�d斍�b���y��<�[O��a�yU-�+COr��� 6<ݮ<@�tSLY9�+vĞ)]}�+@��"t�ӿ�rԣx*��2�\İ?��_ES�v?�e���Y������L˖.��IYi7N�G�B��\6���po��Wtg=ö��D!偖�T�A��o�t�$v����`� �O3���V�<rn<U���UJ�џ�?�}C�7��D	��ҨU2&�p�*ؕJW��2�*�g�ϕnO��
0��Ǝ�9�#�k�n�0���_m��p�OcG��<��	��3c;�)ߨ?��>j�����C�5�|��[��6|A���N�@.�D|ń��o<��V��X��/~�,%�p����b�j}n����F�N�e����i��B�xsX|ր�f�2�@�މ׼��H���-����Gx�۱�2�h�����t��ݲ,d���������ٍ��[����"����%a��`H8��]��ء#��@��Ȯ5��y�bF~�z|��f�ö�|��g���N��B��'?l[YU,�-k]���޲�{�>"=�i/�X��\y<���1��rt����tEF��tU����j��̫w��KC=�>#|W�Y�� �e�j��\JZ�O[ȕ�'�Tg���{q:M��975���B��8\^��-O{��wp@�|��Y���<��L�c�7��t�g��Զ?e��2���(�:'ѣ�?�Ԛ��ћ�v�y�ԛ�g���c��P������_��9pht@%R��~/��XK������aB=?��`�M̘��p��������1� �1L��$#��B��:T5��~\��G�F*�E���7���s �:/m���{�|dM�P��&��YhЎje�$y�&g��)���@8)�����bmQA�7j}�9�ǤZ,E�(�pkh��VHQ�Pk$���zJǕVn"�Uly�� L��gϴ�o{���43l�r�C*��4��4_���Pq�:%��PJI��7y�.�NucV/j�Q�g<�ft��MML$�i	�N�$���`��d��5��}�.���p�i}�-!Q��t a@sG�nSV��&�E��m���Ty�&�Z��ZWH�_r�����L��q@�U����b�6��6a��\HHT|aƪN�YƇ�8��'Ǆ
������mƲИ�_��2��Ekq\k��:���l������M��� �����Ч��!�Րύ���d����*��6���������o��|�>��S >�^��:�S�*2��{�ds#���"��7CL��ݒR��uS`b�xX�������c�)���e1N�!�9l|��g.SM�2����(��D)��>�O��`3�-Gl�=��K1Z͑?oDf?Q�I)�OL�c1��g��'[�< QAT��l�R�2`B������Y��0�˔#��m�� K�Ailb�{��}R�&!�b��vmPt�c���@	u0K��Ȝ/G٥��xK�:���!\Ut���x��Rn��ze�/8$��e�Oك�LsKl[��H����[2��G�x�Ҏ���aG��B;�&/���D�����W�wB,߮6>�5��r��!��~;�ۘ$]��������I�[J��"݅Gk�;¦\�K$��Sve�M��مuܙ��.p�e�A�a�m����8�QI���z��Zw�cI���M��Y6�;�����f�z�n`���筝�V��������o��.�TD �=�V�t�������;l�.>Ԡ�!��Xu�S���[�V�Yй$.V��G63�~�L�k5��ǭ�ȥ�����2���v	�/<��R&\k���	/_=K�gc~��H��/^(���G�׶�M�+_�ͰU��&��='f���.�HMK8aeC�-��t`9��r�t�c�c��������H�����2BEE��\ΘUq�H#���qEeBMyQ�Q�B^���u2�l�D*%f[���e�W�ė[����ބ��w�^ ������� �Qؽ\�yIOxY��W�@P �H�8�q�;�3��G�7���*=�5	@�l�Pg4����8ރ�d1e�IIM��zs=K�h��!0޻��P��x���4���+D=��=�G0c��4�r֭���3ml/����i���㯹n��n ~�1uݡS-OQe1MS/��Q���s1΀1�5�9���!� C�9V�Jh���G?G'��BR0;{�B�����Yp��n�c�%Bl���$��ᣤ���	< ��ܻ'�[�`�o} L$�hk|rHt�����=I-��\�~E�S��l�ߞ��@){vm�y�F�U�6��@�W��ɇ��պ��"	/ 8895�i&��S`HD��v������@��T�
�Ƴ�{�:��khi�1Ӽ��|����>\T��,�z�䮅)<�Q�@�@W���k���ܭ��z��n^�o��C`{*���xS,��軑��Z�a}�����P`V���µj�Jb�:V���	���;�(z
���`�[0~(�.��`�eQ}W^�X��kp=�'<��>i��_�rL�J���(�0�?���*^����\��b�`�/,�=����os��"<D�ތ癣ݭ����Z��Q��`�2�}mu5�a��P�X�	��RV��
i�ͪ6:|���8��1�Q2V��QW�'Mɼ��r�Z�OZ)=s�W��R��#h@�m:ѫ��j���<�� z�A/[����<����믅--�i�!��hvRRrb���K�M�.�T��� +�7��A���������q`-���)�n��*+�=r�m��꟪U1��i��hw���7�U���a;!1��'DO���E��*o�B�RT��������̏ �(����d�H�K.�ߖ��O.,��8ߎ��U�W2V933�	�	�-6���ϓ�)��(�kߔ/�n�ųHSgI{�ǉ�������˃//p��(^O�`m�t�ɿ�|��ΰ5���傔��3&G�_�E�\�G]<�}�=l3���>h�zF�����_�ȥG=�D=Ѽ�IF:��ຏ�i�UdJ%xz��W�����9�Dv���t��в'ɒ�����7�=��j�|T�op�D/�"���)q��-t�{Upѫ��;#��q�삑���RA�Hhr/|� ���`џ�7`�,�.���WJ���`�υR��;r������Q�����AXm�\�b0�S0������9��a���b^
%��."�:��	��r�C�	rD���ꝸ<����#�Ǯ��fGzerEOF�v(�$Œ��U��f_�q��sB�u�-�.O��/&?8:��E��BMIX��H'�e�|�]����Ħ�/H�S�٧��V�l�/��y5�sq��j�he��݌/��y��Iӕeo� ����1���gk[F���c���q�2��9��K�̅4N�ݭ�ƪ,�M�.�M��b5��/%A�y,��wGV�{,�GКD��-�&-M�.��n<��hv2��\|XX��Z�A����9-bxxx	<E\5� �ڲ�OD�^ť'��Ȧ���"p��x[�[���˲ӭz�C܃:�ٵHх��^�<���0+�56�E/�D��Ũ��8���*`0 ��̃i���ϰ���bb�+&�:�Y�U���LMMkڙ
E_��'�Ƿ�0���Ɣj��W#|����(�
N��A�=-�e�A��>>=�N>0>���H����v�V��	��0Z�$*�|��f�ZYY!N��w�	u�X�."|%�YZG5�F�hG>-T�Q��uwu��V�}�J���;���م߼�h����өY�9�*='?�V��%P(T�ULJ
<P�:11�[�_���?��0^��>�k��6RY��	���y��y��G�x������u$�7��kqU�p�ş0J�2<�^�nh�	;zӐ���=�n����.P��TǷoy���7!����d�k�]g�`��B��d���Z�qh��X^�� ��'�b1Ñ��a|$��lCԝԟ�OM�?;�\1_�b���j^7jd�N�y �-���x�A��M�d�zhϡ�9Ɵ��ADh�k�CZ�hj�v�Z��χ��q�=
,����������L�2˃XyM�8(G �eB�ج�o|��8謼���w�kz�����[7-�3�%�r�s�l�KP��_m6�ub>o7�
��#�Z�7hU��<�'D*R��]ID-����]��B�6%	�iw��}۲��� nn�&����f��D�������e�\j�ty��[�Φ)�ܪ�:�,�}��L�P����zY�c�ɥ.z�P�H�����x�#�������}=-44>��_FDn�6N��ʹ8Vv���� V8,��H��J.� ���|�g�5ӬH���mJ�WX�}��6̸�aFk��}�o��FE���H�B��Qsp�[��h[���e<骎!!�%��v���n�g�qjמ���/|� 'i�#��8��nG�`S[/]�E�$��']^��Lzw˥���z!ºa2W!;����~G��O=�����?}@��	Y�27\<�%¢Rv���e0�9��B�]��\����.ZLwE�c�D'��B�8F�}��{�F��g��Jey��Y����l��}GV��uq�'�G����PݕOW��:����G����R��T��=��kG�$�&&JZ{.v*${�{I��S�ӄ2'/�NWRSJ��;�A�g���ݨ-�����y�y���g���
%��R�@����U��z�f�9�����#j:����e㌲������9>i���7�z�=���_��p毒E������f�T��w���a�G5������CN��D=�����g����f���_��}yX���1!�95�3o���_�b'<MWfh'��-�y/�ԴC����af��s���R���>׫�x;�>(,�u7<P�д�1��[:!!�݉苎��/��۪��4mu��l�I���)�}xϤ�۸�.��d�Yt���td`#W���Q*k��X"�`�J������M�d*#uK>����rb�3&* ���)v(���fW�݆�����=WiIt��w18� �`OS�J(V����$�,11Q� �����&�fACv�|���p����l�~��Q��@C#����s64�Pr�������{l�s˔[ �����ZxΈ��L�ݦ�$��h������|g��ǒ��@:q�����n������}��#����=�UV�� ���Y󈉿J��8���$�����4�H�	�hD��v
�/�^;\ }X��N����\7�z�����<P��`���Y�
���iH�98��[O�ݾo;1��	\)Ml	��sp�[Òz�\�'Xt��#җ%S�b����6f�>��uu�tŦ�ݶ����mW{qo=�༴��2h�׷<��&�S�;:4eh	1�*ߪ﹌��\��lͺ��)z��0�w;�Vm$ ���Q3�p�ƥ��o�1����9�����K�c����Q�v��2%Ie�tl7���\���B7 ��a�?�!�a������ٖ�P��8����|�
���1=ey��#�%��O�p���)^f�+L�
��t��.�� ���
p].�L��f�{0�ż��@[�`���(DN%'>�;ʵ�?��.���LBЄ�����C|�t� ���H8���-l���x�B���s����>�)CS�O��#P�y䢧ݨɻ�'"��3��� $�|MHXrn��ˢw\��!Q�=2E��7%e�z�q�jr~�g��.���a�����Z����>���:D옟@_�n`OJO��z��	eD��A6�9�*C1�o���G��W��3�w������U�G�^���)f⤭�<�\xǦ�[��B��^pD����7�k�!b�/KA�_�^m��1y~x���KF�-�g��ٍ��������Є���I$Ȩ��P+�q��S��D�m���h�Ք�@ ��\��{0�Ii�Y)��sTx<�l�A��DS�g�}�o��~~hHy����/�(N�0��x�0�O{���9���@&s��i�H��I���)b#3�M�/�����w�}�D5�8k��z����u=%�u;��o}��%vrŢk��7/������_�y���Jּ�b���(.4���l�(��U���6�~��4�'�E�|}���d|��X�R7��lD�׊�nO�ybY���vBd'��mB�@ߔ"V�-sel�Zk*S[��h.IG���ąc�KT3ڴ�Q��jWrB4�c5*�N���o��I�D�>��״�?\����V���
�h�M�r�)�8����Ѣ��Ngۘ�$��$�PK�n?���C}��7@�^XL���
�=_�Zp��P�hA#N3��@<���9E{#C��I�"����v8���9�UD��<j�EeX��=����yl��L�~�z�7ڬ@���A����4�i7;�6VO?��7P=�� ��zB���5�m՘g�)M���|�l�շ��L 2������ax�V����>��>}J~�/��J"��#/"_[���@�� ~�rk��K���i���iưe:��?��X�`T)���Hm���s��; �k���!Oc(�����zb���+ybl�?��'4:tc(�s?��ٚ�|��cv���H�~������\�kg��Mڮ3	��>Ҿ�~��kKI�E��.�M��@Ko�e{�Jj2� �վ0�P�?Sd�+[FS�͡ՙu�a�!?���7(Ȓ8������K��x[^��o�o=u]?R�������V����U+�a��3�gJ��D�]5��GS3jF7�`lf���uH�Q���K*x�
C~]O�܅]�z��F�kp�ff�?�b�F��
� 7E|�7��1�@�	�C՚�q2vU�F���<�U�t���a��Ǆ��s����2ɀ����2��7��]�!�+o����S㍉� �''�<��k�_��U�%�`~��cgSŗG�0�/�u�t�3p��49m㊿"T�9����2�q��Κ�}��T���e�C��N�Qr6�nM��<w��eLp��z��
��I���{8��l}z ���3	�n�(�1@���3�u�[s�~I���􌱦�)�L�����@��ܴ�|�Y{��|}}�����5d3K�u�7�����/G1��5��@��_��5���^ღ�W��+C���Su�Zz;9n}y����:�W����8C��;�n�?�u����������d_G���Y��������w�k�w��V���wH�Y�Z�#g��;�*�L ߣ^����l�O�D4ey٩߉D�����В��%[��BsV�뚬 �q'��C�(��_����g�bʟO�q(�^okl��C>��4ט��x1l��^7u�vwݤ�C�;�Y����I���p/��4�@T1·]]��}6P��[�1�z�ű6}gT��Br���j=}�B���M�Ok>�_<���O���%%%)��LE��7�G����ݺ�ļV"�y�O����6wv���-�m��hXk-M�B�������ML��Jl��$v��<;F���Ӈ�,��bs��}�D6?*я�jI��Ե�RYI�/��� ���u���d��xe�X��e�;Q0������-�^	E���;���:���5��ıWYf�J]�M9V�\L�L%�������?Z^�O�_�q��ʗ
n�\V�������s��]W��.�ض�i���8�N�9m�>�������I ��Q(�x�y�s��t>���t����K��� S+x8x���u���o������X;E��1����h�Y�$�ϭ];��>�	@�C����EӺ�֙wh���.�]���T��B�V�H�i�����H��wO�ۗ� x� ���n���w�&�<y!��c��)Z��x�q �S�x�2��_u�-��iwX���27H��$ ���\q%�U�xۑV���8�t�%�10�E*Đ1����J�6G㵤gn���6��B����� >�=;�
�N�)�Fه[p��!�V��V�tL�{�kGW�/f��{rc+°�C'++Y�`� �8�����?�Fp�)�d��#,f����������8IKK�ى�

�f��9�+�G6���4`����Ht`
��d�Ϛ����E	JJ֚�����Tz�6�Ԓ:L�����{ ts����=[t��{�U11�D;��J-�C��t�!'�}n=G��)ˋt�㶑�8�:�S���^w�\;\{���V(z5�
=�@�\�#e� 47�C�Rb$� rc�7g����F�ͦt8fN��u_>�"��yQp�x��Ծ�mӖY"Yg$���n�\�<�'*Z������P"�`N�,��F穲��5��#ז�����D�kh��WoW��몖����o3pi���M�?^�W�08O C�ı�ݵ�q��췇�M^�;f���{���d���a]nݧv�^b��o��UF��BEGI)���b���4� ϰkS��ݲ߃G%*U�G�
��Tj5�t��zJ�ޔ���z�$~zL� v� 55j@�4�t75�^?�9ܲ�j�.��ދ���0e8�K8�p���%�;~N�p��Uw5���r��p�ȿ�|{��\JUT��5�K�Ąu��wBC�^g����fU���.R�i�_�N�^4��O������͗��k�l�Sq�V����i[�_�7z������z���w*���+MdG�gO_u�b%�<�꺱N��F�螣G�@P i+��@I�1%y�=H�������Z�7�2L�.��2��g���n�T=,t�-!f?)3�uY�t�R�9���ԝ۞��8 �a%@B]Nc����h
�g`���J;�Qnnl���/T�&��4�e|�;�+��2A�w|�q���i�Y-+-� hkر[z�:��I�9LU맔κuh�\�Y
��t�����V�E���>Mڟ�y*�^�/�h��׼�p�}�ۀ����ŵ������ͻ]��������R�?)(�����+2I���O- z�(���iMXZz}]�����~š���&4�H\0��CUM[�C[�����=�`�/i������������2�_��Z���7�7qڧBi�ox�O/1����>�uW����wo�il�}J�X�{y5X��M1��������~[��d��MIOQ�ǥ%�L�Ώ�ф|? \�"��qV`c��OVC	�sQ�ǗkQ�;q �Ŏ1_�[�:�GNn��ϟ�3����$ Q�s�?`E%�)൮#��MRw>K�Ի�K����5U�!�OK�J#�Ȫ+�a��Q��#� �w��m��+���/oX*��2
��O�.}
qt��L���\�E���X`�o�i��������QQ�_��H���� �݈ H7H�tw�4�-=H��R�]24Hw�=�����X��5Xp���|���{i�;���c�.��n���,Ro�J�fk-��J�m_G�8P:�+�k��0
��z�D���cn	�z[q`ٽ��tH�����ڔ��/t�{0�,�=�Ck ��n�H>������:��ѻ��w��7ʪ��'����h���e7�tyqO�C׼p]�v2��R�y����������511����$�ˈ�i���ƻw���,�|��,<=S�I�|�������N���3Hm��6���}i� ������G�W=$\2$x�#��J`{��N:ۃgX�>��HY�׀ԟh��WYë�hP���j�!��<�m}ML�e��gy���*�z�]�;O�M�!Ȫ���Ի�yf�l�	���,��9]s��ۓ�X�-�Ow�jV����}�y�U��D0Qe���8n܊L�\~C���?� v������6"�	pa���������?�3���X8�O$R!E���V%M��;3�7�_�k%�p�.�﫯�K�'ةUe���~��q���b�z7X�J�VU9~>��x<�\��\�L�ч
��h�ri@����a������pY������ZU�0��sK�A�=�����Ő�H T��! ����� *�-����OOmmЯ�ƺ�Sv����V��|�����uR�k���m�4�b�!9EDY���J�(�z���S3@1�lK��E9.�����];[69�����p��Bm�����r���Ђ~f��;%\��Es�OF�A�����b�,SL�i=�i���eqs_���(��g���(���Fb��3�=X��O�LYC!���lOP��Z��83��l�2�8Q:i4���2����<a��VO���.����&+���"s�N\
UG�S��݋wR�m����㬭jj�y����+���\�*�Se]��A/H�r������ĺG�B	d�A8��c21YGxn����P��Sl#�px��5�/8�ٔk;TH����������]��:��Ǜ¤�16ğ��4��W���E��vaT���B���j��H�>����=|��jjv���#I��Q+�n\�j�TWm�4J�+���?U1lL�d��.? ��j���	��o1%0^e�u�����o�>��b�H.�ߓ��=�6N�� � �Ι�ݯY��Ϯ��q�ekN3*��a1_��KMÃ��LS���*��dBv��p�n'������5��`�2_����B�[��y�ns���v���ߢV���e�D���~�����&����d����>y���q�� 1�g��ƸV��tQV���:����n�Z$s�s�k.gb�^�[�h�5���f�n��o�W�)�:D�T�o��l{��n\�z�&�眪��Sĺϱ��3���s3w��㚿�%4g��]�=X����|�t�j��5��`�PQ�͉�Ԃ��Z�¡�b'+NΟ[��uC��'r�c*l�		��M����
)�����J����US�	�dZs�c��^<��c~gyh:K�J52��dԐ�д�����V�pv	$bpP��� ��pƗ2l\Q�����+�L3 ~RǏ��h��t4��Ŧ]O�lQAC�,�16U����K"�?�ų�yb�۾�n����YD�6Ɖ���;���A<�_4�J�2����O�]���-X���c��R�Z��/R�Az��lߌ3��������4B<��3�;}��4R���T�ux��5�"�'*#^O�g�7B��׆�/z�>�������@4�p�@~�8l�L�)2�q�DE�Ţ��'ϡW��U�|F�UQ�oP���ob�S���c]���ը��m�X\��Ax���'�?*��f{>�\��;�t��Yƾ�����$����!��]1P��3l�Bz�&$$?�ۙ�}U�$Ϝ�r�r_Ub�C6�'"eS��T�T�id+���w//���_zm������/��Z���v�j/��Ч�C�(5�5��yƦ��UoN�5Ky�]5n.N�mOw	�������6Aq���s����
�mE��5��G�>e\���Y	Fe	�w�%��`�����7��iD�|�\���>����*�A
��-���G��O��B ��@W���9�o�'t<;�E�:I���q^�4�.����w�1bQ��9
� SX��{�/�F�s�"�&��������qr]�+Wttt;oN�N�ZX�8e��C�ɨ+F�w�f�0�qk�Ӳ�1f��^��e�% ���WK����o����F���	� �9QҩS��9�;o!ӿh'\<�$j���ג�:;��5�>��_��s?���̆#���ߠ����G����"Shf0�ve�^���S�Y+�*4s=�0{B��dD��_�(�T4�PĐ�YurJJ�����BLL�
n���
&h��.F���rIF�jt��=�C�ʾ4��:����Ҥ���C��ސ��;'�c�p��]��R"RR߾�!�j��	���Y푩u�X�G{����{�,J���hk���.���������8��֖o��\��
��+������QZrϣm�^<?l'�0��Q���n%s��!"W�"��M����Gc��Y���{WBֽ�&
0�J��ތH�2\��`�X��n�[ėR"��|Q �P�H(��7ˢ2D^T�\W3��/�}����-)r5��2>~	s[�Xӿ31����p����z��>(����6����v-5�tA�V��G��("a�G���t�G�K	g��%$��E��=K@��{���TTt�+��!�VFg��1>;�.N
E�T
�K7�=��q&b
�l�u�"��}��>#{�<Z57!����н���t�Jw��ۖ������U�'n�il�ET�� �������Ky��~^�����ϒd>x"w�1�n�z;s�� V��"��"�5�J��i(�q�ˁE���/�Q���K�_��K*(`�2�44�#{��w�����u��S��_�vz��ccc2w��b��a���"��I����/&=��'�5�]���:���
VJ�o�"�Wn.�/:Dn:L��+?kNp9"gH	;�!��)+�)�2��w}�I~fS�թ�A�����s~�ޙ���J��#����FB�OE�����9�_8K�^�9�޳���\z��sً�&X��ћ`	@"��������Y��#��
���[9q��&�u�Rd�_'M��c�;��4ajj
{|��ѡ�h�Kc�ڀ<Gv�.�Z�>v!��B���|xl�ӑ�l�".���	�t�%S�;eJ���ĜI���NQ��K�+�ٮ�z'ۤ���o��)�}�/:c�U��ĄC����uCƻXt��"�y=�w_ J����v}���~����Z/�AdNgˑ�[K[,'ҏ�w��~���\�� ��C�6�7����^���M��ԡ���iHL�b,�\I����K̟�q�"ݮ�7��=�b�v�D�0 �GҎ.��V\_�{�͘U���R� >?���$Q<�<�G�7��8l����ˋ��\�>��Ҏ�+��y��)<�H
�:\}��F*ɹ���uJ3F��9v���F�֪~~��s��g����C�:\���>JK)4����q0<:�n�eʀ���L�#��j�A��E�B��L�mR1�a�S�wT��{����ɚ��Z}�z�@��c�X�pJ�V��ML���r�VDU�.)i�h������^�������׭O����B���\��1"��R$N�J_���ȊEGw�_M	�u�ϛGh��.��E�b"ަ�;�y*���"]��!��ၛ����ʈ�O������;���6i����OTp���@��5��y���N��?ے��k�	�)N;;y��D�,�5z;��^U��N��_�M�Et����q��i��|��e?5LEN�c.��_fF�5
i�0e,��)��BTD$C]�a�l:x�ͧ
3�X.k�#��	,���D�c�첅'������"�Ps��{�}�ފ�nӋ	#A�5�Q�m⓬�3�D�i��J� �!�G�w����6��x����|��^9�h�~.�=�������KӏÛ���2����Dz��w�r����Gk�G� �����0&���+�0��.�l���I��s�FNV1����`U��h�����p��M�B����@���V΋���f|f�o���?Ǆ.γ�n��2�y��OuU�ڳ}&ː3d�E`	}^��ó�}r�>N'�7؍���x��]�l�}@��7��I�lez��i�f:\ѯNk|8�O&%]�PL%�$��Nj���®F��
�w��.�~ɉ6+�����\1f�c��]��\+�˰`����l�̢7c(A�4^��n�i�~=�01I:5Xe�$�ڦR��~�C��݊%n�d$�ٸ$c����U�.����o���Om�0y��~�Y[�ȋp�4B��a?��Y�?�z��~�n��?�}���弯/�60F�sI�O���E���/~��o�{	��`ϻ���^�ę5�@����	Cb���CE�]?>E=d��c\P�hr^��������/�b6,W+0_
_��{��'�<�e����U�?�mʦc�/��9�p���uzk�˥�2�«�����*���"�qY���Ƚ(�+g{��6�ܿW�9>"�5��+d���~zU�'�#4TȆ�\$|<��G�M��|g�P�����2��czD~���1�W�(���]�����3�J`m���2D�����S�scp�D��2�& ڡ���k��������
�E.zx����s�5s�f����v-'���W�c�g�-���v��a�A
ގ�w���kA�
5��Dl��7W��w筧'��7w��V��=>����{��#n0-z���[|x��𘅸��\���c��ӋlE��-|9,!��G�
�X��+Gهm��\)9�>��@��z��Z�6��H}U�o��_DtR2�9�^*Ȯ�g�Ǽ�@a�\��z���#�c:����A��N��� W��h�)�����r�h�RS+_��U�Uj��:2j�d�/��4��a3����:l>q����
xB�G׏/�c �_�ίs,&�VX1���f�	Rd����5���;ׄ�q*/G����Z���h�B�l6, ��'�5�H|D�U���R{����5Ƞ�����u6�qC�Ƽ�窢���������+�q4g����(�Vjb���5��ev����?4�:A:G���悼	�����w.���棍T�~���q��1~\"2R �/�~�5�Ԝ0lz�y��G� m��K�i� w�K��^.�AJx��#Q��]��'��%�+צ1?CbE4wx}+�&>��HQ�-��o�89#�sgǺ3WD�#B���U/�SY*B��-�*���!B�}�:ZC��%*�W)*��z����䴴^m9c鋝���:����A|�n\8]�7��qZٳ��_؋̏h�T�%& �E�rp7�(�"X�1>�*�Z$��R���#YɨB�ƥ�)��c+�tZ����_5^;����f6k�����܌��H��>�^�::k������'ZkST̖�	t���<�hqb8@WW5�d!K���lH� �7-��r���'T��z�����r+9M0~)�
:h�>[�G������{�J���TIWW������2\$-����B˯�ηߞ�/�6�%��󅉡�ll.��p��׏s�˱���.'���m����#��'��A�HY,���.�]�P��Ȟ�0)nlF��ٓZ|7�l���#h�t��uk^��aP���)\z��XO��,����yv��׫~�Z�h�H�����v]�F\>�嶛�b>^�zj�����A_"3��"��`|lj�'��@\�x'mK
��a�o����Tgg2+�@6������1��łW��5w�XЋ�X�Mܤ.xT`��l:r�utE���v[+���[�{c�uo���������KՌ�׏U�ʦ(RR-���X���d��_C�'ss����>�,׷D��bff4�_��"���l�oT��eoi5�����&�]�����6F�&��C8��(�D�S~r$	���������]�A/��X����G�zu����D�2R��J�c��kw5iԀ��h�j5��W�o0}�ND�ד���U�������W�̇i2Bw"w]�PH��B`c�MU7Y��4� E2TI##���+�7VO���X�:u�)h=����鮪������2�/5}c��*;�X5��ev��as��/-P�ְ��5�����;侓i[$c\�urv�\�פ����2޻��As��{���9	� 0r;���:���D����iY?~�w Ʀ�N�¢�u�<�j�H�'�lCՖ�����g��|��ࠧ�?4	%VVV{9�����L&%r�e�8��H#�v��R�-�S���g��d38��ߖ��8qCmS
�ݥܔi�1{xYY�g�dM�����s�J������(�Q�����z=V
�"�ok}�[!��_C������t|y���3��N�b��"�adg*��.֦���궻�'D鑹�=e��D8�^��状������_S�;��e	�wգ�H�}Yi��@�6�<�������*�./��6 ^־�Pe�Ƙ����At�S?� ��7���*�!�y5=[�F�\T_?l�a�QJ��
#6�����pu]t�/��)��(�1hZ*�sg�˩@SM���S�yjH@ \: V�INcg��_ޯ}�%~.'��x���v1�_�f���.|�פ]�lw�.��>�����?�H�W=�����X���~%�Y��W�gb6e+'J��P]天{)۾������#\3]h?b���K/�X�5�l������Lu#:�H�:��W��ل��m�����Ϣ��k���﷪Dx8g7�O��x�
7'�3�:W��`JD�dݕ�(0f�F�f�����hc7��G"9ش�JW���?��#���?3Q��ظt|	��{���a��#��H� QfF:�w6���o��6Z�rE�*P|�o� 3iLn>ЖF1���%1@tF_�RƓ��?й������'9qY�@�(<��:�����=��9�غQν�ڛ��5Zy� ^�`���_�b��v-�������W�j�ou�2�q��hf�s(����p��ʫ����}��h֧�f�zkgǂ'���I,�vv��w���x۝��Ү_ ���Ct���`�/>|�^��	�Wo߾@e)S$|�U��|��Ƴ�gE �[��5�/7f�;5����&!!�k7v��d���":#@�2B@�P��i��!�]WJoػ���9�%'Һ}��42��k�4;Q�6AJ�H��򾖩]6�RT/�]Hj�BAIU	�r�A�@�N��(Sd������P�]]�k2~�3���_��L-x����`5��q~���h���F����b��<���gg��aj}��"�B�M�ڂכm�2	Ȍ� �"O�m�M0�	�R>G5�.��z�w�L0<)=�䯨!�}����Ԍ��Ы��E������81�8��p�t� ���Zy�x0��w�8�Ԙ�qqh�g��M��]�K?�ڔ��V���5����|����{MM�Yfy�sx R}pN��Ki�|�ϖy�[�qjjj�?F� ��I�õ��6�G��]}{�)�?�����ʿ�"D�Z^����[�e`��l(#:j��1�ȼ��ڭ�+M#�/�ܹ���坑<����%�u���s��MHϐk���^ �K����禷4"kR"ᚅ~PG5�|q�ٵ:��h؁Kn�x`��׍&Y�9�L�'g_CH�:5L�4��2�e�xz�\�1��TX_�	wN�Ӎ���ߌ�E�t$�;��@ԡ�r-/��^�ϸ���z�8Y����T��5����{��e��ܭ ��F;;�-dK�V�̚�(��-�A�Vu?�
[a5c��fh�0��Fq��(���0�y/�_b�8%���~c)��E�]_q���g�}i/�l�y�$��� �ky�7�5�:j��k�!��"�H�הo]7˃)Ajc�'2%�Ǔ�3������+�1DE�|6���㚅&4Y;2�'�!�$�Z��0~r]�]�kDRΤ
��v�t��G�z"��<;9Ǧ��=2@���Ҵ���jE�KPH��6�K�uTw��D��%F[gR���%5���fa��~`G�=��r�����="Y<dھ��kV��Q�{�4}�r��"ML�����ҏ��pF_=�.0#��5Z]|E�� %?�c�1�����=�6T���]E]1��M�`h�)��t����;l��ݳ�4k�����0;&�w���Q�d����7-�[zܜs�3�1��MO$��<L�r1c��T�\u}�@����,��U{bgܹz(�\a����a"Z�s]����dh�b��[q`���X��W8�u���Ӈ~��Xx��Ժ��A�%t	��(�9�\��8��ޔ`�Z�D�a X���w+��""��G O/�JTJz�J��p_7HЋyבb���(���c���۽�cX?�Ci�ٳ��A�}7�oL���C�}﮲���',B���-�,���������'
.��a�J�[�-4�d����aA$54Ԩ�\�B�8He��tb����kr��U�;x�K�y4�}��e�Z�xy9l��!?$�t�$�$=Z��d��_۱j�c.n��0l�{B�����PR����B8����-w��C�c�w�?|�6It�\�n���#���:���|��(�3�b�Ю��wY[rսYUWR[��A�vu'�_M5-�|�;�gh�?�����yuf7Đ<!��0_�Ȟ[t�g�w�q�vrZ��#��!Q��m�YO~����ֱU��5{&��!������+�(#xA�Mw���8Q��`#�{8۔7�:�HR������Uｆ~�!�߸��w�e~����	�T{8ʗ�/�ł�x3�Vt�Nmi���ô���$$�(��/ϰ~Rǅ���/l%�F�|�T��tk��\�D_𘛳���c1��Z^hh��e�;/��H��j�����܏�֕�s��wW���w�[o2�K�ھ��tҎ�L�9�ϖi秋��{�����K-n��y�L���d�8��[���v������9��þ��!�c��*zI�Ym�nw�J�tuZ�?Er��~g�2�L���>�`��{����1[��0d�n�ϗ�W_y�Z��SE!�o���v�yTz$�?M�N�hV�$���U����8�-�������y�}�Dj�Rh�.����%���N}3�c~'�wr�8��2mY����������濲��O�J����^�6�*�>품�=��(����z���L� I��	���`dܣ��f��w�*���,�.o!6�(� w���;�f�r>>~�w����Ǜ�u:�P������pwe/�����_�䛱,�,��5��j��ɺ��x�pa_����T�$�1w���]���e�tr��U(��3vJ�&-Gę��� W��}�sњEV�5�p�i^��5��hnqm��l�K���ϧa3��{�lpim��l��LA	�H���v��jԿ^�DL�Ǝ�̰�b,е$��j8-��T݂�g����@J�%]����qMJ��;�/�{�2���H@�������C\�m�{�?\�G��P�B�}�_e��w8.�e�7~��`b@�4���o���P�}�i���XѬ�^w�}�j��L+��o^�\�
�G�s���(��H��퀐l>(L���Uw24������b��tĽ��K�_taPy���جLe	���b_s��?�a�߱'޿?��K�oЍx=��Kv�Ɓ��4��P�L﾿"�a�$�1X��^��M��Q^u�bVFS��t��n��1�[�vU��Κ�{,��=��yq������Ⴂ�|��	�5k�I���&3�4��~>��|]B`�l���8zS��j�����R,�Q �5�̧�B`����am2$q7��:cA�|�:&�g�9���F��6�KIoy���il�EI3�$�G�N�_�y_�������l�d��!�8��*C&���Ve͑v��U`15���Vc=��o'kQ]�zL�֢����<�	3p.�&t����Q�9�S����@r��P��{���w.JΡev� ������d͜��M��|O�v��x�&�h��ͮ.���	��֬Wɿ4�~8#��Hڌhu�}Y[�BҼ� rV�����u�K�.Q�7����Y��`\��I*��b?(?wJ�~J;�~�Xٸ���j�����O�3ow/o]I�7�Ԃ���Q�&S�O'`�
.Z����]�.鋴\���ؗ���`���n-��7un�H�XP?D��-P����v�ц0�)C|]Wdaq�o��p�S���j�;�� �}O������ɸ� {�njY��o�;Q��'�F)�_�Q����B�3�NK�6��G�wϦ����L���������q�E����l�i3�j�ژC�����c����l�瑟�C#迃@�����׳���-�m	%�0��1�~5Ta�Zñ��-�<��;��L�V1y�i U���e�g�"e`�8�o0g��Kbq+jl.��Y����7���pE��;���1��*�.��I�A��%�IZE�ngc�s����Ǥ?�D�ۜ�f7���5�4��S׬-!���t|���̀ϩ�yĹ��5[?���8G���Iş��]xyh�zY�cu}D�Jz��>b�Рv�'\UB#�q��8�`���Z��9ҟ<�׈��u�����-7r+�j����yoq^��l���Y��ۙ����E��SpH�%��+|ks6��� �8��X�4���W��s>��*�����.��n�O��8�ķf���H�[!�϶��NT�d���$�_��ƈ�T�}<쥅h���3�?�5�F��S���fw�� Kg١.s>�g'�si޳�La��7}Θ��� ��y����|�_LOG�x�{�9<JMVa�{$��jⷧd�igxyM�FŎwc�
i�߮�@�ީp��u��Ǆ��Fn
('_�a�9F�������P{��@���'l�YU}L�.��a�]�M�-��K��.�����I�-j���0Q@Gv��ז\r��䞞��p�h[�_�J{;��e����=%����l��Y^9�+	������O<p�s���h6�"�{u�����1�'�ô�G����}]����A�����?>5b���n�[t�~ϊ�������
���dcu����I�e�Ϩ�,n{��U=�'�I���F�E�ȿV��%v^�� �X��օ.�~8CH���|�������ˀ� d^V}� ���כ[#փ]
,)��:ߣ��6�aH��r�_&�����a�2���4�Kc���Hz9eJ>�}4�c�"���0Y*�7���{�n�MXq�9=�-@�VZQR���h�/�{�8D��0�,�uw�P�����Ѥ�)q):�|���ð���	Gyj蓇h��4y2��b𵮐h���I�B�������"�x/ݓa�������Z�k@��Z�G��	�3��k]��0�?�6no��3��l�2�hL=Tk�A]xMf��O�|>��u�Z�%�==\����L �۳H��y�e\u����V+��ǝWBf���^Iu�_�ʃS���J�qQ&�*.�E䁶W�tp
�I_�4yx긃��C������,ѩ�N����5M��9Q������������-��
�@���l���Fr�C_���>5jRR�����XU����阬k�{�ǶR�˓�ۗ��9}�R\���#��,_wʙR�`���;Ƿ�����0u�	�Kcxbx��¹��1����Z���wv���@�[����ġ����O>�T��\�K�=��av���S.�n��%e��P��W���,��S�s�f�B�Tm���N�޾j
Yh�!jk����y$;�o@;;��N{!���
\�u��Uڢ�9o1�T/������ZZ����V�ˁYtX����h&l���@<I7\)$�xʢ�^�vW���=�3����O�a`�w���H(6�����FK8 �C��������'��=���\�OhJ�4�FEq)ԝ/��޾柭\@�gSu�̘��'n,���٤h��W���,6����;�/dFA ���#�\k�혣D��.��U��Cc�5�ARW��Y�=��O�������/������-o���A���H��QNt��^��
��<V�*��a$ �K��ۺ=�X縷��>���v�����o���$	4�pQ�sc�[��qw���ߌ��-�Kj�.���˧�̩Ӛ��B~�2/P��ʗg��!����!}�Ãl�w�j���'�K�=)囜C<���WFng�`.��˃����%��u�ձ?�_�����F���ξX���̝��G������k�K\�lK<Ǫ��r"�A���;��=�S=�.�M���c+0�n���Ka�AvS�G��m�TI����.@�C���䖦�f��k;O���k0'/*��'�K�0������;?�y�qlk�)���k�Mߧ�"��F�9��<jD34n��H�ˀ�*��Q"Z��t+�W�%��63���pѹ����H�K�VM�<C�t�o��Z�墺�
ɧ,�IZ�yET͚P�z ���O�E1/����7$�GVvT�n��F�&�L����@��j����ۢw�&)��pA������SQ1Q���j'EF�g�����o-�����EQ,V��"��vm'ME�F'���{=��w�o�~SZ���x>�+sn���3ܻPB�o,զ�/j�m�d!�t�m�j ����B"�R�<�.y�����>��V���~���̛��8ʬ�U/�AI��?i��x��o��5w�U� C��⻝C���o�qpWRNc:���v�ը>�`�XD�jh��W�V_��NH��b�1�Љd���&�&7D��+�Hݣ�� :Nc�����3&>�e [L��'���@	����K�R2�)�\���g^>U��U���Yr�|���|��ٚ1G�]C�n�D�'��F�@�� �i!�wX���i���)����r 9�F+�#T�h6X�P=��1;��uq>�9#�j�!��kud����;L8�s�&�! ����%�"�Y�B�2	��;��_�fVlu�tŷ�Ǫod�VTl6)��i,�l
Ig�6����k��@���;O�� i��V��-Z����Ih��vd� ��E ��X���-�<C���� !��n���2�߁vf��G���c[�$�3��n����Y�#�����E\{����A�ƴ�������)6��Y�%F���!P�5�K/�p9���l��IG����dc� >�����-��^��~{������r�}�N%��٣���k������w]��('f!%�;z�fCi��N�b�i�_��
�7�k��|/��W�Qn�6�W��;���&8�\�3,�%m��{�˼+D�奷���\����C74m��;���r�[,c-~���.�֓j���F ��t3��gng��-�cZ�uק@��cHjܢ���'}]����I��lV�����e�zNp*i��6�,�S�+*ixMn�!m���I��.��(���^��+��:�ax�[��wx~�_UOz��'�L��/���{@9l��X�<F�����h���/糛��;U<_ۉ���r��� ���5�V���K���3�H��ⲱ0�լ�P��m���{��!������Qjq�$�`�pM�J��/)V�p��2�wH'�����Zal�eA��)=�R1�}K%`�C����6�?�S����ߠ�~�Gb�J��t�c!����$V���n��L<�yxl��)�\���i�U��E[��ʚЪ�d���i���ހ5���N�K�c-�?:� ��KRW�pPU�)v~O@��������M�R<�Lk��t݉�F��nBLA�l��볽��]ܔ-�Np�Y������]Q�Rwᔟ���4M�3е��4a�B��u��Bny�-����/�\�byT�*����	�	�]�tC\Ѩ��a&��;�͸x	��%���w5�������5��W�8p.v���U��[/]旷�N�)������R�u�����t�ұ,o���KX�ͨ�S(�\"��c�n�㯩���ԡXr�tS����eޗ�Β�J��C`_-���%�}f�iRM烤��.{(�J5��	�d#�
�@�ݤʭ��N��Z�A�X	"��cMb�H��dcĽIdt���c���x��Й�|�L�n� �2���WJ�6�~m�#m��p;{c�ǧ��]�{I��y,)�=<� ��-22�i�(��ä=��ܰY����om��@q��ޞ�T]t+#K��v�[��]~�Ud���`�k.�����T�x]��hS��:{9�nA�K+�R>	�eEl�Nu��V�<R�0|"K��q��U?�\�Q5���zb��,��0a�ݭ��5z�#
!I6�����;��{L�k�a�Q25{��e�wH,R�H�D�h�[|	���=%L��jm�����A�'��ҕN}��"�V��a�>2 ��Ҫ��CB��z=�� j���ya�&kR�/ooKm�t0� @�7zDl��l��B�wHF�\L��O��l�Ko1�P�~}HN��}�"�.(Y��W�x5D`���EU��%o�F��f޴  ���y9�#7˫��d�:��g��t��(iZ�`fH^�X�������]K7=Y\��IE]�[��@�Q�@��ŝ&RYJ�6�\�I��X�/jjN�$W��ݺ�/¯17���d;x��D��@���9�t�����A����moF�7�7��b+I�߾^�Z��	hw�=�M�o�B���`�?��茶���h�rH�\p�[�o����ܼU���|�xQIͶ��_EM4t3�7��C3Dr�v�s�����<��n���I��� E�sU�\���3�@x�#�[�b=�-@�2W��-M@@����������})��^����d�ffeZ<��5[g��A�/חlO��<��_<�g�t�̹8�������䊨��\���H#{0)O��
��\lݖn���s�!�\�A���7��)�vj�C��^��\��Ms�f�lr����,��:�H�7a�o{��F �Q#ܟe�aͯ�"��]�?�|�z�>H��=�F�«��O���jR)��GH�����{D�/��Y��J�(���B	��"����^�&|u�Ҫ�	�] ��bi�q;*��|Q���|$�PD[G�E�Ւ��*�z�����͸06�E���q����l�uƎb-Vj��i̬��XX��V<17[�L��mh���9N���uj��5g�Q�J���q���@z�k�
65n4K6M�eҍ%���	G��E�򾫠:`����R9$�'�~u���_�>�>u��ܲ!9�ȩ6ьr�>�&��ۗw������[��\J�ŋ;�w4X�{��}��Y�U6'�L��CP5�#�=�3��$�0�>�O��/�ْN/�=�/I6�9��*��թ0"�kjsY��+��KY�C�AB�❴�73��wܳ���3b~�Q-H��
s<��C�����`�j�u��ؠ��V�^���
�$3�>0�l�/���y���&;��J�֨$CS˪;�� ��]~�d�2��	F0-�Ju����qjrF*�N���qu�]˔Y��)����b��
.��i�r�0���������&��9i_	�Ƀ�J$;9�w ���:�8�Ϝ�үo�u%
4���� @�.�_��+���-[ �6�P�9�,w�I$�C�ԉ�n�)`�"P��r?U�����%����Z��\�ڑ��Q7����<���q��n�hn�}��sF	��mئ��r��] r�xm����NF/�Z���,�ԗV�z�.�K��D_�^����}�T�=�4��er� ������ B�83��B���L�"�0����v�jW1c:�����II�������x�M���FQ��W�����ȱaK��'OE�l8햿N��v�&ŋ���{X�g �����^֨F��F>;����?���}�hK�����آ�yh,��#P�O�����"x��_�[-����(Z���F�t�x�c���He
E�͕�b8��u�ɭ�����*�YW�o�S�y.����N�ʸ9&�ˑP,�H�N�y�>Q��+�����}c��W D�|z��h��!jӨ�����	�-f]�B�X����V�l��]q3���U���^�޺�ٚ�km�f��l��Q'K����=�����Ugꍽqo���$I�e�W�\U�ݐmc�����7�<� ג�2�!x-���_6ate�$uHj�]?ۧ�í�A�A�Z�*��T ���:2@��N�B���,a*
�����a�U��]w�ԯ�iS[�p	���N�:��x)�Ukw��U!`�
��椭�7I87������<��p&!(ե�G���|#M�Э\A����G������z��/i�	��|& �
��/����p"к��^�'į�,Z^�kv�Q��y^uT�����WV�S;���3|w���
֨T��o�Qq�0���`8�_�0hW�����;w�u8f��R��־�����\�ͻ�B�r�e�1�qjer��� q�<�?���x��/>R�[xK��BZ��u,QYb�,Y+��o�0�T^	!d;ٓe��P^�}�i��$�c�0��jy��<���s�s���=�޹���d2uD�y��P�[fVU �/a�rh5#�L4�zE��#0�V�p��L�az���К��!_h���U"������3|��#���
��<��s�_��:��2�n��rʳK��3�Z�C�Ip���Ӓ!rZ�ּ�st��UՄ�w�ӝH�P�;&7���[����%�U�s�~<p�Y�aq
O
]���-��	�<�_�[��m��ßj�V
Q?��q��3>���,9�iL�I��~˸��b����^�Ѵ�����n��/wiZ�{�+<��Xf���j]:�x)�����p��|�Q�q��(��a���:r��i���#vh-0���Ǡ<�:V,�ʀ�#0_7&�����*�q�]�F��r�h�&�����T�����]�u�1�<���2��7�>�{�Ԣ�c&���	w��4�J����G
u&.��M��G����ڎ�6�صZ�EN5�Ϭ�%����)���տ׻��䶴$~�l�޾��m�ꋰ�-�Q*g�<�LX��>�<��m�y��޸���e��]k~~��28��@�m�X%gZ��lp2�x�^s�G��(�ҹ��@�`^
?�?l'�#t7�o��;
~s,c��F�ZWՎ�����3��fX�D�0���������2�fB"���|�5�M���F�����;�0���5u����jaч�����@�4�[r}��a��q��Uy.�R�vˤ�F��N�Bo1wϡ��3}ˌ��}}�ã�;����hR�HE�%��ʔEig&���0�[QͿ�;�W���؉WW�S篇���[yQ�a���}�t[�sY4n�NUU�������L�_/�o�Z�m�.�p�����Ғ�ө�1�,��"���%=w�������t�e�m��V�_�܁gV�)Y�nח���������q$<g'!Ɖ��l(�>U��i��Dm�ٲg*5i6��XLM���E~"�_�E�e��TMl���s5��I<�B�w+��c���<u����V�3�:���Ū������
o{ԕR,��q��-���3��}��8�ޮ�yʪ}��nHt�\�.������#�^�W%��-�n=9 8,&�M����YP���q{`>.�g�8�S��w�ߙ�q��2��򓿰Ar�:���fN�"a�L�Ӄ=#ˋ��D	�c
� "��A?-w���}!#�&#�m)�r�j�[\�)Ύ`�!�2���h;��;M"��-�K��}Y( �H�&���7Bύ��S�V�<'*Y�M�sJ0��F��~G/����^|ǧ���3�FE��ִG��V;k�3�i������C��+#�O�g��y�-��$��
�R������4��v�Nj�{@_ψ�uR��Q)J���>߇���r���K��k��b"Y��Wޟ]�, �j�^�F
�姖�z����殸ڄ���M.��j�`{LC�@L�N�D9>��M�j�M{pK6a'��m7�9�!���E�g5�*��.ÿ́dW����Ry�P��S����_����K�'0������}���<R�"�R�ղ�\�~(�@�c�ϐ�[�Z�Y0��X��`&nmWt�7�)Dy��Qz�0R�q=����:���EL�Q�С�Ɏ
�ӕ�j�*��{��y�ܼ\�e)ߴ���W�U���j5���3������`��\]'G_�G(S��BN�����_�PQl�,;��)���Nr��n�6����:mf�}�Q"+`ݪ����M)���(�nӃ��A9D�Y�%[Mx���鉿 �o4�z��x�1}ϕ���d�:K������v}󋚛�%�%��i�b��;��rЉ=xp���½S �����$�W�0��K�)�(��q�������{�47�V��_��UYc�^��Q��}���G\���e1�c��0�&fͤ�X�s��ۀ�j3��-7�"�(:U���S��U�8~�O}�_������2�mKd�<�D��T�mu�*������ot� _كoA��'��A�ӢsE��!�S���u��[}�X��¥Ԛcjuew0��3�ja���E/����C��c����s�~���{�;�%���k�!�^��<���!Sno��)x�e�,B[���ja���۲Նɪk*n���T�X����1lenͻ%�`&��.�
�VͩpEXv�͘5��/7�}�l�%�;{�q���!e�ir��#��3�i#>�#��(Sޛ҇��W�+�X2��"j��B�,�%AH+LUp�����;��(�������"TmY,��KC+^V;uul��Ի�n���w����Շ�����r_���C��\诫Sn�}��Z��Ǎ$7�?��y��g��!�{����vg�w�󋲎`H�@��t���c.s��������:�ё���K��*i�Mۙ{+h)��]��Ԫt��T��%��Z��6'�>�6�����;WQ��:/�*�~��+Bg@�i�kԊ�{�ڤvt^,쭃������ٽO/0�04˱/9���%H���
ѷ���jҧ=���$ݩ"q)��0����=q�#�(q��f�(��0B� 2/9��Z�@TYp,z~+�E�/8ܐC�(s���NE��:��ͬ:�`�N@4�v�p]��
Ԅ�%8��m���'�G�<�j����یa��#���h��W�� �z�x��3�S㽾��w�1!A�j����$��:���K�=�D����¹���3��,񉃕N:N�}��O
�d0�;.��Ka�B�C�"[R�o��B-J��'��o@�r,��o��s�7�Ô-Q�jt��/���c3�1��s#�j�{������ ��:�`Jl�r�A6�N1s}^W�o�*��䉣/�p)��@ruڃ��<T�?t��:��w�SO{�y��l��,�ʥ�j�L�}.J��k��/�������ڔ��b=8�{�� P��z�����c�X5������ݾx@��g)��KwԿ��ӷ'�"���θ
m������G������[�|��&�5Շ�c�<o�1������d�3�׼���;��ŉR/�_+i�y�3Q��V��솒�~������`0��UmZ^S�T-#f��9e�3zG�� [�A�ڷ�G���V���*lʆ�z&L�냶�v��t��ݫ�:�6>���6�D�:��d�xF4�C6>:v�"�1Z��j���@X|-�� %�~�7��H��&f��x���Z�K���(�]F]:�򌢺��w^�Z�;��%ݪXN��٪mT��-ۣ�h��.��
�r��1��:��I�Y�c�e5���v���$kb�}y�q�Ɖ1�v�L��r��p�|�s,on������0'uo"m���@���< O1��b}�(��b��Rg�Z鸡����S
���6B��q�Mȓ�<!O8A �DqJ�kyYW5v�3���ؚ��NQV��2;�(����>�ټ9�.yX0�]��cH�s?%NT��Ek�Q��`VH�چ,2No�/X6���j��>�,z�t�z}��.n��n�^�=����PJ������[��t���IP�@b�RA�R�r�6�ڍ>��{���>�����83NO����ʅ�7@T
�4*9[z_��Ul�Rɵ"�0e�{J�[󒜳fG�<��VZ�|ɱL����C��|�g�I�x�0�plt�>����}�K�Rp�"G�Ksw��3m���~~=9\vj^7����8\�z���	��5���=�CY��롵�G�<4�=G�.7bl�I(5��4��zK�.a���LD�\��K�F��_/�,��tuE�%�)4��Yĩ�����ߢߓ�!1	�ۿ׹�x����*����k�E����`h�Vq���OF3��u�]�Qec��>Q�����Y��߷U���3��#������C��R��im����u�s�YV?>0��p�>�,�
UVWap��=lk�Ya�^�������˨0��@x��¸�bd���35V)�Kv�Yg�یT[[�����}����᫘�4�l���[���8QKM+\�0y��fЮ.Kk��E�u����߆q����=��%tY���R�2W_�sw(p�ڸS.k���M�-q1
q��!g�]��ƫ�))%����nC/�[X>�������f��Ɯ�+ه����v�/ɔ���1�ٜE�Wo@2g@�y!>�F�J��9�ܒ�(�`��ݦ���������d��ۉ
��U�q<�p#v�}�Ǿl���{C+�n^�使g��!��aE�t��-YlbKπ��J��lz"GڦF��z{�&|@�W"���C/2p��a���(��#Mk�ōX��,�z�.�TT��3��X���Ԉ�}+4V�3�56A=��5���Z����QÙ���ܷf�IM5��c�f�6���T�k��!���zG�zb��xU+�{�=�✻D5ŉ�K�6��Ά�3�>7��K��m�-�T'���.��H\Gj��Ϗ^oØ��7&jj0�����D���4?��4��X����'x�ݲKr����5�bRZ����gX'�m32hӤ��e=�a�y3#�`��N�v2Þ_@�������H�%���x�2�s9~���:U�AF�x^����G�1����(<���&�O5ٌ����=2Pm
Mp��8`�����ec䀻ǟ2���)v�d���:�ׇ4h�1��X {���kI�����ɯz�t��
����<�%�����qf}�=�G���b����v��U!��g�9����Rcvd��R����V�]W�a���t�ap��xW���^ޖ���Rۉ��K�ځ�21x���&�~mcc��W.�bì{'�3��aϰ�飋�8<�/d�1��5��Z�V�`��$jg	Y0ה6�s����*ɟ�y�,��31��b��$��m����ǟ�bE�j��q-��Why۪�̖�e R�-a���2jPmɾ�z(�O���xp v�I��7�Ῑ��[�;g��Mm��Nr�<��Z�Hus_�H��uW�t��Q�(i�u�;	�ܽ,�b}8Y�D�k�Xmk	X�8+�X�b�*���*��GgM�"��Ŀ�@"-�u��L���GrckuI���侏�{IF�+Ǵ�5�1Qc��!�Б�	(O��� ���1Ο{�)�X�;�9�J"����w�zx���-r�n��?@��w��3~O�e��2�IE"�����+���t��zq��8�����X���~�����K�&��ʮ�C��<Gu9��}v��?���8Y�K�G����+���F5�}E6�'�R�qݪ����dЃ�W%�*Z�������Sg������|���?�X���c]Ϩ(m�m��˴��%]XFG�Ȳ/�r����������S
�XN#�����K�[�����I^Ώ�>�ȼ	�X���3T�N�����J�7�u�چ�u�"�l~������К �ǥ.�1G�o�u��=H��n`g^V��Ӑ���"na��Q���Ylٷo�Tį���VNz�i�۪U-���v/�_��fs�b��ɽ�h����ó����Jq��~��ki�;�l��7n8���ߗG�}f�}&}.��?�֨�9���6��	xB�I5��GlQ��+9^.O��j����5m$w.x��v�c��o��NЄ��r2�ﰪYF_~���^�X����A�������$�S��N��Z���o��}y� }��8���b��m��'*�q�Q�\"���)�vc��� ��ӑ'�'�p+��D���I+'�K2,�x�͘�!��	��|�\tM%���D�g6[J�V�ĎGl�����+Y|�ӓ�s9D� ���g�"���E��~��1tm�$��g�dw�m�ƪNtzEԧE����+��_�b0&��ei9�!��-v�)�D]z���X3�r��E�w`6�c��5�4!_�T���.����w�Y�����7���%�I��v�B-�÷?;�R_���	���ON8�1 (�B3l�������;�Z��F��2"w^3��ud�.�"��i�k��ꫪ�~��wY��!�y��������ޜ��M�9���R~��?�I7-�n�y�w��H˓g��[1	�?7��3��3��Q)������
��3��� �/���1���c��%4<F^�}��9��C����_!HS\��������;n�-m��hi�z�Afkğ(��R<��C��ɚY�ߓE��!����� ��R�����\�f�N�M��g�\!�8�O�q����ܫ��S�nL	i!���Y��P����٠��z��Lon��������)��1���1�c�H���|��o��H�v�Ԍ�~�)�\9��<�$�!�,��96n%8�������e� �Rz�Q#��.��l�kt�E\N�������?���Cey�{O@q��Ε&�����<q�����-����a��q��=�����LU {�ko��v����{�=9�ۗ��?�YRd�N-K�T����B:)x���p��o���E��"�%	fϟ���-�t���G�Q���Ѐ*�������S����*n��F���=��c�\��~��f�+��Ζ�Yl���>J����*8�:&8�6��ot������Y������o��V(pRA��m%��W�`HN��J2��@�KU='y��i��9��;I/�~y��w��z���XF��k�u5���_�K�����W_=��{G;>� v�@����9]�cC7q��`��0���x��Q��&*ܪ������jJ��{�[����*���8/�Bf��=���-��`�\I,��Y�I|�A����M�c����V�3�Ԁ���2V���jR���Ԑ����J	��G���)y 0:�߃��:�}#�=پ������qb��]�a�t��qC�\L����uK����iX��8��z��/�[`���YeҺ����Ƭ��%��Z�M��H佧�t[���[�#��v���y���%�Ij�r��u�/M���8������������p���l��[q�~�v�{@O}\'����ճ1.��o��^q9gPE�W� 7QO֤0�Q<ǬN������L� �\!>��٤Dѥ�F����5�
�_�rv��/�uk�p���J��=�{ �annȝ�<�ȳ���?~�Pq�s�4��U�Y_��ߔ���ڠ�t�[_Y=�?������	���4��`�oF�>Q�Ŋ�I��Q��Ʒ=�o�{Ή˱�����+r���滩"���%�?:O�O���G M������7-ң�x.I�/7���\�J3M*=�dN��u1��s\ j),��Z.���N��SJ�s�z�ۭ�4#jc�U�Q9����a�|dh��+<��w`�2���S�;�6��՗~Η;O�s�}#��v�ɑu��Y��āB�o�j�&�"-������9�P��`L���r���#)N�p?���W<�{�ͲD�*9�醁��6P�V�IY��vڶ*��ǡA�3 zv�7&vT�H�S�%�.jvO�{�y��P:ac��9/�e�M���p����#��g����ob� bȂ�[�٬#��S�;O�k�BkQh��*��s[ �I��.ɓ	(���*)�A�H7'Z�_� �k����0�a��p�ף�4ˊ����@$�*���7����� `i_���ɕo��4�1��4X̓���rjH��>��9K��s�`'����f~�� ��$���G����tN���w�a'/"Ia8��S����V�!�iO��n���:�,wk*.��el�	�� �7JHhի�ʬ������e#Cb�)~�3e^`����O��ä���%qI�)��[%���R� <��~@\���u�&��`f+ň65e+�D��-͊9���e[�5���b�Uc@^��4Ǽ׈�jc�Mv��;H�����͵�J��х�^3�V����Ϩ� �K㮕{����mt�0/{/�0~Q����JvY����}u��J��� �Z�p���«�ƻ
\�jM��u�@����������H)�pK��Y��l��~X��{���٩��n������@qEBe��2_#�Q贄��/����"`;	1��nޜ��[� ��[Xi���v���ѧ �C`�����������2A���e�*����і��ٶ�Py\1�
'H�ֶ�6���� X����P��qc�->]�Ȫ��T�Ũ���r ��<.(|�M��|�s���w7��fO���=���#�	v���~�!O�qZ3!M� 2�hR�����c�E	�V���%���$�TL���h�̤u��	"�
$&c�;�$�~R��d��)v⡢{�;�Z�@����������:K2����EE��W�P�B��b������=0�km�����S�.^P��fr)}�R�&H�ʤ�����~D.��q%J�^�5���^��щE���K6ɞpqȘy�T,�-������/��T�'O�_���xs����-����\��b.�5iƙ��b\\*
�m�h������v�d}+��vZ�e�#d��䢻��
�){��L��:�-b�l��߿����Lb�D�!z�l�R~"���{�������<��{�/Y�ɶ�hR��P�{w��A�H�Cr�n)`�RW�{�eRUYS~9q���aK�O�S@��1��.�ր��Y
�hz��9�;�C���#�F�� ^3|3d��!U��pY(_�;|��sqN�\������
t�)���F��]�_��I�X��4|����Ů���Cy�.�~%h�O�Y����7:�����k5}�(�.$��� ��8�iQQyAo���`)�M~����r�(s���{Cˬ�|P%�~_(U��*k�.�9�[<�<?���7�a��;1��b/z���?
Z�Ī��{�  �k����k�ju'����ٻ!�"�5S:;	R��[�-b����������_	'��S1���.\��%�;>�`c�+�`fg-PX�����G9{0P�E����͖�Ǝ���+$�>�_����G�pe-л���g�	��{�(9���tE�UbF�
Y�?tP�jo��C���E*oG�^��1C<)�@��0�� �W2%�����dj ������E�"=2�@WA�B� �7���.��GA�wTO|�:���Y�F�5b�3��#7�A�� �Kl�66�C���\�4Qt,�����ц��#��.0x=�u�4H�/-W��^�R�5ۢ��~�z��������&qw�s�(����?�s,�we>�=ê>֤n��P�C_��Zv��u�Y��۟���v�oVt��V�};}�Պ�	����I�=�<=��.&�`,x-��m�}Ԉ_�.��}�L~Q�2�(j�tD�+\����.���52N~��?Pm���׃�d��X���Wo[EAޮ%J*r�Ow&��sV<����f���a��PWR@,"T��vtŢ��z���G?�dU�q`ͅ��U���ҵ�I'G>�JȼF�N�n����d�W&����n�xD�K�C�O��qw?)*�BI^�ɍ]
�?�g�-@�`9�v�ۍ������:Kwn���W�A<9f�1w����>g��x��H�8{;U�}X�@���E�/>���o����V�k���DU�Ug"�%K�+�}]ED���U�~W���B�j-g�Ɒ��*B�t���3�"F��8���D����կ�|? u>��R[�֐��?iq��`*Ef�V��74�-����w�C��m�\�Ĝ(@�|�W�!;��="��p�G(�*��6��]�	�����~����W,��U��P�i�Y���|���������A�6�au"�DI<��\�3t1?�����}P�,���� l�2S�F\+�`��; \��ۀ��T�EѼ����ΩL}���I�z�7(<������D���r$FP��v�&yn+$�'�D�C����f����ީ&7����b�!7)tX�^�⪘�[�(��R��9_�\6ʩ6�%\��ץ�|�i�ƈc�$ζ(TL��Y?�O�s��;���XMkD�s4m�B{B���Kޞ�v�*�Юj���S�k����f1��Wu6wbx����;6�M�G"�T��6������l~	�=�t���D��6VӴ���Tά�_N�% �ݾVRb���N+r�t�I��u�da�wvy��|x}0.w�����=z[�!���a!{��? ����BeB�	���!�B�ƫ�Z�V#��j� ?�|�� �P��$Ue=��ό©ފ���N�<6'��qϯ:��,Yʒ��b���` �<i��
����p�D}���/E�� ^�f@�?�}A-��c�����z�9l���R�f�`Vc;9�E�G�k]��p���R�J��`@��.�쬑Ju��ȁm�9.�9I=z*Q�f5�W�z�5M�I.u�ZE ���M�Q;�.�k_����kQ���U�l1�H8;�;��#�)����#�@{���f���� �9Xz���.����֘��>��3�����e�K곁�1�s�8o�sY���7�r�E+�$��_��ӯ��ѧ������z3� ����ٲ��P//��R�����<u���H����7���e�v��|B�
�޲e|t�A��y��4�K��3�$��7(��;��n{ '4�_*�x8Pùo.�V�p�w7i@D��"t���,�BW�5g���.�w|����J�׍7D���R.`g7<`��]7�rF�B�ׁ�J�-��EV�U;��h-#u\����p/þ%��ZpH���y q)��e���qk}y�GO� �u]L��߱_\ء��Yd�<n�i����
lO�2&�b�)���A4������f��W��� �w�X!��4��rY��@n�1!�AW޶E�cE\�S\��e���A�N���Sk?�J*:�]��4��%vn��z�ŷ5W� �\�z�
sݗvC����t�L|�@ L�k��L��.��o��s)j�l�%:�46��zp+d嵼�Ţ�K(o�H�L�V�z&���[�Tǉ9
xѨ*���]�ʷhji�g��"����.@u�NYR��^lK��x�xlG�vVz1.no�cI�hE��v��\dYeY;������$���y��g�(�j���tU49g���*fg����q��gQ��C�s5�����}|ڴ�]�B��l�����x��ܕ�T��CeOY;`�̊��`����Hz�շ���\��ό�Ծ�� �!�.�H����?\<O�lM3bw�d]�<����Evw��74F$pj�w`� �M;��!l#��;E�k�U��>۾��R.������J�~���X�Z�U~~Z'��BwxN�iÝJ��l����V�)�ۯ�'2��'�q���\�{:��ZQ5[����s�M�^2$�k3]W���ɋ9���𼒵Ν�9Z�''�	*��K.�#ͻk8��,��t8���D���F�m�z���ƽ89މf�u	)�}/,*7 Ҭ.�6�:g}��w��S�ή{�А�x,���f����*�B��/�w���ZZR�v>�3�:*#T�u��;xK1�"�k��M�H�wZ�i����0�⤃FoP��p#3�
��|�L���:�l��%[�Ky%�냘��e��O�i귇�O�Dht�P�/~�3l��B.��RU.��~�řk�z��f֔Tu� w����<{����>��1z�g:ŋ�x[R�<4C����b`(8s:�H�;�@������ypG��5��X�6���k�1�|��k������m35�1|�e��˯Ky�ݍ6�`w��{td6o�'�}�fB�^R��Q,~�k��6�H)��l��?����v�A��*��g�s�b78���f��Љ*�m�Vժ'�����SZ��^S��WD�ƛ+WT�`��A@ ���6��u��w�M~л��a_�jpB�Y�� �ݏe��Z�0E^��7�@#کU�ϣ��ҿ_��*����_$'һ�r��}�~��M^P�C
^���P���"���J��\�^�૓e�+��B�f!�u�ޗ�eUt�M�7N�&�@�.�s�v�уD�{�[��ocB��#Î������c�2�q�ȃJ+d|]�����9�+wb����c��� ���M������Գ���sg�Qr,~}Sе/�g�+P�w�f�8���-�V��W\���~��J������n1�;2��\Y���T�+�t=�u5{iuX�����$s�%'��e2�q����۷*%��������}[2��M�Y�ڛ-�֓���0�w'�hR���,<��1ԋ ]2G7�<������F�������}֩w'	�����z���;i�qR.+���e~q�в͸c#�f@��Z�eq��f۱�+�������B
|ܠ�{�c�U��.\j�c���Ä��\��k6nQt�k#�ً?Fn�~��o���̘��^q�}��� �'��p�^�W+���4 ���h��͝!و
XNV(Z��蓟��~{'�'��ҷ,�v�"D�+Oغ��]��-t�D_R~�q�����Ph��N^r�_��-e�J�Uڢ��r�V�f����'�z#���7�@g_5��� XhKyHQϣB�9�Q~����i^�c�b=�J<>�p3�y��>����~ex�Eb|�+�_>���p����%@��?����~Qww9��\���3�� ��Vire틑���$ε�� ��3<��Ι�k��00�}�Y�]����[��4-\�
[��j���X��
1Vo�	�_�*�9F@���4�I��p���i�x���*5��g��Y�k��蝁o���5B�j�{�`�F����j���MjGE'WH�6+:��CO�F���`�&׊v�GU��@�������@��tiJ}�~o��IoIB^��Mp��f+�C>�3��ͨ!���J�h�m���K�cǑz����3��4s�����lE�Hu�f�md <�\A'�L��D����{w^M���g��-�P�֗	�ׁͣ��Ђ��ǂ���.5!~*Ë�'պ����q}�
 �7u�`E�M^�#:�n*��G��2�m��~R`5?ЫX�(�5��X�<����c�E�.���t1�&��,�d�`���k3��6�*����P��W=?�ƍ� KrZ�ؿ�����ؒ��I�r�q��»D���J�tM�b�<�j�mp0�~>�vXΫK��8aH�m�z$UN��~�{&um�2��Cr���1O��6pj����X"��o�ޯ,~R�;e� �l� ұ+���t�⢸�Y�EE��0es�qYVHw���L�n�KT*u���pԠ�:�&@�7&u!t���$��\[��Awm��_ܺ'�Py@ɸ����� �1��f���e]��_�(kR���n���FM����y`�~͛��}����|�F���޵��2��k�,�@>I�"��B�ǂk�#F�*)�bT�A{	��M�%�t���4�(��mG�-/��Jٗ}����D�wa���W�`�Uxb* �������*8w2ݟM�{����l^����$f�933����E�z��O�I��
j� ���5[6����+'���$�x�r�����qtzkmc�?�DuCf�&F^�sO�rk�s'O����oG�i_$��|��W��v=��遅�S3�FZ�9�d1!����0�U^(�"�UA�H>eS�H���<�tQL�|$KeZ#�T��e}M��J������i�I�x�C�cQ������P��!O��J2;�VSF�ٱ��ݜ��"q�[����� ��7~���4�نϷ}�O]���)
a�q�f�{6�Q<���y�����g��S�FnI����$4�	B�[nA���Ěl?�&�2S/J$�8�]�v��v��V���p �\T1���ў�4*:�vu2����0 F� ��Tp,��[S��`6o����buG�ؔ���$(Q�+l�*���M��Tu̶�G���'���k��*�0i�`%�F��#�D�x�0�gia�噐�֗+[�1��ئ���+�4�r�%ǥ*��	���_ȫ7&�5P��J��A1*~���I3e5�D�g�����lUߊ��dWζ����$������+��7��/m����r�e�����sy�m��]/�70�69e��t�O�9c��B�R�����jچ��mZ�P�/�o���Km+O�4Z���|*&c5�w�Z(��Uږ���<~�r��fN�p���`0����U�{��v�i���c������>���_!OZ{�(
I�Z]cQ���5���-v�:�����g�W���
�a�U�{�Nw�{^��e��aMsJ�s����ӊu���c�~\s�yJ�g���&����K�2�&�zEH5):RǷH��K^�>�P�����~B}\���D� �� �����7�N��}_�oo}��$��V�+JJ���z7i;��I��j��-"x~�|-���HgbnvT-ǲ��(dK{�F��o?{)@QL��\�]�]9H��'mz�+sk8�j�%qE��Ee`���K�RڔF�5g��(mu퇹F��i�-���v�o�yq��-AF�r�3s�E��9ɪek��g�SY�,s[#�*�����l4ٺ_�$N�4�c)K��f�CF�/��"��
�6�4�W��+��(<:����u�&��I]�Ď��0k�}$=���/����C-�4�7��k�P���`8��8"E���)�@�qY/c��>�{A,?���f���4"dǼ�o�������l��G�������?`F��^�Zyum�O4ױf�'�,����~�wCUG�n�Z�K��K�~��+�YhQx���D�8#|Z����cLK�����o�K����j�]6Z�F�S�G��V�c֝Ȥ�WQ�'24Q��rKԷ$Mθ���╗�C�jS؋âق����v���cv�~+�0�}v�gE;��t9g=��is����<�)����2`�fy\����|nU<��_H��	:�\H Z(Y�$a}�!�c�0�Q-E����W�$�:��`AE�+q
�|���:*�{sb��Zxf�Rr��/\d�
���7E)��1�@���.T�Wa#3qp��&8�������E�&�%P�b}i�5����rη�N�	����h��3��>j�^�\��wB܅�S=���W$n=��1;�r�w�v���M=��e�:���Ҳ}u�Tq�_�F�_Sj��dٽ�Y �?J�'��=�1D�}��{f�z��"�������k�f��s�ר魵1�j�j�� ��P59��m�D:�3�@���q8N�w�� WA�?@��	�'0=~���މ�|ڭ)���
��v=�@Y̖����Nn�ƱꐑZ?#P\��	�jj@�'*�ݑ6�غnW���Z-D��	$�������]��݋�Cr#�T�{؃�߮�yX�y/�a~���A����)ٸ��3#����-�a'԰,�)���1�K�n��r��4Ɋ�N��@�'n���b�E�aU�������5�"&R3�H�z�yᩎ�V�soO��<��8��>W���$�q�pn�룔�����"&0J%�˱Y�����>�Qq�r�.3������nD��`��$+M�7#���"3�B�xV���HbǞU������|��_�yա>�c�@h�����_Y}�ݻ�A�]_���H���Uh*`wN��:z���롃<��}\�f|���ve������C�7&����_����EU��xCС�J�Lm���+���`�/�
��2����k6[��;�v��.���{�#��֪�h��K�Jճ�[l��u���[�2/|�9�^��/��9]�W�+@變 &&���o�ĖU�h�Cј�5����l���1j��W��A*o�'�w��T���")&]O ��bm����[_H"����b����lq�ܕ�J��@�Ow3p/l`�!'��aW�����XX����x'h������?�Y$�X��ɫ����v��%�y�z�Ԕ���D�a�e=��4wW���O�e<�]/�h�|���2ooƿiZ:>�m���pN�+c��-/V�	6
^���͵l#jA ���$�z�8")�+�i�r1Z-����
�cB�&a�6��fu�߼<ԴUO����]�KO�4';�&�,��\r��'J!*_����Ư>�ne���MV!�D�*�XH2�vo�V����a������M-G��:��.>�lH��z��o�[�X��=���c��ܧ��M��]P9_p5?m9&<�(�jv�J�҈P<���㳝oqk[/�nLte���|�k���i��f�jI��6�X�Ja�gw������͐ �ӏ+A��U��<V�Pg�XLupO~'Dc9\�k{X�2m����(Oyq�,��6�7Dbk��험 �b��~�$v�Q�)�S��+��PA$�	��Y ����&�Α�oOl��7d�_̩�f�;�I���G;n�}G�ˏk#���W��A¸���:�A�c,�`�����;! ��F��G�}}��h���A��î�Q�\�B�i���Ogf����vn���렟�t�����M��e}���F�k�}�8����ҝ�]�iAZ�{t#���������������b��8��y}o�v��wg�tj%�{�_���O��3._i�L�[���Q&��[Gz�be�MX�/3y�P�s��e����;%��7�@��fIs�,���>_h)�:ʃcĐS����>�Y��l��c��nlJ��D��� ��UYIw�̂�����L�C$�v- �ȳ��"�2e#3��4%�IwQq�� 3yX��Z��D�$g����p��.������n1o�z]ht����n����/�7&cN����Y��%q��2��9���r׶B�	e�9@��E8�(O�+��0���K����m��#�m�����l������S�X�z���q/�
�:�4�j���H|����I�Ϲǖ��̭7��E�hTr,�PZ�I�@�͆�2�q�G`��߮�[f�������:�f)(?�������P��t4]d��p0Xv�ѣ�Y�Ө]�9of,i�٣1��ʾF�/0t�^J��w+�m�1�ʬ���,����Ԫ�Ȳ��=ʕu}.�ؼ��>ڐ�t`�"%����X��X�Y+����$2,�2�`O�thN���-Y�,o-���_�	8����l3]���*��CQ�%L��H::����ͥ}Y�Շ����	|'�����kq��C�pW��s�����eJ���o�@0"	�g�cɫ����._L҃3���}��,,,�����v���R�g�\���=�zL��5ɲIΥ���gW˒�VR<S�g�Օ{��o�s.�b��<M)F���e$̭�c�hЫC	��u1�<N�0�G��!�M����N>�i8i0[ϨG��j),^9)L֙����^`���Ե
'ݏ�F�C9��mKf�i����B�/�[�;f��_�hC3c2�.��tC��ǝ�4�3������0�\[�ˍ�/O}��e�����;�.��Z^�v�u����4��G�AY��n�7-l��=c�n�T�Dc6�w�Xߋ�~���@���m��@��$r�|��>*�Q�2u��ҳ���(�9�#�?��-g�I�z�C�2b�C�~91��-��k��n]{�x������{9lT�Ջ�ϐ���r���Hð6QS��g'�����ٺ�>��U/�$�;�J�!�ɘ��}󄞫�{9��w���p�<7��-���a��!��R���Jd��I�a����<e� �AK��!�R�y��k��e��#�Ͼ��sT��u�p�	�=�iz�:�#�s̸k��&)R9�^}c�J������;XyX��;��Wa�#͸U�V�u+z��G����| �3�j$_B��Ջ�@�:,v��X��Q/��@��Eފ��L��)Ί^��RF3�U�����Og����lg�'R��j�A�mj*×y��S�d���@�:�^=�'�ٷ1V�⒕a���E�����ҍ��;.[���������7'խ]��;N�ۚ�<*F�p~�}YHd���u�@:--g��;���������扆�i��Z)��#;��{?����>�%��4����<L ?�di�ޭ�	؁ڌԧ	�����U�Q�^}~6�'���{ڜ��	|����y�d��A�f�6+�\O&n���ܾ�:��p�}[=ֽy��b-�&9�Q�0ǅ�>+^g�6��\�yy	S�XB�����nN~S/*���D���O����ox���q� ��^�*��Oٽ=Is�M�>��4����.]x��]��YRY��I*=M��G������z�\�e&K?u���
�/^[W�n����b�k}군�*���R�c���NI��&o����C�וY��к8���a�� ^ן�C�$��c��`ħ��$�ٚ����.1L�v ��c��^���:�����lh��m����̛�^��Jǅ8) *��ᒅ����^�|�]�{!�v;·��Ƙ�?��g�����%'h���v�A��� ��	}9L�hu�@#�ƿ٤���>��f�\����w6�n�F_!���	�Sܸ'��<TǮ���Dߣ�׉�rp�қ����^���ޡڴӌ�#>����u�I�D��~������S֎����N6����jl !يB��e�-��{��럃v�I�C$*�����
�m}T��Q�ә~����MEsɔ�;zn������٤Aw�âe�ңu�1r�C'������}�XƇ~�yvGx'��w~�%�Ҵ��8�V�;�|��CGq�c�x��2���/��`�׋��{i�p9��Źn��W�t����N,�k�#�}�R�=i�o�R��p�7��̖��k����m�-��5q��ҭO ��;���{s�ýF|(���洭N-�����l�_���!��
���e�W����N�`�v��X6���G24�6]3�R%UP�
�3�O|k�*4wWP�H��C��4`7��$����OX71	���z��.I����uw媵��W�	�����"L5sn���H:>HNZ;��.Y[��:s��NJw����v��f"����߯ŵ��������׫�>���� 4�~[��;Deo���>�Ʒ$tAHȢ�E�[���W]r�� ݀.���Js9mfˬ#��
)f��HoD�57Hgz�� ���o��D��g��z�*�H ������6|	�x��
=�U�K���olQNq��Yϥe���b����̄���7����Q�'-IE�f��_���Q�Ѽ����ϛ���Q��ዞ�wS�~�{���Պ�u=�=R�<�چ��og�B�@_g�"Ӧ:�u.*dg?ŝ<d[s�d V�E��J8nx�4�,aoڿ�z;�Ǥ!<J�'��A۽�0��n���
��$5�Ook��1��&Һ��<O(Z���Yt�i}�5H���t����-OV^�w\|ymF�a�e��4&�F�~�v���| iV�8*�Le�*�v�5<X�V���-`b�͓u�����Kp��E�l�v/��CQ�ٮ��L���L�}|smB90IS:�x��$�ɑo�y$lwU���^��&j�q�$|ȃ�f�N{�L�uJ��ޱ(�3ˀe�$�ck�&ˑ�ٖδqh^�"d$|��4,Lm�#��b�wJ������p+~�.
>~���d�?�Ŵպ���A�S	��#4�r\�3�ZNA�|=q;��&��h��{�]{C��i\|���ݐ}%�αx
���n���lC�0֊��e�س�����T���H�,��
1�Y����e�c�گ#��u,_W�67����'��@����+����-��%^��eF?�*C@��ɪF�3��*T�.��φ٦v3�[�?p�[њ�Æ����^��2gDG�.��c$X,�ƅ��:5�k仇޹l��{�%�3���i�>8�$�����Dv��B���VJPh�'�S(���*xJPϖ�k��I����h��|�OV�"��L2ۊv�*�M{�4��7A`W���5��k@H`>}486�D���M�	�GIJm��~"k�u6����a���ay��?)�����
2�pg~��>�?p���,v�-$��2>y�MBA����R`z�P�q�h^�/.����<)������|^qxr�y����drR��i���f(�~/x�V?%��=�W*��:VL��@����N�d8A���L#��χr)�pyvM`��o.�rf�0�������Ҕ f�����H���$��+�"T=��.,�Zd���k)�%J�Ǖ
�B�(�ӪPO-�\n̏����CRs8�_ɟ��2�?n7�&�Y�Vm-��ϣ2V��(h��P�
s�<�����}{��%o��(�%��'V��Se���d��@�����8���*U(	�c%�^z�ya��2�^Y> �j�u�jѧ�$����ruF�5�������<Z"U��,[~���o0�1ʪl<�?�e>��8�m�NO+��R<~�d^�I���~�����^=��Sȯ�� �s�]oSU��Տ�q^�m��(!� 8sNN�e���ܜB���ܳ���S
��c-a'wF	���+���<0��ZE*O�z,���8�-�0u���f3C�*;x_��'�8��WQ�z�����U�i7oqv�[��,�է�{L�ܡ���DrH�#?&���Ա����D�u�!�,3�r̳�"!�SkF$�g��"E�DV0je���]T�_ĐX�
~�ڢxd��6U���HIg�O����G*5O*'	-���gl�Eth ^�K�����
�g���8 �˖�5|�"]��9�p��X�[�H���L�n�-[�:�+�ӷ�^�_rC��F5� ���^��G7�W,8�63��MBY5�7S�<�Q�A*��TO(Գ%by����粭v�'�a+���>ߏ}�}����ɳ
N#A�O�Y��'g��#!m�%
ܑ���`�TB� f���^�4�W�_�O���2���ZIe�2�[?�����'�(�DX�!��G�k�8;wda������]u[�_Zb����̤D�:��X(�Q�kcQhS�~����3���O0��pwDXٲ�[ ���{b�G	�6�3 9b�e�#�������ݯeM�ۼM�K �O���x�D@��J�B���J@��dm��C�X����Yƌ�O��~�ڽ��+�u���0 '�1�U���{s�SA�����n��;���>?�L0�%������Is�$t�˾Ok�� �ڮ�*$Z'�?���ݮ���.����l��P�T�͓\�Y������W,�Pc.w8���*Ux~��ڱ��dd�Rd8�_�=��P�-#����WP��H��G�ث�y���L6�!��de��|8���9���G�����:^w)�\�?,L���kV� ���PQ>�c���>d�	eu���}[ZB=͛�]}��֭
��M�	"�<mXB �����O�f u{���
��6�[衮U�7�n��/d����	��*�8����Y�)nw��)ۀ�ٝϵ�>+��~��߰v�a�|ʞ���������"����|�ha�S���?\���}��~�<zٗd��{s>�U^�E��3�s ����,{�#_\8��dk]go܄��a����3#���e�a�<�����}�d��Ϭt�	�P����0�W��.�qe*��.�J��Z�ˆ�枣�i���	�����M}3�@����B�48���{S�vl�.�
Kov��-�':��蜁����"�8���zv+h�6-4@�߰����1:_ŀ�
�nqü�f �}V:�q���]r��:�쁒P Ժ��Y3?�]@��ӵA>5�mm����]+��W��!����|��W�n�ܔ7����#PK:6Q��/B^��kz����S	,3�f����T��l���i��="[��-��4�:L&�rb;��$ᜢE\V�n�'��/�0�!�r	��ob�zÓ����g}���/��Q�Q�RcovWG����a����@�Up[=Zê��
��u�A�i��6�X�C��x{?i�$�D�s���,u���6�huZ�
9�����5Ϗ	ӑ�E|��چ1~g�st�ˆ���!����a/���������L�/���.	R�E��*ݒ^Rd=Ѽ~�ghma����,91t;��\�>N~�n�YA���&il�,n�v���R��ϿnT�w�Y<�/�������?6��5��S�d���"��1���4�I�8�S�E-�p�SyT���H�Z��W���(��ۙ,��7כ�֙��.��:N��kC��C�p�'2M�T"�}ԁ�"e5�]�;&�MiB��.o��I9饽�,���&m;�g]G�t{C8����[w}$^�k���侰z�(�������X�`�C��`��j�ʏ ��O��VJ6�@s���M6i�3�5��"z�=���9�e�Z�P���r���P��]�+׊>z���c=P쏛��c�})u�������C&5R�ڼV�PQ�N�����3ԉ����6����G2(�l&�s���������[�l���w��2�[��H+؄�A�U��]���;+vU��)bGy�����ޜ���:���� ��4�ä>�u?ڞ����-���:����ޫ�k{퉺W	W����{�.�ϓQ�U�>�D�à�Qq�j����g��nx_��ci�ݙ�I?���`���pF� �������犓U�19U�Zӽ�uJz����[H�u���3���N�88���!&�ůr�p���d Xz��!m�j�p�]���r�|~sSwvX3�x���
n�tJ�跖��x�t�82�=zE|�%(�@�O��d����WoR}�K�݀�������A-ϔ���$R��9T�z�B�rG�0_j'�pa"�倉�7ȹD�@XO��.K�5�����~�pTAj�'�_�s�~��A�}Y� mh_�/Ɍ6 �=h�b%	Ɇk���E��q'�il�}T"Y�p{�k��t����;m�>M�z�'�-�Z&�f?u';<�M+���<1�q�����
��4���q�m���i��WK����B
�l�ԑe1�w(@jZ���9���ξ9�\2���\�FN?��
܊������?��`�A	�i��ځ����,���Uu�Oy��ql����)Y4�wK����=��^E:�1�>P����x8?ZX5�^���4��W8�U��4�ډ���H�$?�&���S�����9`�ON��=�p�݊ ��ޭ��`�����콩��������Z<��&2�g7_
^7�ߕ�>��"�^t`�x/e?��t�q���� �x".*y�C{�Z퍪KpB�Ex�C0��F��3|pz��R�=T$��uvZ�U�������} w�ҟ�����0�u��a��~��<��]�A�9��{���Yk���V����A��*#���%lʤ���B���6�]�!�:-�X �̇t�&P������~��#T�r��$x;�D��	��5������n'￿�&��V���$D��	CMp����b�`����^Ӣva2w�]P%�S�wQ�|A�&A^h�V-�M^ ��B������?���qLҕoV�������)�c�*��������D�g��n��l�0I�0�$�����E���tA��7o�n's��j7Og��A�Uo�&I�Z&�o�Ӕ��%� �e>q^����wr�m��c��/k#ݨ�5Je��٣�'|-A���
��60��` ��|�b�H''�9�|T���n��σ�/xCV�%�({�����\���-Ҫ�T5DՇ��ն�'�f�������=��a�L��?��RU-P�*r��n�+4�zQ:�M���x�>�>�����D�aI�ߗ���N�O��㾆��?�7�:-�9�::�L\��p�7�ֺ����X�u?b����p��O/;y$gkW=Y�K���#���"G[x0~,
�<����S}y ʬ��Ϥ��+_w��8f��2�L��AKj�9��<�B|v`�P�n���.y%pCT5�O<NS}��@�|!ǘf�z��G��G-:��la�?Z���r:�9z���!��4F�벬=u7˴���gemOX�8ǧ��בM�=�z�Z���=Aϣ%{�J֮�Q?43��Z�eF�`���mE��D�R9���[�p�6�q�b9�7��ma[��o�ǚ�׈q�ű(�]1���C�8.��/�u�d�
0��S�����͗����x��x�Z�����<um��w�����Ȭ�-�C3=Mi��cW�Wp�8�CF�Ҝ��[��φ:�����_\dTV��?-;}��{@�������0%㝦hɲ�[2 ��#��6��=�C���X4���^N1�pc=]���>
�C�����{�6�k�8�vI�5O,�1S�B�~��0�#�5�F�Fg]M���R�{�h�8K��H���ГӶW�c�7ڷ�����߮��2��3�D���l���3ƌ�bn��ܟv���aܽ�����a����`�z��dE�x����U
ɽ����1��u^��mo���"��܏��-���9C�ij��(��-�"�K=�ҽ���y�R5N_(vvi�*��j¯uA�k��h[{_�g���J�w�g���>B>'���N:��`�*�zR�D��4m�[w��¦߬����<\�eެ��rst����?"�������1��o�_�K�DT�4��a}h�`H�O��6���Nf��u �%�ߕܵ(����f�	���J��L�q�nzq?Bu����uڻT�6~���{D8�#۽�&��%^&��p�VX��<8��0IcN�Cc��B7��Kk������2�lr� C'ym.k�(S�B�%����E�Ԗ��l��h��R٤��ș��p�u�]�n��<��<j�ҊU�N{�^-�5T���Ź*�P���w�]G�������z�7�5;�~��sia{Q'_U��~q\y1����K�-��2���D�o�p�?������n]-����W1��@RX�wS��1ɀ�T��x�f\D8��.s�&$߬ )��ȓ��.k�aK֩�hё{n����h��bN���oMr܇���,�,�XNCT�p_�k}����Uɬʡ�k�̊��L"�ח�>�i�4f�����l����<[���e��w)�+|��s6#/Uq���V:������%���83~f%,[Q��R<��ې�&	9��T�Ƣ�%] L9�秌VMU�.P���>��,�Ζ��d�WC5G�7�Zţ
mli�waM"E�m��8˹8���'yf7g��6ZP Gxt�z?�ְ��y�2O��kko�io��4 f�}S�V81A��^�����:��4���yP�|�HA4^�����'n����7H[�E���O�Qju�Qg�r��齱;^��z��˞ɷXj"z|zq|w�I�V��z��CB~�節�;+I��96�b��J#����q�F&��eY�q��h���}�'4g�2����礣<7H㫳~UI�+~�*��m�쎗iq{h��)��Gn
��]"�!����Ԧy�o<��ӕ�ۣO4\&3_�
�VE����*�����>2ߢ����.����0Re�@�y��F��ۑ❭��ܣ�s��\��76Hk����¨j�P�6,s�h1�3{(\�n6�v^�k��}��A杓|"�"��]�AI�	���l͗^ͼP���M��C���p"-]�D����F�)%��8B6��!�%��]Ϝ��8����E�;���j�m�2MI�/���{��,��B�Ƙ�&��)�(�^ΚK^^Y��_�#,us{|�]4�|��)U<� �Kj~%��IF��4�t [��2��VE���(��Yv��~�|��u�I-ipr��ԧ�w6�Y#�[qbfjyr�����в�+*�#*QǢߺn�\t!ץ��u��/��W`!�l�n?�ʬ�GÁ�����k����ZuA�ʳ��@Ȟ�k��K�\F�ڐ�|d{�Ⱦ��3|P�2Z��YqP=#SZ��Gg�{�����_��҄JB+����=�n8靧V�5�v��Lu9󖿑���� ���!���gWw�l��abPS*����k����_2�6���Tg��Ɛ��q��̱�J�ş�Uݓ�{�h��Mx7��4΋{i�fFz�ǚ�1lh�S3��Y��e�A���=U�E-��Y�����
Sj��;��0�cCǷ��kD��<UB���{{W�\���Z��;�I��r}P�grʊV���8�k��6N���wי���\��׋��wf�����\~dK�]�5V����|�_�G:NW��B{��?��6��d��ڊ�.�槚�Q�������v�䈪�s���B�O ��gz�'���*=}կ�!���m��8?;D�7<��>�']!�����U?5.OQR`��>�_L�>3�R����
.�o񘑘�=B�WE/�x�:���v���7^�<�M�����@�u�-B:��K����A^��ff���, mx~��ۿ�x��������C������
�o�# �e����K
؂�%c_�Y1�+3w�	��B�&go�J�gLo�6)�`gC������a'b���x�E{�?]5��3�Y�QRp�����J������a0r�����xPpyg��dsy�.G�^�?�F˅��S�?� ��|ZN����z���U4�p���F���'����o[)�����p� �l��j�;�+���P	�q��+p����߇I(Ar��%0��YH�mQÌ��T��ΨㆸΨ�o����;���Q�� ����r2 `�r�c�����q����P�K�s�I����V�ݘ�|��;o�kh��K�9��x��񰯦���s�_现���n�C�DO���B���ԟ�^S!O�n�N̰ho�O��6�I����h�\f�;,Gw����B���>�.���2_6��UHӬ��.ֹ���Omi�����̾`z�ed�8)��]�l;s��Q���3 �.(�����]z�:��@ݝ�������
�q"���[Z���fo,����/��.E.z�=ˁw�7��S�7���-����j�����DQ��1���iIkW�L�4�P�sp�5˩��"/��Uv����o��\�99��,�������i��FK�Wx#�9�AGVV.(W/�+7ڻ��l%T�	�(��NBL�C��xЋ�j��yL\�p[Uj��.F!��?��jʢi�^�#��*�$� v����'ۛYN�VF���~����4Btx/v��J��������r'�d3�طb���e�dK%��Cw��Y��2�<LNY��b3�4��֒U���S�*��g�-,�Fi@#��l��%����JԷ�_��Uգ���)�d�wr*�5�5I.*�p-ӓ��Ǭ��Σ	��R�]�I]?���MW�ؗ�,�ɬc
C7c�����&�	X���l�u��k��6��|<{�^��d"RItf�-�X;i����'��'6���G{xꊲ��p����"�[�����N,�� �]���O��
��q�z~�ÜN'o�/5ԩ���Ǘ��P�%�{��/���X�b�T><�/�~��=s �5�c!�B�O�L��f�aS������`+x���vf�<��[98������GW���6Nm$�.�-<�Pe�V485�W�o��(�<?=w�|�h߱��œ,�c?����|2;fｋ!��)F�A�N����	u�O�j��A����'Qi��i1�ߦ�%�v���A��"?�	`�JOx��ҏbQ���g���2�"�u�f'�m*���2�)k���6f�H�/܉@����ԛ�ܻ�ʌ
K޺���S?~b��n��f���;4�H��o%/��*���k�QT��/u���v3���p����r]�a9�1�cB�]���zu��	ޫIF�©#2�(���R���r�)Ԗͷ��:��}��cy���Y�)q(+��+��Y���[dȴ%�,Z�~���u���[���R4
D�xy�+�|���?��f��Ĥ���/Q4�i�=z|�7��*/���.���ug��Z6��CЃUM�xݟ��oA_R�u������M�� 2�mW�z�,
��k��5�1��?�����J�n���ڂ�W{�k�ž��}/�n�']Ԣ9���۵�l�p�*����#C!_�qoiw���TpB0�)�ٹѫ$�s>�#7e�}�ڷ�f���$��������W8l70��e)�ß~|��1��N�����$G�ܽ���+Tk!3�!~����'{��"n�,!�W���h�<���ސ,��M�@o���0���:�j��&7! �$R�ke�ͽ�@���!�H��r�ݿ���h�-_��-�j�)pվ�*F֊p�F�`u�v�$?��m[��~ٜE�RB;N�D#�F�@�;���i[�Jӽ��5��oG��ĞykV�L�����|A|�}�7��fb<�o��vG
Gڨ}E�0uY��C�88��jCHO3���ſg�a���}[�����n����۲�SɎ16g[���$˅�;c�y��0��Y��X�GDkA�\Y4�Z�Y����B�W;���*��Q'*�F�w��=�ϔͯ�5�O�p�4lF%�b�e~���T�H����8c�䎲R��܉����^3�����^vk>������;;�x����+iOa�f.|t�H����S��ytˇn��E	�����M����Ux>H|(�O�P&w�0xW7��Aȯ%���akm%��:��ʻ�0��7���5ot��(ܥ�����R��Z�/5�̄�^��A{R�F���d���t�$h�i������ݜ���p��k�56�n����~��Z:ߋr�%�S�m��ClO�w����N()h�#7p�V�4Dk���/�Q��C� )��_��ـ�����b�\�E���l 鏙dDA�E��J�<�*�5���C��;
�"��2��¢Oq�K�{��3{�X�y�.P���������~L��*�E%��Pi�o?����h8��u)~�b6z����,M��]�Ÿy��흙�H�7 vEV��6��uE9��y�.��=�9"A+�}R�<P���ď�sSqy�����X*=K�������ɺmP�:���o��s���s��0_RIf������^�d'�}I�8M��Ne9L�T�k-"�;Aɲ:��d��W�|8j`P�S%Σ�	�qK����/��bv�A��
�J➣�d򑿍�)��*fU E�&��Jn,:��-Ol����=
��mgx5���ě�4iȲ�JC��?6�wΚ�c��k+�D_�g�t�����n�&�-o
ͻ+�����w�2d�0�aà�c�Oܮ���F�U�o_���?C�����:�Ӝ[�;)P!�W`���u���� �I�`u4_�ڰ�t�l�ȯ��6��<�R� B3�h����!����U� �x�?1��qȭ;:�Tн�IV��Ԝ����['�����tU��?���becs�0_���{��Wf8��'o�LB�7W���?T�)�is��'��v����xB��شxu�-��]��S��Β�W�`�b{w��	��Wx���^p�4�4��$��2b�ܱt�l7S%� ��+B���N٥���ȡc/�A)�Ydc�,��"����q�ç"���&��X��M��̚��a�m�;IWK�ixO��&-��8�ϊ�DD���P���m:`�3��ғ�t��@[7\4�a���B��O"=N="�D��Em��r���F�m�ڱ���+�R�t���4�ԓ
�@�N�ܮ'�=y�������?D���hv����w���*^��l��BQ��ְ����s��F��%�x�eX�R�lڇB5L���g��n�jF2���:�2LFKyJ����7m1n��
w�k�D�8�DȾ�5|�z屹����?#���]8��(�#U�9/���K�R��bY(n�����Ter�9Q&Xn����pk�lk����bHd�C�}8��c�mrvk�l�0dL�&���ʗ�:��i��?�{m2�G�F/F���z?��gƱ��-l��ݥ����~{?��7U��D��W��꼮6���)�$��&�)�����Vq�.����3.�K�k�̩%$R����J���x ?Ie��\������~l��$%�&�R'��l�9[�L�6&�� ҃�Q��{bl��X��X&�i���#k2��e";2	xzl�8����֩j4U�@��(Z�����4tnA�M���[u,�ŋ}���9�^G$Jː�kϪ����{�� �:�6�����qvś���7!�c��{���[!�G��}�	�O�������n�_TA?� ��w���?�?%%�ރN��M��2��	t�i���	����f�vX�����W0x#y�O�u:T3�ۙP�
U��\_����l$���#���x���i��ka��iQ�p�&������O�'v��I�Wn��"5�|ӿ���tȫ���M����o��U@?��jݷJו��[]�H�P�U$`.�m�lB�#��f�be2�}���z^ ;������&��\*�][�ъ�ֽ�zi��Oֺ+27�N��C���A�W����c��Zbd"�ȭ����n~"S��[R̽o�!8�b�\�� �	��j��P�~E9v��54)�ciy�a�*+���+N�k�˓sߝ+>��K�����l��t^K�h\{7���/-Yl�G��0Q�����D&zj�.I&�|Ȍ��&_s��ݞ��4 ޴��
_h��,�����}V(r�ڔ[�>`��蔆���A>zk���0n�_(�ْ�m�Q�q{���Eof��g�t�Ը����oe̓�>��UAC^�27�҂Ŧ�oȰ�h�|�{f[�H�=yx�j[[TkY�=�-�X˗�IR��ѫ�Y�[T]#<�"��>��H������W�� ���\{j���kΈ-��c1 �SX����+\��FE̜�ǻ�~=���t
L/�w�gaW�v�Ce4��A�S����W�������3=e���ˇ����y���Q�8�W��/��P���'��c Q�lQ�o�D���ψ`x��_�!�@jWC�W�y���Aщ�g�<#Ҹ�t"VW7Z�	�΁��蠖�����2Z���H��H�Cw��Mo��f�n^R]A����v�����.��F@��fU�~ٚ�,��V���`��������rV�ԑ  �{�'��i�\���W�!-<���0�O��v*�����g1�kIɆ ��� 4UȖ��u�~�5fL��y��i�2��p��{J��פ���������hH��0�2c��[el]�b�x.Ư_N~>-pP��ƕ����[N�Y���"��-�*�VC�O:b�^'E6�7���9�J��*�z������`;��5v�Mgj�����lk�2<-%����i�Or�������Wg�M�r�����"�B����H���i �Nh�����!V���	㴆8̐���⌤�־�G59�JK�3���;�4�2jc���YÐr��2���R��n�����R%���E�Ǒ9�X���aYd��b�?�`A��^��0[�ǈ�a�6.I���eGѫ�M���5��W"�&�Y7�ήl��K��A�]���E2��2d�Y����3ZI#oPE�F`���#x�%�Խ!���E��4�V/�Tfބ�G�a��٥���m�p�S�h)�Im#Cz�2�C�*�"�M}A!����;�Q��o�8��޶0�(��+��>�l�Oئ4h��ʻ�� [)i\[:'���m�l�u�xQ�����#bqBS&qq�پ�W�u}��
/_\A.��_մ!M�bn|��f�����u���~���ĲT�I�������7��Q�}�v)3*K�&�5�ކ|��;���X)��k�-����3���m0�d,�uW٫0�)���!��hF���c͋����v"�>��P�v�GN��dq�6� �5xCr�7T�,k�HD�b����3������I�^k�����DztA��.���C��^>��V����:�(&�f��o��q��{��A���g�a�/M9K���|�"Y�#"���`�� �����Ozy�GZ�޿=!�����)|�X�1��2<
�_۪�EV�<s�������i#�� R����t�|��0o���s�0#�=�b
�{��E�s��6f�aa�9��l�-���:U�1��,jZ�à��������뚍7d1?������^f�'��_�G�C�_}�.{�Н�_M#I�8����]q�ՓYI8�r	(�č#Bn�*Eq�s�Zhn&���њE��-��t˕�D���e���vv�Nyh�?U������Sd���[;cΉν�zI�>~;I��M֛f����V?�'��Ui��7=�&��V��3d�N���]W�?��� Fǎ����Ѱ��Owc
���0�_j�?]%��b��2�ц��(-+�Mb���m���m������zH��ӓ�X6t�~rA���*���5�����LLĥ�_��}E#S���Q�l���`��8bS�H;`�j�[A<e�ZsP��8�W� <M�s�-�^�r�7;?�k,�A�pp����.F��R&��H[Ӭ�vk:n�Ʉ�}1��G�v=D�*�]��)G�Kn���(&>7��o�2A����'����CpXn~V�q{Wf#HX	ޡ����K.6+	�P�X��Jeބ�K�a.PZ�$�܂/ki��AIa��&�ݣ�!��4�[\M���%�;'�����3��4���C�dpw���·�����]u�=��W��Æ�#��A�>sq~�5��o�+��j�xkL�cA�a词�4��A�Y����:�3l(2E��@���{"J�#Ah�i�:0�S?��H���� L!Y��:�F�U|��pG���Va�eJQ�'7��7�������7Z��S�e)�_Ң����f��Y/,�Dѻ�I�V�=~�%TɸV	�������3����R���C�[��"$�ٌ6�v�X�@��ݟ�ek�##�gZ��.���q�5������ ���*���_�)�>Yǐ��C�.�#m��n��!"�9���ə�fA�������e�#�Kz�K��N S�0�XD�U�#���Q߆�UT>}�m��*��t��q3ej��K^d��IM>��Z�b�z|�h{��:"칡�u?�p�x�G&���}�k�G�{�v�!eE`
dJLȎ1�g�RT̀Z�,��)3�3*h�Ei��u=�=�M�~o�;̮�V̇�X��-�P=n�"j�d���n�G�i*�σ��;W
eeU�������Tg��K���YF#~����Cb�ŷ�@�!�FC��o��d�?\'M��ۉ�;N�!r�&!���&�<Z�v���B}�#
�9��@�H��\��ձ@�S��WRD���<���]�����K쓾�X��KԌ���3��k��n:���S1��O?�����s���3����F���5&QU�=���l�O�(Ȏe,Fm�ҡT�c����^�c��i(��6P��`<�P:�����( cĴ4�*�ʓ�灨X\��̑�{�Ҳ�'W��$&����:Fk������D"���Tۼ�w�Hr��Y���Sf����
d����}sbB+HT���*8ʩ����{�Z���U� ���wŗ���I]�p]��+������d�4������XQd~��:@�K˩m��?�8�%j3����þ���uB�V����g�}���37m��'�4{hD��/���ξ��'%GF]�������O����G�hH�v[���G������ea�b���tCR���:�N���)��_�L@S�H��y��Ǐ+>�P޻�(_0������w�u����娴���q�1��Y��@�3�²�A�V�C�7/�X=��c?���D�.T~wF�$K�Z�w#���x��t=���`�G�h�k�#�i������ 6w:\N����w�)!X�^��
p�	�M���I��eڎ��{��p9IMg���֬A��@c���k�=[h|޾^�4��8�Y�#q�9.��
�%��!�1�V��������M���b�ߛ
n����U�Uydw�u�� ��ʷ��t���;ΉJ�m"�M6��i�G�����FW>�w~�c����ϰ얊���<���is�h�P�Ǥ��9�ٽ�����E�� L�4.�en
�ԧ�7�������
d��>)p\x�k�6�B�=u-�Y:�-�Ur���yW���̬>oϥ�BV���*DE��zy��B�
�Di]��U �`���%o�Fg�L���kL)%Li�����������2�����>E��A�bT&�Z��KA��%�Bwd�r_e<%j$ƀ+����ί�h>�=ّH?g�o���Yˍ�_��[����x�!���e��R?��h�E{9��.�P��jY̥��.��-���n�r�I栊R���Pk(9F�w|��-@h��Gb����|8�{=��Ю#�b���ڼc�#%]��))�� ��Qp,�K��m^<au������[�C�_G�����jr��zm5�����l������X�f�ey�>F�GRMj$�n|�q�H�B�m^����S����ju^��`$2j�[U��Y�~���v�����zB$�"|$+���� "�{���FCA���#��l�����,܎��X�l�6%�y�7��3\lܩ�~�)���G+�-�x�;���g^
�A�-�h!�F��[��0'��/��覽��,���Q/�T�w����ug��<X�󎼲Fe����]Mtd"AE��>8l���[��-�+)�h�]S[r� &T\��u�,��L�Iw'�ʲ���#f����O�P5ٮ�2G���3���C�,2��j���J�����n c^4�o�ї��d��e� �|KIֽp}e�gX�K�L�״N<D�
;�h0�zc��l�H��2��QpԾ�0��|g��}oN-��+\���}?�qQ������(cBBU�?6���n��8m>y�}��&�������C%�.o�Za�Q,��o\��-�e��Ә*���t.��͡RJ6���DEjL�KS��+���5s��.V�'��P��_���|[���<>�F�?��.�	������[��g��t�%�z�>vK#�8��}>l+�2>�	J��S�kP���F�G�kˍى�\؄�	m�;&{l1���o���^M
78_6g�Z���z~ �;����֥����f���kF�O�FZ	G�!H�m�@&�)����cN��Z"�4�^��05�q�����2b�����翲/�`����޸/P���ǻ?b��̚��:6/����N���^Q9�S�Ch_�<v��ID�t����w�x��JK��)N+�9 Yr���B��o;!DHb	�����r�=F̂c�,ʆ�T��7�%^HpphM<�����Cm@D��8���.�?4�q��ff/�m��ib��Sc�'ڒ|�
��Qew���xj /o[�/�A�>����S��m��R��.�xx�a�#Z!Nn�!�N�58���6�lU%����C0��-���X���%I84.�LY�v\ޞnѩ�;X� ��.��h�
���u�B�ڦ�;���<b7RM:���Ȭ�+o���t�`Yr�U��3y=�{�������S�!v6�N<��_X�����j��,l2D����X�5#�Ȭrz�w}#x@�;'�k���#�7�/>������G�����\3�n�fy���b��.�i)� ߐ[� O��/��ꚗy����e5�uU��Y�Z�Z�.��U)�@4e�eA���LT���!�[���<��v�	f���B֨�`R���F�;�D+b��f�nD������Ğl>oV�������L�&�/�����v��86׭&AL�b� �asdb�L,uɲ�4�z��8*GH/���f.���n�T>��DN:��$���uV�V��W�$K@�� ��<d^G׈6��3�x&(�X:a9��ܒ�t�������Z����*Pޝ������n�;u!x��9~�d/s]���O���E�5�c[�{��A엔O��h��V���ׄ[�l�Qܕ�id
ޥ/l�H���2~��f�H�<g�b�< -
�!h�rO(0.�+cP�(\�ź�w�i���[�����6/J{H{�dk�4�j�܋ۯ�<j���X�<��������k�D��%
�1s�p�L:��YN-!7s�+�o�hiÁ�J+ ��<d�)����ްI6�q�Η	�����?�lg�d��Z�Y�7�E~̝n�߸��kXm}e1�i��K�'�m��|�n�N0���ݮ��\O�帖�Hn�~��\�A_�&�+��N�����!h\��%���Gg�T�l��jx�7=�e��a���@�jdI��j�pD+��Q(�%	E��#u춣 �
�H�H�Cn&����TM8�H���c��-?@�e�{mٍ=��p»Z�Ɣe�B�Mb}!�����c-�>��%؞	:y.�l�u�U��}�a�Z;H��c:�&/�*��;�S�/!���`�NAifb�,,6]�"hq/p���� �L�A��Xÿd���}ƕ,A�%n7C�*$������I�<���͡eTޭ�Z!�t#���y:�ƞ�y���FZ8;~�q�h#�:�\�FE����<���:5Z%�RIO��܁%�sWK��.��]]ś\��Y���\k���z�:,�U#�N{��!E5	�.14� a���p�Yi���|I��lx�m��6�� R�����]�`'3+��侷�����y�����UN�`[)K�Arnl��,I6��d�mq����KN�☠�����y�3>m϶N�;J�7�	b1��pv�|K#t/��4|�`��#���}RG�94j�boO��LM]@`�Hrw�{��%?�����J����!��K��uJ���[���*iL�7�3�/�F�8�-Y�_sP��Y���KӴb�3a���=�<;��Q&r����䩳�5d�&�����#j��c��8	�72��˭�=��]^?�ݎGԳ�;%ѽ��bh���8u��E��!��}Ys
�8_�3ٓ���h��#F��N�+���"�'�6���h�K��k3����(�8��T�)&�y7J
�Ilx�ԶR�5Gu1��e���~ɭ��$
}�÷(�)2f�`Y�٫E��#4�}C�u�K�KD�Ma�O���ְ,�<�K�:Y�l�m�$�6"��0#�N�"�'I@�j���U26hZ��'�}CSt�1�1�nR�;��3��/����J��/ى|�[�?q�$Կ�2�U����i�J�3D����r��r޻̶�>i$�0%����j;6�$���I���K�����ތ��G>~�;�o� ���M�
��qw��m껼�L�X}g�e�p����6(Z��U��BGS(�,��8��R{�L{Y�?�|9�ҧY7��U�X�4ɠ�$�f���p&���o��!g��Lͼ�_7I�b`<7�C��~�N;��t^�7�4I(���\�T��\!�4���G&�K�&�#,k	v\��s����FNm��8QƧp/��+�A� �1���ƹ�~wa�v�2"���`���6z��c�6<�*O� �[��p��i���Za��.��Гߘ������� 	a-����]-�gh�7�]V�7Q���/��u����ysO8�\��-���n�$oeBe%�B5ͤ�zXLe־�s�M2�	�x8�^������v�{l&v�X9Rs��L���r�f#�Uv��ʸ����ߚ׭��h�3���u���<{\ᘩ�	W>����]��X\�
A<�-�Xam���*9a�*�C_o@#��6Ω-����(��I��	�a�9�����w�����=-`竨'݋;fS��oak}/�'{@>�'|u/����ɑ:���9,X���5�^rrp���K�~��%�#���-���7�E��7{Z�uH�Uj�=����f��X�05=����]}�>�P�{�D�7K��E�pQIW�F�Ϋ�zh�d�'���Ϯ|��&�����v�$/$2�f��ܼՁטq:L�9o�]�c(�1�E�gI��J�e�DB��#����\���)c��2���I2^��Y�-�=���O����g���ҞK�U&��箄�������bBO���^}��y5�M��eQ+4V�IO���^�/>oKc���%N[ˣ>�|�\���.�im�-�sNݬhy������`�K"-A���Z�2����_~^�E�w˽  "UbTb���c�E�]��z�S����H�A=��LSO��{�,˥;�#\Lk�D�z��=EE���"��x���6J�[�=���Pό�X ]n�3)�'���74�q����&RXp����=�G��AFK;�k;�8G#��w�^O�Y�-!�i;�G�4Y���⤉[�?w }i��T%Y7�]�RY�	yǾ�M��X:R6>��e�Ug���W���m��Ze�!mԙ�&@�o��*;�JC_����x��ն(�wƲ~d�I!�� 4�[SO�J؂�8}F)�}
(f vq����|Wi�����e�umEbИ���\z�iȸ�9�m4�V3�0���R32�^E��הK�����5�p'}��A#�
�R�zD��Ŵ�b`X����
��)Qi�#���q˅F9(:��<�ERLXQ9c{=%���@�#���S��!��g���>~�+%�mB�.1%=�������M�X6�"X?��4ظ}�Y8H#���g��Vr��u��ॅ��H��8iS�Z!�`}K|��������)Kww���!Ο��)bu��93�	��^�=28��f����
g�,�7� oI���ة��8%;���R:������� ���g��G�7?�^�L�,gG�֏\��T�հv�=uN"ZB�������".�*O>'�c�9�8�z��g�jN� 3	ALdZ�om�K���zNr�Z�i�Y��|�w+��T�����&�+��V�(�OJ3���am��1���)K�o�Z����[}Zz�z�������gw���@m�_�
%�K[+��q�s�� ��:��|K�$�'�9Wx�4�������Ӊ[ܴɠsU��T��v���516"SƯ��(�C��B�x���t�R�T��o��cB�N�۠���)�7�J4���h�K��&����J�TvR�(<��v�5�᭢e9N��%�tX���e�G�}�����u���?�c>�������sn��
��1�^��6_ށ�ǈ�@�%�l(�c�p�bk�7��/emx���[M �=�����#���ȲcZ����.��İ��3�v���W��r0k��C�J�����n�:��_�"�>>���+Ү1P���P�{���
�^�5���ܘ�����e��*��}X�N��<����{����+�y��h�x���+K�O]t�.���E��w��[	:9\n�����)a�����[�#4/���j�kh�c��b�1+�s/�6Ú���߭,3�~��χ����9
;��F���)��Q�u �A?Ty���T�c��w˭��b��D��vX�3�|X!�[2�t��'����d�@�3��%�QD�uM��V�e�h�7π���j	�1�Êm��_ � ?����F3R�O����3W@�Ep9��Ca%w�{�p8a_5	�Ѝ�e
?�v�W�,!Y(���_�'V�Qd2\${�d.K�q~��yQ4/�]���Zs�4���[���3t�}�Lu
Y.�m|�_<Ny�p�&���9���s�Ȟ�;H?S���HB��_��l��� ujz�ƾeT�6^��ܷ�	橿wdg���^9����6�M�f"�EիJ�q'��}vaY��P���X��)�M���Q�["ݡ��e�F{}����F"���ȴ���:		�(�cZz=I)�d t��X��?�ʼQL��D?�ylQ�fQ�{\G�)��c~�:: �	�K��V;�ȏ���\	����ѧ~>��E��5ߋ2�>��𢲻�p��V��:������3�~�����f��#L1h�&��Ȭ�����?Xh�5�xt�]%0�tIP9�մy��o[�mV!j��ȟ�U)�M�g�f T����X:�����-F+�G�m�ͧK[��6B�~D����x�|����;��0N��t���湱��Ǝ��=(NVnz܆�����y;�����a	�|>�1̸���,�)u���TU0���ɏ���N�����]О2�su��-�G����v}X�{�Kޢ��w7'��p��]>l��\��C�4��p�z�V��h!�.Y�ǝȣ����[쏅��cXK�7�P���H�}]fA���d>M�'�΃��֤C��8l��&�Ӫ[%��>#zx��u��8���h� .~��8|���1:=)�+�����9}�C��]�v�JW÷�KY0l���>��A�AX\�����{�d���}���Q�r���?���T*����(��A���K]��*Zr�yW���/xza�S��H���VM�o�����U�Z՜%�8�9O2�Q�����U!xy�D$����suNk\6��IJs�����Q��lK�G�b"�_���B��YiU �=��S�䮼��=Zʻ�"a���oA� )B]�a�.�
_u���_ڊ
����X���ۺg���{c=H?M�/a
ML����G����p��݇U�R$4�3�,S5�*B���'��)����
�/�pd|j�4�A�#8�.|X�2��O�Ʊ�K�NK�_�_s�o������&"���U+�.��|�Ge5v��w���w@��7�K+=�$��̕���
Gp�	!`�E���ǥ5م8��fD,-8,G��DC@m��D�/L?�Lع+T�#��U�1���d���6������{k'�~&"�6�=vC��ٹL��"vq�9۟rׄ��&�|�),h�e�2L�6LW��gU�dǶ%�4J5�2Q��(:N�c)�f�W���|���'�O�&ߦ]bJ�=1&�Pۤ�h�����g��h݆k&�G�/vb�ڜvEi���(o���)�9;ݻ��AM��OE�E�.|�%u��� �ҥ852��ж×bh�����A�����%*7�T}�K��]4��?+��X��}���D���Z�B����c�g���M�R�s����	w�pr����ݴhֹ�?��j�]��o����w� ��L�o��蘑e���/9L�5��V� ݝP2���F�	X���M�����<p�Α��V��d�6KJ&��*�ڲ�`��eqW( n3k�q��,�}�{�O�L}H����ׇ�<~�R��1,+�R�;&f���h^��ߚ�m�M��ڎ]�p`����j�oo���z ߹�G���F�:li1)�v}��/���8����	K�B�������bɘ9���{��6Po�I�jh^��إ(O��g���`}���J�T�b-m�xS/�p*:J�s���_񫦂jqZq㊻���QzKv� ����t����+�kO�"�D����^@������e1%���s���ݶ.C��>�0V�o��?�8rȢVC��Ա���94�6�n�n�[�y�,�S��A/B�����֨2[�Ɓ�$#P�����,K��V_FB�B� G�G�j5K[9��\	X�X���Ŗ�^�P���p����
J�*9�榿�\s-
n����r7� �͠�����t��!�÷l�}u{��"��G��*�F2X}�}��s�g�E��_�"ujh�W�V4f��<Wg䥶���.������a�Ŷ�ñ(��]�0o�1<]�n��b�ɛ4�7���+ �T{4Dh�3�m��h>���;��Sc�H��~�`��%#-��Z����������Z$b������ͮ�L�$�/� <�^<�[ۙ ��/V�W�Zvw�w/��׵T����a:�2�G�P�1}��V���yb���~��?�t��[.yO���g�y=�"��4��Pަi�S=%��(���V/�~�%��/Cv*��#p�6��p�k�����M��޼�㤫#�,��\��	bozx��`�ո��o"�C�I�ߛ��TM����5��j?�D"z����z�ơHN� 6ҕM�Ɣ=Q���~ra	3�֦�N����W&���6Y���̓\����[���4�Dߗ �!*s�a)�s�cD�d�s���ո�� �@�5*ʃ>�{ƕ�B�ڥT��q�oѵd6pf�*���s��N_Ew��eB�f��~YԨ�B���}uu@x�`��zq�A�U�����I��,��������&�|�V��5Ą�e���F�����G������ի��Qgt����[2�C�m���ݖ%��
���a�M�6_��d)�'Ä3焵��O����[�od��-�\R�(S�}�����kS2���	�p�8:�[w�[��\I�c��r�I��>�e��eT4�g(�]*��݁�A�*���7~�&��M]"=1��"m�ط��5�V2Pa{O�6��V`W�q2xӀYI���i=�L��eג��sژϷ�qj`ͯ�a�3���æӜ�FW4]�E�+��,@�b0Z��"��knԈEՕU(o���m�_&�K��M�ki�����X�[�6e��ӕ�]�{�|9,Ȣ�s��gw�b�O#s�Η!��+�6�V��4������]�$\����DIX�~�o�:(D�:�e���J��Z��q�i�|:�a�>�!�fK�4���*�<���0�-L@P 5�ҝw;R~z�U���e����`��[l�)8.�$� �r����ԋ����<��^�e�n�u���O٤b�&�oɣ�d	K>C钙a�r��F��}F����Jm�����^A�� �yCk�
��U*h^v�G��_3#��)%⧌@lT$l�ߍ�t �&d�ک�G�:`i��A��c�o8_�;i��OQfq����Dl�g�L�Y������#�\��m����5d�t��]ǮSm��|:&�'?��U|�$��3��L�^���환�B�K�b�	�8�g0�N\���Z�t�S�BB�h���̞��1�M���p{�Q�	�"��s���Y��Cz;Q��2|��EP�gB��FW�a�&B	�Ȁ�bd�ˁyS�<�pvp�K�h5�ź������,�����cr�?�G��%_���Vo���+�380����A:Ș�V��;��*�\�E���s`��[6��}|��T��&b���`��A Bx5������c�E�o�m4�i���$��⑚����%��ᐠ���l����������'R���Дs����b� �I���f!.У��"�%����SBi���A���Y[5�Yv��O����u{R��q�߹P�&]�$�W�?%�?W�%�m�*�B����c'%q��tMqw��?���$����K��B��< �1p���J�1��xb�-5�ĤͰN& ������G�k�.q���ye�a:%�Ʋk���$�mMe��u���Ũ{�|(�����xŬ�]�b(Ŧ]�Y�	F�	7��#�P��Ԭ*��l�vSS����s'?�&��>��Bs���1����r�;�X��{�b�>�J�pr��r%g/~�ڬeE����>5�mb��T;��Z�E�}��CC8�ٴK�/!�����9$	�J�x��bg�5lo�>Ծ?b����~�͖5��+��Q[��Vi���q�:h�ȉ%}�T���kk�Bo�_o	�ΰ|�4��8A�_ �W�����{�?Q���܌Q���A���N�C)b�$�ո��p�_Q��ƞ��[��x��ڳ?+nx���f|�q�_?��Z��v�rܥC����j*b����v���m�9f<��.�;0�xǨ_|~!N������+�ŏpN����X�k|�WJ?�h뭏U�O��|���d�|�%JF�k�3�n�/�ޤr�N�6��v�s y�-�
&`Ż�s\K�C�+ͺՃ̝�[�!��d{�zS�V�¿H��\}tF{�˘Y���Z�!U�_��{ʵ^�r|�ԏdNS���ٛM���߅�d��e��j�/�?%�D0I렽|�Y�t�%Tr���}��j��OE��be��Q��;��A�&s�@�z#�^0��Q�R;O�%�N!�l���ӒV�HM��HԿ�ژh��^�K<��.���+�[e�W;-�a:�d
`��0.:O�E���&~��]�U�,;���.|�.;xxe�-Y��/v7���M�9���q��Q�D`�,� W�ul�e� v���O��3Ƒ��|8���e�Җ7�:v��|n�t��SsPw}��|-��/_e��~��|�����sܜtg��4��M���6h���WB�?2x�}�Vu�Ӌ<�׽C���� _	�<�O_��[!�4���yK4 ڸ�z�:Z�e	�H0��~[XK�9ZS(�	�4�F�U�%K&jڴf��`&�ɷ�۔��$<S;s��4��Q� (��Ds�0�o�l?2Q��j�U����tK�5\������=\�m(�[��ه�\�����tB?Kyg�
F�~��~�s����"�kYT���U��՞Rs+�;5�6�*���F��!{i�� ��Y�S�N�����������E	�Xp�����-?���\!}b� ����DŪ�=׵W�����尤�����׮�G7�4ʖ7�!'���yE� ,�}��&�܅k�?��J����4:��܏�e /���U�<�12!T�	�6���*t;�#��].6k����Y���fw�M���b�z�f�[������6;W�,��t��ޜR�,7�&�!Ƈi1�Ȉ�O��|*�рio*1� ��U��W�w���+Y����C�W�x�g�T�:���[R>��SU=�Ъ�=zR�8��ɃhK�a,蔱�*Χ9�[;���c�ø�_`�l��Fn=�;��+D�M�]x���@�3���0-G� ��4�P܂�e̷��L�I�A�N[	!l��؛�!���"q�OB��a<A-�_�8���p��ˁ>e"�q�N�MX1ᔜwy��iq����	5��	�,�$_�2���1	eܑ����ex�����W����F!�Yw�5y���Te�L3�k�>E�����~���m\6�q"�х�`���㤓�.���U!]Y�ɫ����w�8lm-֝G�lDƃ�0;��f6��O�����3���T笽ETW~��
˞��C77v�1"� ߗ��A�"���S݃u$P�5��3b�����Q�g+��������@��Y�2�d��#�:S,-�HnA�
F!,޻��R+%�f�~�;ڣ���]��KK}�K��~�U!,�B���r,�Z��hr�7�V#�u��6he��F��[Ea�{�U�����`耜GِVٚ��hu�Ɗy"��H��-��}�X���%��+R?�wd2˩N�����s/���U���Xw�q�Rlh��4��k��a�E
�����ZE�MȜ쨸,�ܟ�b��׳6J�0���2�NAL�!���`t��!�)I����b�Vm%�} Q�'�-�n�Rp���][��Cl	ɳ�
��:>S7�����`�5t�I�G��{�n�(�uH�]��wPr�̡�bB%���\�Pm�"O2��OR)�i��,��"`Kk�&�4	S��K�X���n|�>c�����Di�T�ժ�Ż���	cXѮ���h�1'$�������\���m��^����?:�+�#j毡�qeQ��L+5<Q8 !��p�_�*5a_�E���x�������-3��p�f���j���aBxk��ëi̬�s ,+C��21co�������Yh_�������t���]�`�����f����/�3�z�ĩ<�%X�)��F ��قh�i���PՕ�S�P+ ����֮2/��W��M��P�>S[�iĝ̣��=F?6^zd�-�8Z�8T�W�vN:�"of\���phl�:�a���}91M���"?�73o]�mT��_��o�І��c�(����%s�32�����!`�7+�� �I�M���?��t��؊~��b꽔��Q�F�~�eTH�ж���S������)
��)�ojJ����[Dr��w��	�k�m��!�3A�Di�O��.��WDd���+�B��2�
Z�C	[l�eP�VORk�l=���6q�۸S�X'QMBL]������^��7#S����r~Y��!j\eq*vY,��GOoy�}�V�7��5v���E1p�� U���+�3�Ϳ@5�;L�}�z�'b��+���_{�`���>	D�ɞl\��+W���"���C+nT�_�>����Wr�4AAF�$�W4G�ej���{��(:�K�)��^>��}���j��о�1j?7����I��ۉ��E�� Gkן�H��X�m}/8(�5�0�B�߂�B��Ԫ�R#�>(-U��&�7���X���K��_4��-t<s�iB��\o�À�Z"�2�I�K�%���J��U�����ky ��=��Gҕ�ԝk=�|�ӛ���`����"���eJC�t�%X���\ӯ�Un�(��n�.u{�ઐ�wS.f���;@�9��~n:����UR���d��f�M0Z��^?�FX��j�x���d>c�Kw5��Y�tEk?~�j�g�+aǧF��ju��k�W��p �pL9�ŉ3�Ƃ�f�MW߻Fa�'��T�/χ\/����.6d��K����C���������'�p�=�'5u���sB�"*�Zx"t��l���$>�xzA�o�'A�s=�G/�;P���eɰC�B,%�0��8�+��LQԊ�98l��\�l���5+ ��i����e�+�	�7�x��IE�f�
6�!ċ弹Z���P�����M�78�=���h=g�����7�-��~���	bBm����iܱ�jE��>ׄ��i+cMf]WH�tG-e��W^1�fnze\ �?vp��iO����**��"(� ��@n�;hWV�Z�յRx�f��/,���7�aּ��ok�_��2�Q�+Z��jYŰ �h#F�(���0���C�`g"2��ސ���XV�ro��Y���M�,$���{Q�{N&�7���N������'e|�@CP9�T`����%��5�>j����Rw޹��5�c��Ts��Ί��͌'�_M�H �#�Vɠ4'�j�z����2N��S] �t`��I$,�؊AI����_�xVGw�������	N�;y�<�yU-�D�zy�#����=?`0 }�t���?����)2|J��:%1̪���V�Ӟ@�e��WC�������3W=y��	<�ɯ&�JϜS���S���ha^���_�D���ل����45���Di�Q����/2�}+6a�0�f����~��6l�H8#�wε9�+�T���~�y�h�s�a�ܰ9u��:�����rG	3JM�]ռ[,�D+r�}+v5_���>����q���3�Z:):+���~�K��\ȃ?��_�Q;O��'�:�F�]�J�#���m�7@x�"ET\a�P�,*�L�-}������]81�<V�����d��a0[6K���?���m�n�>}�0���N�I�-�I��Mo~�O��S�l�2~O�Mtt��|aH���d���n��������>��O_�d��Jm	s6.�����M�z3��5�d1����1E=?_�V=Z�g��4�e/��1�� &����Z�U��Dz>����@�����|�3MӬug�OƬ_��� `����h�PB�s+.�Q�R;��?`4_�@�')	����S[ȵ��ja$ G���5����YH�	r`�۩��#���ŗ<$��#b�{���B|e@��i��u�U]�j�R�C����}ejp@��j��i�p?t�q'FXF�~��y��8(C���v�{���b��7�z��ۄ/EB\��.��[�c�򀜫%Yy��	��ԝ�x�2�)%�S^�@��̎QN��a�e��r�aݭ^J�͇���<�s��^=�t���A3�'#m��4:xg�u��q�.}��d|TY+�r�Q�6Ƅ{.5lg�I��
���_q��m]��]ؕ1���¶&�(�zm�%n�h��ؗ>r��p��l5�6�Z�B��k�	����2]�#�ݨ�*����*�����ŉ	�'ԢY�������8���z�R7�Z����iJ�	�Ma[y�g�����ך�����e�ԢvŨ������dsZ飝~��Ί�*�e(��o{�.��6f6N���[�!A�z��Z��M��1?dm��S�6�O�~��Qt��ZO�R.GBU9<�c	�nC�m�*�睟�~ӳ�/�=l�um5|�}��<E`�n^�T��a�y*0cUg ��죲��r+͸�,��Hɖ�l� �������P�=;�l���Mxo�Yٓ��egN3����O��>�g���ء��ﺰݳQ�OK��$y��(CE�nmR=#]2#^��[!݂�o��<����JȈ�LzV��5�c��s�� z�k��m�x~=/��x�-8��e�4��v�a��k>���|�a��*�"�����J*�O ��(�R/@\������������!����D1d�O+%���䶯ψt)ٖY��I�u�vvڔ��q�mW~�lLA����P�\�
�O���i�p�X��t���P����yD���i$]�g͔7�2;H��y8r�S�v��@	M���G?��Y�Z����8̗m�4������Q�Q�����"�v9���F�M^�;c����
 �	�qZ�'rr߰Y�9����M#Ja�~+}��Fm��ܿ�m[z>�zi�*���&;>HS�e��L�U`)L�k����L�ߚ:��3]7c�G�[�q%���ʨ^F��<s�8}8g,/;�� A;�z�X�'����#[4��B�C����'����aT�=:��k�#j�a��׭�����7�_KtuX�Ϡ���T7���W�q�� ����-V,����(	�*�F��t���w�f�� 8_Z� 7��4�-�x�ַ��}��f{�1���+�0n��f�q�^��)��B]���J#���A/�v��O�Ӊ�n;�	�IYkO��&<�f�q�I�p��y���s��T8T����%]����;�����UD�>�%����$���n�C�SP�NA��A�;�k���~o��?�r�yf��9����h8�`���U�Fg:��U�)'�_?���B��E��$�����nQ�Č�V��Et:�fa��{j��k�2���u��S@v~|�9���vZz��9<s̪I�������u%󃥐��CʩԎ�=&�@�[󠊂7�O}�� ��
�\z���hU�̝a�Tb1�)��}�4�Zl��$��Ky!��vq/,��Y>Hv�9�)ZπzX�C���B�M��u���c�@(�M�)���s-9m��q�V�H~׾�7��(��k`���Ic͇���`�T���kM�beP�@M�yH�V�&~.�����q(P0V��%*�1=';�y�p��%�d�U5�	�C?�W�3��6��7�.��؜�F��l�QR�T�Jag;Zӆ������|_SkǅS���JBV%�K����"WL{���������3%��|��.�v��,֤���Rg��S��	�yVc��P��Ƨ�WRe%O���Ԫ�7B��Q������5Y�����2ʞ�^a]�n_)%a����ɤv��I��5����m��j�YwS�@���n#�l���Â���`�6Jq�~cѨ��ȝo����,J��a`��'[[ķs����)���Fl�j2C�mתו���L���J<g&���g(�X���Ϯ��^�]۝�5��^`���$7���,f呔w�F��0KvE���X����ͦ� �ke4��n��'�{����ۄ���ӎ�-dᖸ5c�:��|�,���w���k����U��m?��V��K��(��zx��?A{vt�3�%}Ѥ�3W\�l�����M9���ٝFX䨗����2>�L}	���u�c���c���T�FO�����[+�&\ � ��>@{�"���y$�	���)Ž�����G9�1x�=.޵�9���	<�vo�U}��9/S�����i�!�yHYM糾Ox5�A
A��E����x#�oM�Eb���uL�wj���笠4^?�Q���eT|�A�G���:�ޫҒH.��~4̏k?%m���u�U:�u`���H뫣3��ͯ�Z�Oo?�>_T�y?#taT�e�D��od79@�AU�v���\}�EK%�n&ڎ��K�2��;vm��g���A�n�#���A4^\Dhx�R��Ւ���g��Km��Q�΄�^��y�x���V����$j�\��.�ћ��G��2_4UVd�54w+>��W�Nv�_����<6��������7d�ٝ ����b5���\J��z��Po�9F.���V�P"s���x|㩟���Քg�ri��)�B�^O�g�_����#y��ۖoЕ)�h��}�J�)c�Db��b���t�hU/��OnfsC#�ZjZ��;��̦.��>/�U�D��8�F��U" j�3Y7m�1o^=J��ׯ�xs�L�D���"�!3|˷z�NjѺ?C�p���ZZ;�~�[��"r<���*|+#Nx˄�L�O��u����LPѢ���v|��?{2Df���2- m�G�\DQ��ok`ա�ʯ�Dc�Z|ь�^#�m>u|���Gb��q�_��|$ꩅ>XK{�I��㵣�$�/6�$ۖ��0�K=I��q3Z�g��2A��J����Sg�|�w��IT�A䈐� ��w�]����c��űO�?`�z`64��sVE)>Cʭb���a�ԟG�>�|�h���5�N�vLu�o��i�~yR��bDN^l^vmD��F}@�+�Z�x���I�@ԙ��� ���a�zb��Py|����Z�x@���[�wO����H8�e�^b]��b(��5"�R��]ux|{v�&?J�������^G���_Ӏ�F�q����vP�r|ٴ哀l	D��6��
0��b9��3ͱo�b��P��04^�h����P�����_i�"
��aH�:���~�)�4� �d�C�t8R��<�f�#�q@J�0�{�����
,��Uj�����Xph~
�^2��S��2�o)�ѩ�{2�!��D������>eYXğ�>�D�>,h�̂~A��V#dq�Mh�hK@B�w���v摒|:_��5CE��>�m;�M#�3K�U��AܞR@����B?�����+�(��
��笊��4V��G����DɄO�����OʯVˁ�LH������kZ�עmِ{q|V�<�R�%�%Ҷ@[�+�����M�H�(;���wGZN?�D�l��
�z��$�7czEyw:wl+�/�������m��#�_�g�a��9��]���@ꨌ?̭�"	q��
:j�h-C�DE��� u|�Z(,7|X����T��&�����������y�i6��ޖ�]��|WY�,�^�N�
�s)��`��xT�(�"��k��L��R`m�;M}٩����G%c+K���Tz����,��X������ǎ�i���]gMTYt�5��Q6�J�/�Z�t{ʰ��7��e�j����E�P��y�S-�ܧ�Ʀ�����Bi����
�׍6���V�m� �:�[H�d�1��6�D}ѐ��gA�O�ړ�Z�JF�?@��	�E&��4y�9R0�(��&�M#^fgX�5��!s
\�?�L�����ߍ1g)H���3�L��F����R�m�_LM��#\ O)�ڄ����mWVp+`�ߐvn�*UO��L��gD�X$!�õ�G�j��c�i��9]4O7i8�/��5M�]� &�Y����*��z�'��W�l^���I{�0�E�t���2%Ҷ{�b�f��G���r�
��\e�B�%~���Z�ax�Rg���&u`�|���%���~��x4H;�g���vB�C�UT�ج,�._#z>�*�m�/0=���QY��&#n�F5���`��}$t�s���7��F��e�b�TקB8(��Fg��@�(�)8�4-��
%;����ˌ�?7]H��@+���,���Cpwv�����m�В7.*�y��q�6��ؔ�藉�J�p��M�V�)x�n`�F�IZ'�]�?/�	�V1ԝC�� ݧ�F|�B���F����[A�l47�˽&���w�Sc�[��Smx���<��\�uJ��9���t�y�2����#�[wP)A����N��)���"���&.��#��iz���`�dv��%�'�ئ$��jC�cQ�f����l�m��(0�n�/7GS�K�d޵���0�F8EbP�����-�	��+?I�p7�@�fO����d�5K��ð`��v�D�cK��<fVN,a��=#Q�����seN*����R5���@��L�N���'	l̋��g�V�JU��i�/[A�_��H�K�-�3ּ�Vq�!�h���C޷&�y�W��*	]������72'YG�+y6Y���*��"�W6~��7k�b�z�M7�(�a|�uv]z#����Ǚ`��f&�����`Xⴧh���R��.���ň
�s�:�.� �:��%��m5����۔�qk�ʒ(�%n��;ҷ�\�F:]�������jϠ�=*��[��A,�J��8�Ð��[���Hc_S9h'<�_�)Eӂc�02�ŏdR{�vW�a7=���� �~��!�e=T�	5��7����3�¿�����#&�|��W~�G
�ZӢ�h3��@�C�vJ]]���E�{�����y�LFM>	��y�N0��m�/�Ħ������rX�c�~	s~5�{L|u�P|P�C���z��o�D���Z�����<��2+ZK�h�0Ȟ�*��� ����g"ъ��bh�����AbYX�R�qJ�,mt�`9�f;��y���N��%!X��.cXq� ��\��'q!Ѐ�x6H*y9���#��%l�^o?�E��3�:l.�l�[�ȿ��V�*�h|y�����������[>���!���^�Nsz<����X���WK�nB�,%(}b�%~�K�!�95��.�{� ���}��prG^�e`t�6�˯�{,�r��?��q��^��,�8�t�ޑ���e�_���9�)�n�*�K�%�����+��ᐮt�ֵ�_Y����L}���8)Ǚ��FZ""���6=�m�
RK�ݍ#�̷��B`gAknZ��Ú$$5�m��Lhn�}X��`�e5����O-8�NOV�����×d�嬪��R��M��K���^�D����;Q�+̐����{��U���?�Ǒ�F6����8~'��N����q��^io�|��XG��kۆ!P�uP���n}���辺F���{��/=Y�j��(��r!3��o��ד�����<�K�9b\6�-����t�y��@FPlg�Cm%�#��OI���w$����qPh�JN:'���W����`Pi��܍3�Dj�g���{[��R�W��>�eqFɗ$R��\�5���,�z��>^�}�xSj)���ۃ�U')=6�"���RNa����#�B���4�Ugf	���H[)V^����-��n���r`�ltٲ�m��Y0nOr2C�n9���n��em-0.��V��kѼ��[Z�.� ��c��1�a�Vb��7ڗ�������KI�ks�iN�M�D�PR-���Е��Ȓ�F'PQ����"���S`��x��ZA������e繦t��d3��_�i� DHe,�Nss.�����b\�$�5�Ϯ���M�x,����29�T����y��ړ�ש����j��	�x���vg5?��{�nk�lb�EKߑ�̩�+�����,3��ZZ}��%d�פ���0&��L3��|,��ɳ��_	�}C���Shx ��'�솃����j��E(]jM6+{ٔ\uP����[,�֟��? v�-�ל�`��d�M��HUƤ�p6l :0�ْG��#�!ZhiV[�C�O�+�>�{}���zK��n7����>6�?M�U.r�Uj�/䌴�����U�b���J�F��v�C���!%8�<o$�:�E�3�9�vD�d�!X^4�_��΁J|�w&.U��Im�iz!?�\:E�&4�L,R��ǱG�0P��6sQi`���oӉ]���hHn�:S\f���a��K�v��n�d�5q�_lC>�(Xx��@T%(�����`�e&�CR˺l�6��g|�LnU��+��3v�J� �1B�o��Yn�6o+��^��0����ൊ�^ ���0��s	X�rC��;h��N��ԛ��X�Ds�8��#�pb���.���9��]I�Ȓ�u:0S�)|��O�	,/����1�E�,f����1���_m����$��t�=!��V� (�j�}KEb�I�@�P�^f4�IhӔ���gd�������|6�� ���&uH:a�~H3)B��b�v�ͨc�z��&B:��b�NkS�e�_�J�C��\�����V��"�=�a}2�q������T`��<d14�e6C=�C&�E=dG�j����}���4���Y޴�)���KjD`���Ĩ�*�;�tc4�(���;\T���НLE��'�
n��s����s#�d3 �������8�S�9|�F��'��%'@TA��x=�����10�'���6!8XF��j46�ݖ@��)մ���S��h��n86��Y �U��R�����a�����T��!���M���㇞�1�+:�P��쭱v�͋xؿP����(�����Y�0c��2�R�=W��i2�7��͗��L��:�P� |<W�w��l�9�Ζ��-��}u�93J�ߨ���>ni�����E�k�nY*8M������\D�S*�ҏ�wtdNl�r��e�BU�^�^�.�_���	|��{��o���R+�L�n}��:�5��;'_JuF��?>�Dz!�C�_���݉ף�5Kե�Uz������"�w��z��٘g��9�c�Е�h��7|'I��vs�e�����E-��/������E�J{�C���=�I|qua��i-�^1��pk��Ȏ�[TM����8��6f�~ʤ½bk��R]����ap-<�����vr9sh�*��Nm�:>�-	]#�!ȶ�)����*e�ǂ�n����F����E��ԡݸ�,ˢ��>댑��lQ��lo/���ԃ����	Ϋ���;F�'��m�.�
��f�?9��n��ꕴ*v��Gh����ޅ	dG�	��7�����K<���5����\d�e�g�փ/ّi��R<�Q2�-3P��6��8J�v�ֱz�N�A�k|�'E1Ւ�d�`׭��C4̆�ۭ��1�@�bI��;�n���C�4�s΢�s4�9��M۝Գf`N��t����i�_�o�:.�����f�2xܾ��E@kjehj��������dkO��>oFM��o��6��a~x�0��!0�[�6��{�K�����g��bF�=�n�	�l�nT���S+G"/�za����g����h�ů�>���B��O�=���(�B���G<;�(���"�y���N|Г���Hg�����w1{DS$���t-�8�Q+={ن�)Կ�tW*�)����ݡ�E¸=����}��p���
m�p�´�p&��?8j�+o��/`�ԛ��U0�|ZY�M7D9U0&=���a������k���Z΁6π�W\;*�ԉI2<��O����{�q��K"e�	G���AJ����(�@<Nf�&���'���+���]]�� ��Aٲ����KTp��<;8t��4&NZy�r���b���vY��ƺ��!b�Kv!途z��m��X��6�XP3t�=��`��v����q�j��¼�%��Pn>e��N�G8]�.��w�@U��ҍ�/e$��m�U�ފ�6j+P�n�65��74�%����}_�Dh[�ͧ���&�����E%��J-��j!^�rS�9ԙ�G+�k��5�KZ_3�6�횴�8�χ�,MV覒b$Q�4�9�Z�Vk:��=����%E�Ɓ%g�Mϖ�;��A{�4�����VY�ں�on�l�/��p|z����7��ٯ�6BV_v�c�	�Mc��W�"y}ţq��{�9�[�`�k��%R\!�Bw�A���W(����j��z*|]09Ф`��f>��ՁF	���n����y�=���t�W1�њqB��b'JHJP<3{�H@��^�)X1,��WU�߄>�u&1L�?���;R��ɨ8� ���qH�C����j ���=�M�=�(�5���*ͥ `nS|3��9�5B��0�`z�<���ON�f���@�y.���E�X	�U$�����&{=U������A#M������P��Iͩ:��Wa�6n�(������ht����4:�G3��UX�F"Z w��}4�~y#v3�k�����2��L������#����ԁV�+:���]d���k�L3^츚6i�j+�۴9J������n�I�>�%�.(6�1,M$���"1_j0�AiO�J���ґ�`�[���d#VLC�ݶ�cZ%������w�ƭ�fA�eW�As������[�2B���c�]��Z�6Z�Ғ�hJ�p[$S �p�BF𩸉.t��O1���*����=���4"y;�C�!)IfE�[_U6�)f�����[��F]v�����-U8�mp�ƼS�������~`�l����*-鳹.r��s��,`��$g{��Cj�NU8�>H����7� m�`!�i�*2'o#M�C=Ιg����Ǆ�3�ϗ��:n1=�|����a �~�v�����,X!/\ҥ��� ��[q�娽.�0EW�;G[-i�+8�-�kxQ}sJy@/	$!��ZYџS��nY}�!�U��d�w�Rlఋc���n���G$Z���{uoƹ������2S�J�E�g������D�MU��#��B�""����I ��c]�H�Rw�>��K6�Hd��
IRHi�b���i��藈ic_�Z������!�|3m��@G�1�D��05K;|�SO1��Ͽ?JF0"�����Wӱ}��'�a6ݐ`�T'��AiRnX)����B�L�B\�J�6���8�Rc�x�ˣ���+J��1'�̶t�(9�����<�}W:�t�,�Gbv��Ri�	V�x̵���`��E$����=Cd|	dS����B�w.�i�3����Ki"Eψ
5�¤R��<&����5��N1�����f���K�m[z����ry	�Y�ZsIdS��PxM��i^��|��]h1v��K��,v�א|t]	�3��|2��\2��DG1W�������_[��z��BB|j��3��]�� D1L�|Ɇf�q�W�h��a��E��2���D��ӈ$�6,��>C� ���a�|<�Bt�����4	&���Z'��.�zG;���V�pǶ��>��`M�������� ��1�9�����Ӈ��A�`��Y.+��х�t�2sb��Kn-(�w�|-N�����s-0�*R!�'f�"<�G#��D�-�]�&��	�!�$�a����k�j H�Cݵ��qY}�ƈp�w{����xI��ψ�>�یt��+8WTZ���^����H��]�����$����Za��GWWPȤ�2�����%=27{Qy�%�"�`�T�s�N�ϭ��٢k3�����I\KvG>��eպ�d�Q�^��D/�$��^�o�궋��*�^��wա���>[NC���e�����=�l.�K]5��T66�ݦ��e��ҽ~=D��&�M��Sb�����oę��y(�G>�*��<u��ӣƅ�E�Sˍ L�4�����Kh�o�������I$B1��וj\�>��Ǎ�!y�~X�6�m��~�xA^vZ��?`)�7�UY�H�-�:J�hg	뗄�"L�h�<8M-��P��;oٮ3)3�J���[��݀x,&����h���"tک��N���'�7a�;�p>�I6�x��Ƀ�VJ[5L�M���٢V.���}�\�cX����
$���}
@�=��am�/	���©Ce��%�J���F;�ǳČ�v���ܛJtř���Ȭ-!<y�|_-D�~���xA�4��h�n�:o�"�A+U�2_��>������忁�t������X��(gq�@�=n!���D�^�N��fIK����D�2�'sw�Y�t�U��5L�?x2�z�ɝ� 3\���[�����i#���=���0h���q��ߥ����O`B4H�8��_Y�������\݅NV��M��ػ:�A��R�`!92��ݠ���Mp�i�k���m��x-X^^~�g�;�'�;5��"i��9c�.�3���/��A?2�֙�ԒڄDS@����mQ�m�/�9t�J^Se��-|�?��_Ǉ*�{���0�v� Qtl8�.�ܡӼ�jF�5��5{�ܝ&f[֝�ҙm��K� ��~�h>�k9�	�XImo�s��w�^��5H���t���k^����D�6�wJ��� ���0F�mqX����!�\�8?;|D�����kL�y�d3�UYs[�YVy��v��5��W�F�4A;b����\W�ak���^H�pj :�12p�b�١�S�����d�jG�Ys��ϷG(��ڍL:�oo]��Y��c;�w�WP%�)�?K{�T}��������學0z=I�6��o�P��l+.��ɀdh�{���2�����=%A�"��%�
0������j&����r�ҩ�(���?�����n�J0�q��V-���-6Nӆ��^9��`�o���m�ZKM����I�a߭4�ϲ�+�f0d$�	W��SP�c�5:�c�0f$���,�k��Z�V\�y��읆p����W�����z��0cSB�k����xBB �����'����(�GMA~b ��g_�&[��8�������H���^TD��y�tS�Q�s,\�1�6�nQ�kg?f�qOѱ���-��F��
iR�Yg�"��%d��m��@t\�v�lnh {�y)+���E,���Z��;�~�w��M(գ�i��鲚��E�*鍂$�Π6��9����s����v屷r��1x�R�(�R���nZH
�^Z!x� �Z����W�('�/��r)[��n�ۄ,)����^y�j76��x�^}}_�_B�E��>}@�ب�f|,�	���_�ϰ�ۅG�#�6$�(�Ev�������Y�E�~�j�s�l��][Nv�n��G�/߫E\]�)y��~Q��d^智m�S[�U�o���������pW�WȺv��-v3� �XW��rzKdE�'��c-�HtH5�Hw.�/r� ���T�!n@7��ް�hs2)@��K��(��Pf����O��+4�;Qo
�(�G-�������nӚ��m�U~�>0*-¿������D�ym��ph[����M��󦹵 ��Lv�;8��p���۽������!o���f���ҫ���c\Z�A����h��
��_R*\;w�����;�/N�B�x��ri�4(O��^�W�g�-z�3�fH�X$�Eٌ��yg79s��ӱm�UM�Oc�6�Ɨw�,�]1bh`WR+�Ƙ��c�]��ο������d9��Qh�34��Ȟ�>���bC�=B�+�-�f(n�D��V���+m(3>� s�:��=�������:x }Ñ�I�}�W��/�/���_�����6V�ur�twJl��+�!bN`��M�c9m�dI[���}��_mQ���%Lǋ���~�_�4�:=�������Oo��p��V�+T`��S4��n4Þ��x��^9>Ǽ|4�*(�#\Gw���q^�"��9���M�8��6�����؉Ij !��ʌ���D�a]���!	�ر�J`0�ʖ�fˮn~C�P�j����Z���y��qA[��1}s�C�/?ǁ@��Ĩ|I�y҅_\7?a�CX��#S��m(��'
��y��~�?��8�h׋��0=H�f��@����1����Ex�J�>p��'v�n6���T�+��)wA톗�����������h��99�B�ԬW~/�:�e�G��i6Ue�<��U�6���'ڂ�j!��! "�W�D.�� b<��RY ���Elŗϛ�֟�T7,��LB��eN���r(��x_���Z�~-��%��Zw#�K�,�Zl$�i@ip|�e2��_��	��+���J뫉�*��K�Z���}:�E%Ǡ���=�9o��A���zۼ8F��o��%���N2�)�7˒�F��*�����|KAj�uV��`��n��!�O'|ٿ�^��V�n��+]f�n�n�~X����N^]� �}i$Pԫ
����B�6��PŴBzd���`�:�[H�/?� �poLP��B���E�m��|�ϼRT9E~�_�	��o<a�B��D�ԛ3��v)����ڵ��9nN�&�4�o�:��s���.�
H'KQ�-�y�?CNX�n�=Q�c.ȚK�8˴�y���*8b������j�ҷou3p���vN��
��6߾h�:�5��h�D�1�d6�C���$l׺)1ŸF��%�h0.>�
{��L6	���\��hr��B����13�ߢ�AI<�ұ����ϰ��2K������&��y��g|����ǥ�`�BFP?�C�u��AL"S7lp��B��m���mcJa{��ry?�)>��A�7Bf�M�����ODӮ��w�ڨ���B���7`ݘ4:I�l8#̐���5k���y�샅������"��$�PO�$� ����~Y��f!���cp�4ԋ{�*�������F�J�0dp#�pF�1/:�:�J-�z��%n�|�ի�-HXTa�K��g�_�]�x��e4�S0���5�����ˠW��:�����)1���_�]O��2	0Z�c!�;�Qq��)���9�l8Rk��|�-��>{�9깎4�^T�v֙�\�	����wmu>�y��c"��m������t�/h�{}]�Qx���)��G����H�@zU�n�u^����u(���[]Z����ɎǙ$d�Т��k�<��W)�����ܹ٣&2J���j������>�����7�:T�Js�C��C���5S�7��x@�U���R���7���^A�N��|������+'H[��S>$�'����s֋�d���-�1+�_P��~vk��&���soz���2Ρ����!sm�A���[�����w�����w��A���t�af-�E�O�l�}��Z�F�����M[��8m��J�"�܁��:�r؉j�'^��t-��R���`��'L�lk�:]��:�����4 ɩ$E�/��dZa�3/����'>�$��C�d_D�I���)>j���d�A���X�)rV�J�a�6���:I�����8��+�-X�r�9�I�qz�������a6�tDh�J#ab*2���2/�ٺ��5�nH��)%0��d�ĩ#�7`��AsT�q�b�G��u��3�3��ĤΔ��)aG$;9�5)����_�/�V�d�K�;����u�؏yPh*�:��:xl��ok�y�l^`UT-�Hԫ$��Sy}�n�)����I�K�Rn��+G8'�Z锆�	�	���[fS�墾c$XBz�l�,�`���O)�Kd8u.G� �0I��U���@�Xx����01�b=�̆��2E�ѳ�{?}��΁�7ϧ��;Շr �WԡU8Iyo�5�

��(&�ș�U��Z�:=����2�u��O�;�v�&�.';I�6��]m�]�M��]!X�ؕ�"G�]̳ߤe�w-m"�蓗�c��ؿ�Jvo�[ﱏ�Ǩ�mB�F���!
������}o��J�,*�*g)�ʹ�_�f>�B���N����(����ؾ��_2����V��ha���i[��$��or{�x� �Ⱡ���a��hA-��m����R-
�����<N�˘�\�`K����Q<��Y�H2 �9�0OL�gPxh����K��KO��J�9��7���[��9�SP*��=#��Q>�������Iy��wo�,pw��aܼ��=��a`*zZ;�����N\��9GN�>��8f��;�^C2ߞ��_L'��G]7w�{��r/M�[���R�$�.i� UP�lX������7t�1�Ѭ�v�u�]#aRl�]1��:L0�ա��V7���#(wp6�bH�J���][!kI ���%�ED�H��݈�y��f֥칆V���w��ľe�r�Y#wa'	d��en-�s���)oq��K�J�Xa�#��L�����81���+�Yʣ�k�$���N1�� XS�s\�~�a���YfkKPa/��.���1�����H�[���م�����x��;��P�hpg��#'(�5���?ڽLp���X�_"�&����0s�D�������H�k�"U��`���΢ѩ��c�8��_�a��x�Ҏ�8��¾��������.5��(�eac�q"��X�`猿O���*o(�#��i&���Z�܉��/������ \�:��<7Ԕ��.Tz[�0�R� �YG�b�G�V�DT��'��Z2�(̕� ���{���5�`<��͑�H�A�7t�n���D�I������
��s'{���H�S$�?w�X+g+1�	�,����V�b�x�@�vg���ˊtC�W��������?	L��8��4_7��8��)M���AS���M@���<.�e-��^3�V�����;���#�}�X^�Y�����Rb�{w�6O����g�{ޮsb8Z	�xg�/(�)Y��!9Gk�����#~��`yj{�?�bg�)ha!WR��e��2��9��H�Y�.B�h�!�����͔(������`�����6�> _�%��v�k���&�����DP��߬�q�w����";�����)	�����~])����u�↿a���j���AO��Mڿ�H|=�5zoUe���oD��q� if��k,�*�3�H�N�������LJX&�������-0�^M�l����JK�^]�x����2�C��H(�]����ᵛ΢N!6�?0�u�;@o����O�XBo=�e�K����[C`�,���N ��z����da�>��QP�>���J��A����HBk����?�03/ЏD����8�W��ED�#���ĤK{��-�|,���?������J�-��%���?�o��uGӧ��Ȩ�ǯ��1�����ˆ}8B�,���ӕм�c�it�J{E����7Y/��nր\�?�SlHf�H��q��LOdy0����'�mP�a1~	&J�y�?����̜�}��be,��j=-ݼ��"��I�#�����0�. ��Uʐ�K��Mz��:9Zb�N��8'Y�܁/R��G��+?a�D�����K���{�*e�`�<!�&M����iL=U=�*��ՂGr�q[�]�G(D��f;���4t����*e�*��;q揁D%	��C��uYv���V�l���Kd�����z6��k�h<�α���qE)�Z_��q徙h+$ڊ�u��
��]<�� ;!��"1� �����6��P��ɞ�/H}8�w�2��F�y���fvܧ[�9f.��(NT�|�j��~F!�B;�s���r�'�g�O(�֓��jz�����k�to5�=9t��i��vN\6I{{��6��i+���Oe�����9�ӽ�h��J�#�n��U=���&��:ty��n��.�<�{�}�b�r �MC��&�����6ZCa��{����:b�����0�T/��1�l�¦����)g�]Xē_"�J~!)��v�I���No��˯n���ΰ'������OEM�� j�ї�s(��v�����j��J��*�u|R��1ڟB']����}:���%�}���3J�u:y^�0�J}��$I�����`�!U�P�d�"�t�*�h�A�2X
	��C�\��ڡ�\�=�����Z�ҡ�q�mn9�����urňr&Yp��H�wGO���&6{�k�˔����.���5�L	��Ij�6���Gm��c�*J�o;���֛?:��}��c��ݞgs㶷�݇}!����N���3����#����������X$ϣ�����K��]�湺�ߞLѿ����|ƹ���%�b�������%I;(��
��\�u����X-��e]��%Ǹ��F�⛉o6�|�}l c^m���h�rT9�V�K���a�m���4Ց�,�oeEW�3o�gc���J27߹PW|ډ��ߣ]�;lNp�v��Hie�Fy?l-�Q��� ����	����mvչr3>�a�����2��`5�3�,U��1w}W�]+�RT�_5W'��W�����$�� ��Zh��l�v����S�|me�D:|S�)�kX܀l�h���VKƦ\�7���w�l�:6�X��Ab?�ʤ8����-��^BD�.Dv���O��J9v�"�"!4�#�jU�Dtv�V[������l
܎�J�u��|q���HW�ƅר�y��֜���q��t�9k�`�F�o�5 �$n��ر:SA�m|����\����A��ݙ�i��]$�8��(��27�R�2Zz_f���Q��f#���?T�J�,�m�f�~�f���#���%�e��J���������ČzmVxe�o�"{�R�K�^�p��fg���KGo5�33Kj֩��T'Q=�һ4Xj6Z�X�a���]�;���m�T��SD4���������o�3t���|��gQ-�`ib��Oɓ��i�w�!�=tT��ފ�K	 a�ۘ	\��Y&���SL��k�b��h��J5Th�7[�a>9H��*�t#��|�_4d_g5���%QM������φ�!UI
2W���D�(���Ю�{�3�t������3�%%^T����������t���'�jܪ^�y�W%h��>s@}[@"�{8h�'���V]d�S��mͥ����Z�#H��^��nG(u�� �}�9�`d��#ܾZ|7����\�!CG!����}��>F[
�Z�T�$�M�`�3����Coo�i������ѤT�~��y���P�k[�#/��� �Uz��]ҧ6��&j=�ߚ���Z��_7�B�Lc���U�7xo���ۨ�k��ӎ]V�i��w�n`�h
�kE��O�澬�k|+�I��YG"�|"'�F��,$��3Gh�:��-��Nr��cZv��q����M��C�Ʃ�˘�ʼ��=�]A�ǰ;�g��q�+RdF�sx�5�꒩��,+�eo�S�<O�+��<+����5�T�<z>�&Y��*q|Ғu���s��imq7��ZoQ0 h�GW@�JG� "r܏�V�è�ٵ#�\9�f
"j����s���a ��+�@�!K7Z�S8�����W2��yȄ�HP��-t����]��ܻxdgstnp�?w�u ��FM+2c���E2�]T�U�����wI/i��&L��yKip�!�&Q�{s,���9�'P�*�����������JaT��=t��?���0��}2r4��S7�}�T����k^�{\��Cry��堩l�H�З�F?��d���Ɩ� ��`Y�5��սgr>�1���^�����Zp�)�1�g��W��'����W���%��{�njl��-����0��v�Ê$�|m#U��UE�ػb継#��'��_Q0��4|eT\M�-� ��L���������w����0���ww�3��Z�יuz��K����9��8�y�O���v���כ��K�s��]����تh7$rP��N;�L�׃O��S���
��Ϫ\�96�}2�\v��MR��P\���ݷ�=�=�]���Jz��(
>y���.Q���.�'c�Wg�i�h�S�� �t=����-^�P:+{}����HYB�.�6�������DT-��o�|M<��`��o��̷VԻ�������OO'V��6��HU���&h��>׽'b��)AJ��938nY�<�b<��N���8�[+������Gx��놮��FWL���<�)&V>k(���mh��_/ f�����;����}2�C/;���au(5BAVs��m���ꍈ��~�I󞰹lb�5۳���'<w�g����m�If̉����3,������'�<k
h�uZ���0�����V��������]o债�;mC�-�`��� ���&PY�J���,�Ͻ8@��'����4�7����w�sl� ���g��:`�-����:�]i����7k�k. ^���G`�W��y]@`%���uLX� P ��	�4Ce��û�!类�H�f7Av� v1z*��WN���v�`+��y�* ��6�^f�,"�#h.��ǰ?WP����&�v�^����2�����͓c<���d�_I��������Q��bEKkv�*�/�<n�(s�l�e����wT�h�^T��������$�}���I2����zf�ksg:6dL�-X��;<ld�{��s����e���j��	��q���n��O�%����8��ܡ�䝈� S9z�8���ô��2� }���
*V˵"o�ыr�2��_º**�]2k���8�D�v]<�����F����+���{�U�V(�	�6����8A�A�r�]��n37�PG"�h�!�8��ݸ��y��� ["�?w��@Zթ�ʟ*�5���� ^z����g���C�t������)��G�$�e����Y�ev-]yK��H�͉�����&XkW��WՎ��`Dg$��^OW�H)3տq��=�.�K�qO��09	M��c\N��`0��TL$�K�T���\������&��r?���x9YM���44�biG�:ۦz���x�D��!~0�Q��Vo�7����`��l�+oӭ�R;���AH̳2=F��ШD;�hx���#��ۼnlM(r��ނ�
3���a�����Zn�����^���O��|��}L�h�Z5:�JJ? �-��d� �B�����ê���N���}���n��m{j(�8)}cGYP-�J:e2H?6v�T�W�G�&n�m��ya�V�@��Ǆ�$�S\0�ܹ
��<X�8?|�"�
n����NOZ�<��u��F�9�?#E�����O���"�K��`�)�%��e���@�#��~��I2eԤ:1�T����к��j��c5��֧�x��N�8)g�(^0 @�I.o��jғѴR�fx���u��QSu�~�5e�n�������e�*C������k+��P)/�9��K0�����P

�e�&x<q�7���a���O����G��Җ��#._ٿ�07v����� �ώ���gA����YU�ߧZ�K.��D�Xg6S�L��k��s8��|�N�D��C�~Q<o��9��^|C�G-��UʆW��m��J�Qsɱ�¥�~�m������+{8�����0s��[^g�I2W�e��<kFv�L�ڒ��5�n�^�*�.�P]���������/��<�_�{�C��;��U{n�h�?˒�dn��R	s< ����8:^�C��Y�h�7�=$���Ӂ���	�ڰ$���:�-}�jJ�c2��^Z��)�V�4�C�\g9��79�]�=��q�|��������։0��S��䩮	��J|,t����8�J:��A���aD+vvZӝ��kH���_;��ӟ%�M9
D5��嗑jQnk�퓄5�2��I�.	�Eok�,]�C�Z�v��l�����( ��<���kBA�/��91<]����[ѩʌ��+(C���N'�&��%�%x����Jxn����3jp8>�4Oے+L����ߏA6�:U�%�SKwT�ב�M�>w�,@����b[
�&<�s�!W�����Q���M����j��g�g'r�@Y$��ď���[@��8�<W��W��ȝ�1i>�V��>�Z��\{�98�,νƹ[n�yd��HS�����4����GK��R�mR���]�=�<9��a���.'|kD*�>��)D2��f=����B$#�х���Ӗؐ�L���ׯ�Pԙ/�ȩ10��6W��Z��vC�0<�UX��x6z�C��h�JYf�\��/O��z�F���F���yĈY��"��'H���H������N���C3}��@��ibn�.����*]�MX	P���~�ʉ�kj�R��z��E��A �Y:>>r�ɉh~���w�{�a����?*hO��/��8�w�`>�����z
#�ԝ�R]2je\/Si�KA0h[3��T�� �W��k�|���FG��a�����zS M�1���zJQ�+��̹"�z�%��M��0>3�\a�MY�����<���o^Ǒ^�gV/B�.h�s�=��<U��f|� y�0)�0�&��L���G32���RR«��Us������D�FL<���M�б�h�w0A-ҵ�[u�
gp�ļE��A�K�,dn2�C����Ne�j�5jG/H�T��Ԓ�r~��^� �|&�&���T��L����X-�\*��Z$q�iEMq�]q~R�N2�b���Fv$ _&�C�C�Tcy~�6�Ή�� T��� �X-�l��n�^��d��b������&�bg���GF��ݹ;t��	޾�xn��������`�_1���?"�\ؤv��dk��F��Ѧ�t���)�ł��yu�?�`̢����7k��Z�ň2"�~ʭ��j�h��z�_�]B,%�[���+6I��LK{��^vi�Z�)cvX�FP3��ֱ�=ଜ(k�l�g�:�L�h�i�ވ�	ʯ1���e�����]��4v����ᩩ%>.�!��܊
�z�����xL�o-C�.w�����~�����yR�T�݈ݏ����j�2[y��"��XU�Iܰh���ǰ��3͎�E���	��nL�g�4�+���y�6f����;���"好��)�|�~٩]0�ϸ��d�F�)6;�Y��*v�ഹ檧�c�y����}�cj{�}���(�g3�O�������+(+._�&��kfzگ��(��f�)�@-R���KLc�8��ߓ�w�6�}�LaR� �-+CEi���D���ͺj����W�Ga�5A�n`'g����"Ŋ�����V�W�Jr.R�B`H�|`*����涔ک�) �$g2��c*�?�H�kYY3��h,$�FP'N^K+2��4����z�Z�� ���Mo���f-�6\W� ��"��َ�X�Q�s]
p�3�� ۸ ���os;�np����Z��4��Y��'M��9�&Jjmz{�ʺ"R��>�'Y߬^*�����pK_.��+�fk�#S+�tlZ�̧SsվSb�2�{�ea������^��\���c}�c�@���Ӽ0,�S|, Oy~~��f��ֶ��}{{��w2薻�nNJqt�.�B�q����X+�E��%���9��y�6^)���y�D�6����Ԏ?^���k��	pƩ�s�����?��[��Nb�wRk�1��)��4ݻ;������M+�x
����_�UOu��@Ax�4߿M)M	%v�ޫ�qo%~�ݐ��s5�}�1���T�%���f�< pG�[P�ioo/���ܻ[�Ɔ����I�g����f-�t�9k�7	�n�k�^)5��F�fc;��!��u��1�Ic�//=��Sl���>Z�u�
�O�Y0-�p�=��Ɇ�#KZ� I�$m_��{��Q�cK(�m�!jwk-8���0�C��K�М�#����_5��7�a�7z��7>���8�l
،Z�Ch��M]&o�Уʶ�0��e:=rI���@mgp�i!�pE ����~��]`e�.Ƒ�EEM��r�D���*-mj6ȃ��o����,�ʡ������e>�j�e���jl������ԝ��*U6��&�)��Ө�d'���kb��Y�"p� �N���/,=)TXn����h��
ܼ*�ɝ���_i�Ͼ�f_vs ^�B1oL�C#����������4sED�<�m��N;
�p�l��ʳ%D�s/]���L�DJrIccrK����nIj���)&	^�E<$k�&a��J2,���p��]w�G�����	�D?N��m<��'cͷJ޲�<5�c�^�
a=��W��S�2/�oT�<|n	��x"J�i�n���Т�&fXG��P�}��5J=�2����h�vZ�0`"�gf�.-�a��	���}wW�~��������Q͊�+)�8����՞v7n��np�^|ķ#q����M ��%H���W� h� �9��ED�����R���W=)��>v�of �Q�w��s�umN�t��
S�r4�*#H3���Ԕ6.���J	���z�
sx���^�b��ܞ�d�Ew���]�����]]|+�$ҙP�p�NB�,��&ˣX��Ʋ���x�� c����肬��M/[����bfn.���S�<X�/�H��΃�T'�v�y���2�ۅ��c����t��#���7��w4���lx����T�ũ�28��;~��Z�E*IXU��Xy?�`��yP�����S`#�%��FK�hy��Z("ӽ�kvv��
�v�������
iX%="�|����5����z��g��/�M�K �e�#�"��Kc �B�x��S�e�gl���o�@Al�L�6{DO��]CH~£[��@���oz)J���m-�a���xT���*����T$'��d�e��4<_�F�m\V�K� �`:_<�Y��8ܘT�� �����|�r�f���i��$d�$[N�O#��7n:
���Q#�`t�s�xJ�	|��&�eX)�T�?3�dS�pk��8T�?�i�7����#�L>� 
�'�M�����Tr㲭�#�T�i�,l��Cȥ����-��]��:J�zU5��=q��/Z8�'].���ץRE�~������aꗙ!Pkrr3h�G�뿎�Lɖ(T���#�{Dj�w9����I�`�e+?x�u2s>;��F-Z�{�:��AʆStn���UUM�5N��%ieԹ�T�.�(��mGس�t?��>a2��t�1��������ɧ���	�ث0*�-�O�E��Hb���Ɖ$��eC`�]�H0w�$�Fܹ�1���ʼt��sФ������@����̜�=إ���57wn�>4rc�����o��}����w�J�1�Y���Pm���mZ�U��y�QW�ԃ���TN0�������N�� X�a�� �䪤x�q���⫹�~��1�ېu�7n�I�^�%���jW�d����dG2���M��W��zx�9�~�ajJ���B12�n)l#���dË�N(
��_�'b�T+	� s�:C�ҁ9�{�`��J��TN�Q��m�jc��Ρ2�NWε���h�����(�f�}N����Wp��⦷�"�m�km
|XÆq�M�,{.
�ɉ����`u�-��Tn���N1,%%�˚߲��H�]Ȗ��n W���v�*���K|�RӪ�y���ü`&?��-�2����䜁��i� I����'ѶKq�p�1��7a�j����I]ɪ��{����������o�ԞW��������챊��e ���=��V�{Gg�r�\t���a)/c3��_Z��4ҩ	]�|QL�v�T#�:*��W�kL��D� ���v�C`��c��ܧZQ����C(�r[������Zn�:I�+�t3�"Fׇ��a����B�L��6�F�5j�1�ŝ��@�d���ؔ�c�Mg	���s�ϑ�v_��H˒�ڌ~�
�Yq$$ڿ��^XXȶ~,�&��j98�d�m��&�hqh7Y��􍊑Og�B�1�E��5��f[􎢼!�u|:m��Un3��h�B���E���\�}�@��AѾײ��訠/p�5ŧ]۫'0@	����$��@
D���<�nfs~>�D��\���N�3��<��"	rXd��2��_a*�ws3��Ύ��ŀF,���͆&��s§I� q�OP��7 F��ݘ�;����7(�]+Jc�_Ó��u{�$���j�b�x�s�[:_��?m�UV�T�I��v�*��Q��2���<��ԇ����J
�4(�~R!�<Q�{�T�O�����b>�����;(u�v�O��f<������Z+b�3-\�:N�O"BD�c:D�ْ�;���:�G����{�=�j����=�7)7���::D���v�������Z(��:�xo 茏iY�՗T��9ǉ���T��ja�����l�TLM��V�sN(��장�������G��Ѓ�J8��l�NC�#$�V�&�N�_��Bͩ��>�ñ'�c� 9`x+M�pH3��)�m���a>��ѩV��#��c��d�}M����&��D�N��N��[���)?S�~�%��N%���i('/f�X9��3�H�\I�݄��K�\��{�[w�Ȁ�LY~gZ��o�
����!P��H�`��[���^��{\�iA���V�IM�n���Wv{H䓷��3��`��3$���i�υQ/uZ�X"'�S�(}�@��F/�L��Q��՛���8? -E�ZDx�^��>nԄ���>I�o�~�t���4�u{®x�΀9m M��5���܈̓�[�J���nnk�>{!�Õ���M��'7����ux�NW�7UF�绐���{��**�����k�b�B���jV>~�;����A*��T[���3>��#�G�B,�v����l�+",�p������x�PiGA��8l��N�߰�jW-�՞2�V�r�mz���RQ~"�AR�<�^i؏��\�Q"�,O0���%at�)�hY�9��y��p����.9�D�Zh�ځ�0��g+����Ř�u,e�<�!b﫥m�2�7�o���q]��#���1��i��b�mu�w���3�m��Ә���?��1�� )t�D�g-O<�|��2��B�'�	m��k�O���@H*�#�mW{�NB��0����Tڻ��ר=�$�}|����r����Y� ��\�������΁�\��l��5�ȼp_�2(t�J;xK\��a���#}7`��Q�%S�X��.���.i�w�H*�\����A{�zaF��d���-��T������5-��~� T�s�n�]v����%�V|���,_7+����ݣ�g�����$V�%���J4B �"v	�᝺�i���� ��ĵ�j3���^KIh���߁�|���W�S�&h#nkL�:��[����,�`��>w�>�R<�5jx)J!b`a��v�PiR�2]��r����)c^}��SE(C���_/4׉�w��M���#��[_�������¼�1�랟j��f��)
���y��T�8��e�T>�]��4O�r)��Т_Q<���"��4L�����)^b�L{-I)Chӯx2St��>EqC����	v-�g�+u����'���ot�������	r�s���+Z<i�iL|�PF�0ӵ.�i��P�y������C�B��B ��"/�Ы�3���Q���o��쩌"��Mf�?��2������I*��
�;�1�6D�[iسĪ/��J$��6\���&�ی�n��x<�R��ʭ��l��˳zװ��IY�`�5QE�kY*=<��.�V��$o0�1�x3'���g�.O'1WT��b�c�ZQZ]����|��'%4����� �jv�c�B�'�ُ*��� f]U�.|C���H�]�E5��@�[;u��Q�c4D�Â��qpTo���L�*̙���o�M�ۭ��aߟK��2���z�d�V�Q���$�9l��?���
0����,y>�G8��Ovs����e�Z��9������yv�X1���bQC� ]g����Y+V����ʃg��/s'�?w�)a[�VT�h��x�$,�t�t���?�Bf��6��l�jp�����F�k�:��M+��l��g�Y�?�Hq1�9x���6������&Ҿkh�����dP�������孍�W�,_�I��6�p�<��p�|aa��~���S�]���o��y��7��-q�(�rZ��-�>�M��!�\�� ��RJ��V�VZ�����d��?��:�$r!����T<,��5Ȭ����12�K-!HǭK��-��lݎ_}�׋8����0ִ��.�b��c��H=s�l�J��-|��<��t;�D��#_B�s�Ҥ��QrW�� �ɐ�K��ܮg�a�ىɯPת;Ͽ+����Az{Y��j�&���9K63��NC��jߌ���V�1��u
�Z<��F�rU��0�)��z�i�"O�>[�cǥ��g�C}׉�Xa�tvŅb��WF����o9��S����r`{�~�)#M'�-��8�"����^�i�YfI��7�9Kσ�AUΝ�&�ǋ`�z���(o7 R��<'�LQF�bb���+�ꋪ�����jG���)��[?p��֪�j	잴Tַ�9E[�kŇ�?����N|c/�����>���Ĕ��0���L9d�w���x]���D�գ��ȳ��WxT��n�a��}�y����M*,m�moT"t�����pu�u��u=��Ծ���-�e��oI"��o+.c{��d�|v�
�0c+�%�v�Y�jIZ��}�i�M\ߴEܱ�;r1��K�]'� ��q�c.�u����y�X�;6�f���yLR>��ഋEKo�(��G����UJ?�H�E�ſ_�q ^�f�]zŋL�)p=�C��嫻�=���!"!b����m�>��1Ҋ��]i
�X��r�c��˓�yA�jS��'�U�Z
��Y*!V��=���� ٨���.~/�k6�̰G�D�}�zR�� �:CU%�@n����&�C�f�K��HA�_��p�e.E	��6S��!���̸۝��O|w
�@��T�,ǡ}��r�&L$�<����؅g
��:�{ťsR�;�ܦ��o|�w��Ԕ����
&GS'H�-�Wڇ��&o~�8I۫��1�O
�*6�KG�,���m5�����K��as��Ջ�;J3��)�r;���Ʃ&�]R|���4J�TE ��i�'�i�M
�M��$�@�"����NO��(�m�����42	o�X�L]�i���v�{�\$�O6��lb�^��#"�y�e<�}Qx���+�Z��^|u�4|�$�{��S'�����@	��	yq�u��B�a=,�X1P�St�f�#����qy�%�_�w_�7 $x8X�x]���r$���X��j���S���UU�Hi�jA�RJ�X�U+�H��po�^L��^2=��<���WN�e�t�
κ�O�n�1V��6��G��T>(J�t���3ݰ_m��)��eΛ��8&5T��A{�ޢy�A���?�\���9�2�>�T�Y�v�0^������@���5��ܭS��ٗ�F��X�j������Ƴ����W�ݟ*�|:#���?������'�A,Q�uL�b�J<	�|zSRM#$���8�}a��qhޭER\:'�L��B���`6I���f ��I��zZ�9O�^�<���N)[���ק �C%���o�8B��$	�q���|����Y��b �f67�V�P��"��7�<�	X�@�Z(ڄ��)��#�^�W���`'��O.l���1��Q���� ��������t0�&�Zk��b s��"3����[�����̎�u'��$4�_�Qt��Ư���,u�M�9b�ؾb�DxH�t��6��1���{���2�-��DB1k)��H���r�`\��*�@�ꜫǝ�-"y����I5
d�I4X-F=Z,^��x���:�R���Ƀ��ޥg�0_Ec�;@�u2sn��Hb;z��Pʾ4_dښb7D��8	E��E&M_^��p�����-lu���Y�;��H"ؠQ1T�J3LQ6D� �Tzx�lu���U�Ev�����٣��\ӿ-�M��X�	�Z�]P��x���{�G$�y SL���w�[�_*|����~��Ao;cS�>�X��p߼�/�_���C�Zߎ��cV�Oze����n���X&`}?��ڻ''��k9�$�0W(���C�/K�h$2�t�b賃��imS�P�b�������$H9��#h�o&���)��^{��+��&����ߝ^@z��1-v�8�[U:��*Jz�Y�����ThL��Q��)��c����f��k@5�pZ� 2��T���{=䢯�s��?Ɏ���i_���HBB�`h��0E��R(>�-�phI�6�&W�siԶ|-�l:I#mfUȈ�:@�.�;�MH&���s@�x�����C�҆���Μ\��a�Y�U�Um]�I��<���X���W%�1�FC%zM�"H����s�p�Α�y�j�7�����W�ݗ�E�r�1��/l���*L�Vc����w��K���s�x鯗��L��]_�"{=������[����w��E�o[(eͅ��Ć��9�.Sq���ÜB$�:��J��p�v}�[JT�P8#�b8��M��p. �p�y��]�|�y�w����B�n҆yg�+ݓ��'�"�IGߏ��&V9H\M򹛻Mw>𫩁a����k��B�i��M'� Ҕ� f��ix������KjL;�nN�;��J~;�>����m�]�-�aX� t֏f�©�85�_���-V����������Y��bi�/�TC��Z���N)k~|�e����79A��n�]1�4���:j`�!Uw�����tv�}�b�{a�ngi+�c0����P���Z���1Ŋ�iS�7o���/�v��l����vS��*^V��ΦYv@���6�:�16!�I	���j��O_VȕWܞ�WԜ��3��I*�1� YG�%�@��蒘���N�qɞ�)s� }i\H��bF�x=�1�6"�H/*Ͳ�?����xP���p�SI=��HSo<�7�-�p!m�r1K�<n�v�$bEw<�Y�\��g	L�v^��YsfA�q�BZ�D>�:�CƩ2v25�%�^��LD=�h�g��O�c����u�m�k	�*�t�����)'O�Kmk�q�T)vQ�{FQ� ]�M��&!fI5��zS �WxxD�[����r0�ZlQ3q���j�B�w�o8$u�\�&6Z�b_�&�!I�������9S�큣Q��`>h/s�.�j���0����.���E2h_VfaH����f1m��'[�W���������,��P s�"B�_�1�J2F}���x9���M��1��9�)����@LL��m�n�H�.K�LAѣԖ�6����mC����2j��UE	�����a��!U���<1���er�������h�)euZ�=r�M3��|��N�m���E`آ�A�k�nL�Q3�_g��Q5���'��Q�2N��
Ҷ-�1�����v�����]5�P/�xq��@���:��79�"#銡"MrSզ\-ϳF>���__L��h	B�7ۃ�2ѓT3�*}��RG�%Y�4YU��C����t��~@&fUs�
D2�6�:f.;���G���=ݓ�2��`�Qo������D�������;��a�ZƁ��F�_#4_��!E������_o*q����zr6�}g����"5��"	\�|-�P`[z��ڲ	v>�%*�+�T��^STM�NF�#�K.�=mӲ�T{��3&ҳۨϗ�������f�z]n~]�j��pd\� i$��%{�!�C��%˨�Y��U�<z����Y�0d����ʒ&�z0�eq�ǿ2覨�vW� ��Ic��H|<��W.�|�%�b	��^I,0�D��d��&�{��k3#}(!�:Ց��:��A�Ƃ���ͤ�'AO�t���B�/�ұ%��+���uqjO�¢��Q7vф`�Y��"a]�RP�Gn^��"��l�+�WsY2�#M��m���``�J.Og��w_y�̷��q��i��[��M��!n�1�x]��L�����c�k?���M��A���p�#�Sd�H��Mڏ�C+�jV ��D��i�P�U��X����]u�G-����j1�r=Z_��R��}���$`3�B2��g��KjNנ/�0FKn��;�m۫�yGNfx�m �����}b��0�i��D(ڙ ��;"���ץ�=כyaG�',E�I�)�`K���z%�7I�]<���'K��/kg�?�TК��f�I�1�M$K��6�w�h7�&�.a�#�)�tX�e�쫽I!���ǜ����>�-0��Xb��J��Ч��ԉ:+?Uט����ge�C���N��g����:$7rS���e���ʹR����o�V[������ l�S�r�&��=��d�/�nu������/O;-C����S�D�˗\h��[�����QNT���Ά����$sC�DsQ4J��O���~>�[�_�S��r�rby��z|�免D~�Z+M֧�?�%��G��^1xv��A�z-�\A���2�?��{XA��lp4��2��/�#�r$⢺$|����M��N�D�������N �D�>g��� L|���������h�!LҸ��JFw3��/��(fVJ9[�����L�t4y��9և���k���G��}�iζbUg��T8%��e$.i���<�s��-�oLX6@0�,!� ׉���$�!�U�	�t�����Ӭc=Y��<n�w�D�̟��W
r�pQ���!��?1���ew̌�z��!g�j(&�m;�O��bF��scc�*�F��k����gM���9 a�B`����m�]��`$)~�A���P����-�b���l.��UF�i/IK�x�I�2I���r�[&�l%���(1��P,���4�# �h��~ޫY�Z������~B����RĹ���%X����y�R��Y�}��a�M�7cn&�gةP=ě'���_ %���8'����WO�����sk�W�M#��(K&�s���O�X��L$��0�#_D����5��A��:�����]��c�����8��& g����zAh���1��r:C6�L���F5�jx����\����̷S��	�J�	����5����r�7�~�K>j��|����$�A�W�w��[m��COT{�E��Bg�%�V�;͔�>�a-���X�1k1�K��S���d�)��]����<J��`�FV`f�pv��p���e���T�ePH�+�w��K'��l_�뉃�Z�� i�} ���I�����4I�$d��>e�ڂyi������&<`0|�H�l?�	ΏBYP�[�JЖ�o�V�Z�O�u����A��?+�i^���}���$JƱc4]�U�b����K����%�[��)W�x���l�zf.ۙ�x���X�\~PP&������AY�r~�d��	���E��v(��P�ߢ� S9!�T#�4�ЮC=��<��C�Cw����-��8ķ��JCF��ɸb��,��`ұm�ڥ���|*�����nT��_�uj0�$+���ޒէ������&����EV�-��*ڌ:tV��m �� �$�i�^̅?'�^�Ǡ��cHt�{5�S,>�9���.	S�߰��?���%�t�U:W�o]�F������Rt�� Ab���.�ԯG6�'Tn%���������D[���|�Gc�n�pvU�$��Ĳ���2��������������8��b�������^)Σ�u��.��S��	g=���U+T�(�l��=��>#��֭�%#&:�kwL����=ȳ<��M�[��:��|2�LM�h$]=M��e�2e���q���n�FCn��p�%x6+��%�?����������N��q����I
���:�qK���ɚC�u��u+f���eQ��ņ���� xz��q��|l�C4���hhU(������f�xM�k����3˲�~���VV&BRĻ����@������h��'ǕNN�n�.蠡J;v�/p�Զ�/U>۴�������n�s�j��m[�o���v�ma�7���t�t@�����	�-{�n�59��h�OC*�'���[��b5���p?^x5��Ҿ �� <D��f�7�}�!-F�AnS�^hnc�E7n�]'O�5:�a{��Ģ��C��B�yd�W)���*>�1{�֒�6"�Y5W2���7��.	v��ᬰ~��9tqr#3��o*��}�h��J����9wV�5QMŚ����r �<k9���lP�:�+㭣s(ʑ�jP��'��m�D#����n/e!\,�8on��Ӿ������vź(�BY�'��!�?nj�GI�Dُ�No.���0=m�$�����_C��)��9��ߢ�0:fX��ع�1���=|��B���0^=�9��ﺡ W\`]��d�R�_�׹��.2��vB���	�
v�8)��P�".l�rߪAH�v�M�a����~\LB�
f�!�le50����q�g�A�+�gv���<������ܽ^�tÁ&�}E/�f6��6�q���,D�l~��֫��j�K���~l��n������w�����wPON����7$��H�"�Q J�|��U��L\[o���1/�/%�Y���#%W�4E&��r� r�C,����wq�`�_-����{�HٻV��zI�K'��\�OO���ߎ�%|ܬ���y�;�64"����U�u���d��DJp��($i�Ϣ����6S窧P�;E=
����>��������O�"
���>AA��]��436����?��2V��G�+x��v�~��WV�d�oV�|�9李Rkӵb�p�Ϛ��6������ᄘ��8۸'q�=����p���Cx8(e9)�ѩ1s��~��v�U�I��7��1��m�.�����`�\?��-��y(�+�7��Ѷߌ���cˁv��!���Taˉv����y�s&��b�	���
ɛ���w�#������bA��ۭ)��r�٧��{g�i�eS��_����|���G~=�}��iv�v2�>��x�1��Uy��o� -��nP,����0��8��X�W��S���z��,'�MG��=�����߾:o�o��?'Z=�-��,�1��y���mn�\�-WK�����<�Ǌ?x��޿O�M�B�b-��L�X#ԏ�~��dB������'���V��j�r$

��e6`#��t�V���ԾlW�]��I%�d_N|&g�Z�=t����l��ԉ��hp {t,}���(3zXw9��Q�Ϋ���>L�r�F�ɵ
�ß�RB�hr��Uto����3j�����AI���xVXPa�Ngwe���?��~/}��Ұ���g�!~`7a�D�|ᰩ?Uހ�bȞ�?�:��G*Fj"Ӫ�bw���,^�P����j�u&�v�)�@���#���ٽ�eI$�	��/|�.�z�9�h-��5��3rL�֔���g#������\����8:'܅,ө
���~.A�
��h��b�k�9����U{�tvo,��j�ؚrq5ǩI��;v�aDؗ^��Qw���z�����|�O��y�:LS�"7�)'�ԵԨ^>���B��წ{�נA����kK+���ީl*�[�Z2Mҽ�=��ӭɫ��Rh�d\�S>z��S�ff|���1d���V	y��rJ�>�����x�s_�Ʃ�����qz�m+�l�O��¿.��ON���4�K��b�v�ˑ�n���K�R�B�?S���������PX7������n3��sW�`]�dX����ӱ`h�R<j�`�O�����L���à��c.��y�q�g���&���H`c�}?X��%�_8J�o�;�0�@!�!��Z:��������I� �3�a>��+�O��W���+4��89wG�I�)*5�N�$]���� ���?�|S8cރ����8d/��j��9c	�yV/x(������^�`)���d6�bz�E�o�r�j�2���_��Q:k%\�����)ե��3�	��lv�~�A5�%���nH��v�V�����"mǵ&�&7�޹}j���e=LO0��͜��a\���/�p�LI��f^i�!�ഝ�R�pJ��
A�#�ֳv�n^��o4������y���=��.��"LM�G��G���>������H�:���i;}y��q���v��;�g�4�f�)���r�T��,�^��6˫$|\נ��l�q�#��ئWcP9���O��V3��z���Ǟ
m��wJ�,#��^2dHR!���0Y���&\�p�F�l��VW1�X%���4��=}���������3�s�������6�L$��M�{	7��<g��Y��c}���Z*�*����N����#-e�����n�Ǖ���Q����Z.Ps�\l@����'Xs����Z℟l.��� Q<���L��64�8H�q�n��~6��rS����Q1(���P��I�鯌f9R���m�yU���'ʒ�^�:��<��}�p��*�@��UF���_ ��O����|�:$�`����Θ�� �(\�Uw�9���AeMv��j�g~��)�
#v�S`)&�x�-`^�j�՞�h�,�d��Ԥ#�U2��Z7v}Qǅ>E��̷؞�X�V���i���WrH
^�#]"��8x@��������}2"L'�+m�%͊*�^d�H���r5ù�6�骜��5H�¿..e��7���hq�c�\����.�w�t��(2�k^Ť�/d;���DN�֊��"�hn��v?��׶�|�:m��:�f��9t��M�~(ƃ#��'��1!�b��7�E�l]��x������^��	�/z�i��,t���!c��y
|�'9��!���z{" m[Kc�{47�ɸ�I��U��~�B^�Y����I�~�\�)v�@]e�J�ꮃT<9U��X7B���MQ�ڙ9�N21p���/��7@p���4�u��JN�h��1|�~�ԪX�DO��x�N�A�T���l�-s~-�5�sH��T��\TќY${q��9E���E����#4�b)�P��N]KnIٮ��X�^�&��@k����g��ly�q��KYaHN}�}*$�Q�n����G�n�\u�`f)�K?�\�?:7��w�=����G3��KH�~�O�*�S�;��r���c@x��)J�jl���Jߡ������Н.Д��X�:�~�r`Zp��f�/��$D+��������CZ\��w��9Fr���ԽKش�?���KA��jq�RuFn��
-��]yn����'-3 i$����X�-$����e,,�Td��^�Ὧ�բg�2�K��`;�Zb�9��S����������YB�������$Q79wi[�^$��5��4�\�1+*���?b?��)E,ߥ%�S(��_bV��|�B[6�h�\���;�@;�ތSk/(Z���� Pݳc	$�n�T��+��A���N�s�MmKk��j,���F���A3�V悂����y]�7����g늦��Lv�ߚ��	��̍ԩ�@��\C����6x^.�m���b]:b-;|��Wb֪#Az��0P4����֫�vUp%6�y��Ҫo�d��Z����Ό񠳕A{���{ğmMֲًp�> *fs���]�?��ȓXC{=ҍO���ډ5�W/�\�-.���B�wڻt�����K-l���A|]]�1�R�4�Qf�`�����^�k�R;'�b�/Qg��B��P�y9}Ռ�U�8|��ƒ��!O���XN�mo:Z }ܶ�'��Xùhe=�]9���v��!��G�*Q~�/?1{��d5��^ߊ~-q.T��� ��v��^I%By�؉h��Ew���C���^��`�[��.;��
���Η"��2G�#�3w�����uK�� s6۱w�u��t{v߽�_Xɜw�����۫2�����tP"<]��/V7�� �����n`n)>�0Ƨ\�Zoq���G6{6P�Uc��0�H\u٩�+���6�p4BḠ���q����PG�����o}3���*#Hsߣ��ӖG�s~�E3^=q~�k�Kz�����0�ҘC[��ra��� rs^��-�H�o,c]�U�����Ƙn`�| Q 51�[��{H����Ko����
w���Z�+#[RX�C����1��uJ�;���Su����c;�^ 3�������8;�?\�{��\���δ�����Jf���eu���n�.QuG��D޶��˖��3®���a�{��ԾtL��J����
���z�_¯R���ӽqb����m��@�'�[��� j�_uE����-��B���l��;�5a1�$p���`ݻ��ȧ�dX
�4&g���_k������ظ3�z�d��w���j'd�"S8��a�f����Va��c֍R��������L�&��?�^�A��Q����u�}�p��-|�8fJ��?�<�̛�))"� ���P����v(í�zF1��v����h�w��j�{F�>�H<{odX0�*�����L�~zb�04�R��B�xs���2+~�C��ٸ�ٸڇF��\��'8�E�o���Gw���ץ#�L�bv���<���/�u&�\���B//��{#��Wk��N��U�H��Mb��ɨA����G~�/�4�!�U�W��3��Rz��̺訩3\;�t.����r�ry�t�N��!2WC��]�l�Z��a�n�jј�S n��Q��ݺ��~V�Uhs�Ĕ��F�I3v��X�~�nVu�(�_ F셄�I�������B�j�k��wgM�����:>o��W����'DdU��M�����S1jw�3�9-1;-�Mf{��8�v�cԪ�M�^�_��\Dg��D�a�!��+Dz! �c�L�Ѧ��Gmv�ᇠ�|��>+x�U	�?z���S�//ص\�׫��FIfS{=E�_�n���Xb�GG�N4�rka��uU>iE/[���A��9�z=!|d�8F�xd�n��9�9l���ۧ��]b/VPs�iӈ-!�ᱵ��kH���a�Β��.x�����
�N�x28j�VF�ב.ro�@7��������S�ը9�4F�?I<�zm�=�"ボ�g�H�5hN�d���m%�ݫ�p�	o<��sn���D1|O)�<��e.�K�$��o��/��C%��!M�	,��1����-��Y˹>�V����Ok�NO�E�4�䲂���(>�I,��ʧ$����E�_o~}��d_HT-��l$y�,:�;C#s��ҳM="�-1Fι'�ᷬ7�LW�!O����~���gƩ���l<39!��	�ڗ�Z�)�j_X���0&��z�,7��-i|>�ܓ`�ZL�ո�!�����5j��:+ZΘJYp]V��o�Jyx��1'�.f/�]�?|��Sy=r�K��-l����xZ䖭�v�^d�+(]]/m��tQW?P��;
��K�|��r��"=��GIp����q�W�'O]8.kX�.&���ewt�6�*$0Ю�w# � -���̾�� �k������<�� )�W�a��3�~:�3����-*ymo��:g0jz��k�4Z�g-�.Gzn[mU-i.k��Y�]n���W6Y����
	���O4~'RN�LW�� ���\�ǧ��"j��d(c��9*���PM:e��瀎y�߂C�U?�OSݳ9hA.�4��!_�1p��g�-"�܄baw���}-:s��i�Ml��E���Pʰ���~���qn�	�)���&����+y%F��ᄸW�'5bP�M�T��uyB\�����]����V��#4��9�YM�uhq�9�#8.��cȂ���&�g0?�_�*(�+[{{D�o�>�4I�\u#ĭ���SY��Gۙ��k�g�`���{P{?4�_�kq�bg~㋱���g�6���%��~ւtE���Ok��q/��9Tf�JBq�t�����τ�ѳ�,6����WjQ��.Z~�0R��r=��(F	����H�(c
��k4�幨K֣F��i��Tz S�4�__'��̂�������r�΂���(P\)��7�I23WpZ̾�_̤\�Yy�3�Δ�t���ف�+�.��w�b�H���t�q��7f�
�|��:5Q�%�y�z^<��`vd�%��� ���Jf��h�w��H_���>͓i�� ��e���8$�J?�f���H����R]ge�J�v�D��r�ύ`2��=Y���'\1���1 ,J��d�e�(VDTK���7�#��N�������)�[R/�nNh�sz�&k���w��j������A����>7<������a����*���\ˍ��o00&�)���_<u`��	�B��GO�pvOP/���JLgA!�p65����q��������%o+�>�{j�������PK   �<�X4q?n  �|     jsons/user_defined.json�]ioǖ�+��K��uk/ӓ�D/I���V��T(Ҏ_��>���{a��� �bI�>�v�=w����Y~�H;/wV�i�kLy:Kqgw�KZ\N�3��V�����ח^���?�y���{892L�	�K(L>L_M'o�qu������|���9�-�b���y��~��>]�|�mD\I~�\����ڱ,(p1��%BA\p���|��xw��A����r���ߏ�O�ArI4��G,���
�f*��b�	�l}�a@�w�8��rbi�$%��0�2I�o:w���9>�Z��x�kp�s����,�w^��3[�L//�ܷ��6��JR��e��Ͽ���՟5º�W���+|��a<Y.�	�.�/�_Nk�o�g��P	cA�J)++�ѵ��{��y��������T_����_���Џ.�� �>D������O��`�8e����ON{�y?<h]q��&������Ϩ���o��?��o9�_��?�����P"J{�A{E���p\�ǆ�k��u�@���i1�H��qOxI��_�gi�|��X��}��]^��������ՙ��<99��E|ථ/l9�+o�c�B;EO��%�<� ��6�Ro%}���Hxҁ��ЉX�y�4Q�ӕ�r-fȳЫ�Fz`r}�.Pz2�Z���Z�f�V�+�~�k����[�h�����\�h�7�'�~l���Q㥼;9�`��f:)"���	��Z8������:�qg��7�<5Q���>Ͽ���߸�\S���r�1����"��j�6V^?o�87[e��EZܑ{�sgqU߃J?]��w���y�-a�h�Z�&N	A I|44s}�<�n�S�'����l>y�>�	��>�o�a1Gݖ���6Ő��f�� 5O�jI$d�HH�+<'|FY����4&|�"`S��mb��Z!��k�~������9>��*0o���T�l�0�I���j�/э��Xðm
������$e��`�{>�[�.�c|#�"̡����`�ڕb�Eh��K@��sA�������o�mR�2���ϋ�#?)3��~#�6�X���~�6�X����~ЎҦ���T?hG=Sf�{��M(e���M(^h���M(^j����6�x��C?�X�S�����T�M*^h���*֑� �i�ڴ��~^�6��`���/N�_�C���tY4}qr����1Q���/���4^
m^�Aw���B��ч7���1wJ�U: �;HK�%j�O��l)�@��;"�.����_���s�́��rG�+&Nݏ����7|�cܮ�6b�#�,e�F�H(K	���;��R��Ad�Q�[�l��;�6]�l��;�6U�t��v���0�Q��R�a��B��B�Pt�s�z��m���U��MA�e�C��h���$4�#�a�?�ieGZ�n�I9���Zv�5�,@�L�#�QU���/ndGZ�����Nv��5�)@���eG�Y��ԁ��H:�
�Ͱ�Ցp6��k�>�_�f�
`�;L��6���������S�
���L�0
(���L�P
8����cP@26�e=$����.�aYAX�Um�	�䨠�kPK�B5��kPK�B]��kPK�B��n�A-�
��s�c��F��QݦW�Zz��.AK��@w�ٵ�-�
��f��$*tX����@���(*�w��!XQT��2�ð����e��bEQ���LǊ�B���E��.�aYaTx�e {�&F��+���� ��� @(@&�E .fG���Gw��f�Q�sع?��w����i��ǭ%� "Nd�׊ѼS8�os!DNRҞ�́�d��G��g�c�b��f��j:��-��o��c��u>���/6�����e�c9��?&���
�H8���&��$����{��kS7����+I�惦t}w'�M/��m ���t���!���p+ڻ�ۧ�|5����]���Wͧ왺 �]�p�`$T��-�����QPy>[�L���(CqG���j1M����uH�{|f^����ѦE�	�;�z=�C\�Y��|��,^L^�/�lr�f�M;�_�}�^i5*恢�!"�}"�&Zf`�#,-��d!hHh��Zb�$:mWL�
�A��h��o-$��V?rA$Ӧ���]�5���K�O���oD�T�#���OekpomX�,�X@�&�0��VD����6&mc�6&mcR_L�g�ˮ��3zr��WdV�����	]N��x�Q�(�L1K�T�z�s?R����f�0Hz��� H�<Ya(H�������(0j�w�x�x��Hg�UJ�z$ʇ��ǈ�
�{3ъ~�+a�zt�V �� �.>k��IĆ�7�4sgc����"F�Y��U��>���M�дM�ʡ��S��O�s�(������4��ݻz�gLug۫V>*�lHb"��_�0i��0�.�H�2\)I�w����"S�C�,1*fik�+X�r����M�x�3a<�-Cף����vZ;"��nNcW{��zWQ3u<�9�`̾W��� ������v96Z�۟_�/�h�	��F|�jS��g7����q�.�|'�O��}��%G�69 �|��R1GdV�h�g�eԗ�TF"(CLvcb��
�s�
�܄�q[�&h�4���16�U� ���F���cN��gR�[c,�`��9\�Q[��*�~ YY������ǘt� JqS� �i��!R(@*����@b7��ݘ��W�K`���Pf93��@ZƉ�����u�G�{�ظ?y3_��߻�r����Ҝ���>�!���$GB0��)^�lj9:��8��C@Jbh�$���c���)z�t��уq�J���
��޹����,޿�*��
0��[L�OeTd2��i�&�Ě%I��ܽh�6�
k��}�����}��y�+���2����n�e��v��[w��H�Q)C��	b�gH��y�A3���jt[�n��6�O���||�u-T"�g��VG�]J�)E���djJ�,"�{G0�DhM��H��q��9{���s1]YM9�5o��FZQ��
�B%v��e����aO�`PԪ�VU�u�>e�/�X�@���0�>��a
J�YV���
�I�Gu� Xi�����o���l �*I������t�ۘ���xL�p���Y@��g'n�۫��yR�g�G����)E�	A�T��F�UH�I�.�"D�z��i�ഋޢ�����$�V���#�DA��yl��RR7#&�V�ZӪ��2��G��-h��z����>�S�90�������P���\4'�ZO��&�V�m���շ��6W����^NN��'ȍ�w_?O���6\6���&�	Td&��@���HդlN�)O��[)�%ϒ$�\}� �	�d��LZ/���U�^m�{;���No�!\�M;w�?�c��� K7(s{Q�6¨�5�t�ʬ�tg���T�Y�NN^�׿Hj���_���׫���s���S )	�2�k��B�D�`i�9�@�t��uK�-]�t��uK�-]�t��uK�-]�t���߇�ǯ��l�H��� &j������	�Ԑ}���!�Es֠Lc% "1&{"��	�" ��Jd/�SDf��NBo� Li�2�zb��/�g�g)��y���y##�^�BsEɋ2�W�9��3��:g��E�#� d���w@t��\K�l��Ó���gU�%X[.����F��� `�\��s��Z����ޅ�q��Z�����y����ɛ}��qk_�4r%a��e�D&.$t
Y:J��8��[�R�,������N�����o�Dܺy�)�`��>bV�>�Y[�i��-�����o��>��G����WQn8��^�n��ֲ��k��b��k�zSE'�c7"l�l�l��[�9�-}�pq"�%�D�|��@t��@L,Mr�ؐm�2����$��Ȝ@pu	ܬ�C��Jy�=�a�m#�ls�&��,�����P��&r�Rb^<9�`�\o�|���U}����I��AdX�Y�]F���D��]ɨ��TnD`�#h��[x�4�����T���i��[S.�M��#�������i�]G]�l]�qⵔv���K?�X��/F�p5>*(dwʚ��q��9���D!k��Ԝ�P�~Ke�#�ԃ"B2�GbDr�!I�zY��M���=x�v��y��8�������@W������u��-qh	��>�K���� {S����DJ�kI��Q���a/=_L\��y���$&�`y����!B`��5M$[�0K��Sr;�zlLT�Qd�R�{�(����*m�!C�1�I�<Fk-R��@�T*�����9�`�CC�ߍ�r@���p����L@k��S��� ۇ?bT��U7L�������]�7���]�{����PK
   �<�X�|=@�=  Ȍ                  cirkitFile.jsonPK
   �<�X��(��8  �8  /             �=  images/02932828-f6d4-4923-89fb-67d65ebd103a.pngPK
   �<�XWC��)�  � /             w  images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK
   �<�XK���(  �(  /             wK images/1042b8f9-2e87-4dd7-a644-1e53cbd80f37.pngPK
   �<�XR�\"# � /             �t images/16f29068-8fa2-43fd-94bb-aa3b1aab738c.pngPK
   �<�X=A�'>    /             '� images/184639ba-f95c-4173-b99b-7b38d7e1948d.pngPK
   [��Xw�'<�  �  /             �� images/192efd05-ebbf-4f69-b47f-23f46b924e86.pngPK
   �<�X����7  �  /             �� images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   �<�Xv��� f~ /             � images/4d249bba-3190-4770-b321-fb8fc027a237.pngPK
   �<�X��НR5 �� /             � images/52cc771c-8bcb-4758-820d-da79c3626c72.pngPK
   �<�XT��"  T$  /             � images/53cc934f-9b11-4097-8823-694d19808ece.pngPK
   �<�X��_8
  3
  /             B images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK
   �<�XH�:9�\ u� /             �L images/5bcf48fd-3e7c-4271-817e-97f3eb0e00be.pngPK
   k?�X�F��^ ~% /             �� images/60a08d3b-0b7f-410d-b1ad-60796781a205.pngPK
   �<�X~��k�6 4 /             <� images/663b53f5-e86a-4272-a51e-f5b809259b46.pngPK
   [��X|�K�?  :  /             
� images/8210dba9-ab36-4d93-90c5-eeae848c0250.pngPK
   �<�X�IM��  � /             � images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngPK
   �<�X�� �f  y�  /             � images/96fabd4d-0b16-452b-94e2-688cfcbce531.pngPK
   �<�X�&�}[  y`  /             j images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   k?�X��$W� >� /             �� images/a253aba3-74e0-4776-8a4f-66dded74c7a7.pngPK
   ���X���-PC I /             �� images/af9fcf8f-e29a-4021-9780-388d342ee2b4.pngPK
   [��X��D>  ?>  /             � images/b521c326-5f2a-4e46-b9c4-2671f5fb6bf2.pngPK
   [��X`�/��1  �P  /             �  images/bc683665-cba5-4f6d-a6f7-879f54c58290.pngPK
   \��XvO�XM�  Ի  /             �R images/c0f01ec9-b7bd-429b-a997-759c27a1505b.pngPK
   �<�Xp>r�  �  /             + images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.pngPK
   �<�X��g)�
  �
  /             d) images/c1fb8ae3-abb7-4800-a199-c8a1e0562abd.pngPK
   ��X��&¿ � /             �4 images/c209dbaa-bae3-4d96-a84f-55b6458b16bc.jpgPK
   �<�X���]  [  /             �� images/cbec1558-c992-4de5-91c3-4ac90e5ffec0.pngPK
   �<�X	� .W /             �	 images/cca7adb9-3a17-4e0c-97e4-0d979b0e08a4.pngPK
   ���Xy�kWq �} /             2% images/d23d5e93-1caf-49a4-82f1-46066b67b28c.pngPK
   �<�X/yR�c  ^  /             ֖  images/d2af519c-c065-45b5-bffd-6bf239de2b90.pngPK
   ��XMi��.� w� /             ��  images/d9f6b7e6-de48-4348-9514-eb3e948015b7.jpgPK
   [��X��@��  ֈ  /             9" images/e8a1ea1d-d840-4bb4-a734-95947de726d9.pngPK
   \��X��>}��  .�  /             b�" images/efb2c8d6-2df1-4fd1-b4a7-6ff478b87b86.pngPK
   ]��X� ��! �3 /             }�# images/ff7168f4-0295-414d-88fb-5470e87041c4.pngPK
   �<�X4q?n  �|               ��% jsons/user_defined.jsonPK    $ $ �  8�%   